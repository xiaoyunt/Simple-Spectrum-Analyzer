`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eGXH0q3ZxaANIAaRJzUbh+VRBLY+VHF27xTXr/RjTeD5XzjcuwgcmBzRfR2cdMYm22s/nNAlUkmo
nGe3vsYX/g==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k5/j/UP3U3WpkypdNUl6vjXNIzKJqmQ+JSlp/eATTRRNSZ+HY4nWVp8I40uywv1YY9MPHs3/tvIi
BN52d4cMGtErawz08uLwxNwcCaJLikWjg9TTdRbux6VyzbBy4ocxHcoS11EME9iHhpNhAV0tkDiK
w8gRamX9L4EccIHeUnQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VTBciBGz3VW7wuy+U7xgwRHfs/nTkshtD4PImrruIcq5+pVhOLRyyTOkIe55KjWVL/GSSDvpqjDC
0VZ9GTti4G1S24b3b/cc3y1z8oL200u5AP+gamj2JtYTk2yZ64155YpNSY+BZEZuh1i5xTwIi0nq
MVtFGl3vb687+f8vcxpEYeOXw7o7PQqwA5APXGHUYk1YSMbjr+WzTjqup5kh97455jrxx/ZEmg+z
Mm1RAwrRhOx70TIrH2qQX8HZhB4Morq5pQkv/twn9Ifp5V1AHRXBmOfF0cx7HwLqcUZYTl40zgHu
c+rVABfQfhMHtGPPU4yfjUK047ziyd08ymjCow==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TwcpDQq2+HgKFiVI3yOuMguQrMFr0KQCkLs4G+qXTfTuq3AgV6bz45aT1biH6vU/s/dE2VPAfDM6
/VJXt+tzWH4EUeTdUFkCVCeQB197PaNX6cp7S0BVvJNlPKlvlOUp4NdBYLBeKORfAWiCBmZ/jRZh
yCNxL+kS5O0QJHb3WAiCkW1nnPRt6I6WhR73PfRk3YvX/S3JD8hIRxa2RDTjimPuaBMGf/UrLbU1
eKu3a4n0Ml7ZcW+vkF57fiEZdBbG8i5MOVw8bSCi26b/sIoQnbO+BfbNrlIf6ROdvd0bfI1FV4fA
2hgkzpcWfrOvY/fTPEPleor4jJbh9S6227EoSA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t5fOG5ULfLV9LpC85o8I5alShvD6uOfwPd6I7/xoS9xWPezOMTlWbU/EWBCdhMkV7mqUTgN5lRl3
TlIcIuXXxb0YN8716vxm+8H7h7eQ9qGVmW6n9uSDchmN/XH7ZOxmUVJXrPRNYqNzVr1IM2IOBnZX
lfBsJ/zwmNY9N9y2Fp0+QmxSRXZqF7XyQqv/e+nvXse7dX62CVSLCcESuOZ4eBhxm4q3qgFUaOR8
F9nthILoLYvd5IaFQUw3ifF+G3D6Jj8pComAQHq6W9Imorr20bZDw8iFXIqlpYU4ECNjkWZ+69Os
gnZHJZbgB41T5oH3EzCPrt5/nh/912bVmr/CCw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OBss0bm0Syj5wzPsl79oRR7ZmSTsZC2ip0/uxY9fZmAb4fNJQJvnsNhZXlqOWaRWvMwVCrt7oSRR
/AlWb+7f6x8C3zQWeUkpVYnni4gfLnfyfmJ9gc60BswODtottkXqIH6tXikFHMbphLNdDMOlkjtB
0usPOtrxwCY/C0PmHJo=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eEzJ1isBWwPO9/C8uQLJvL2a7PgtBCRRJnWSvdMR47Wy/iUGjsqOQzVRyary8kRtwW+JXZ+vYGEu
UDZEA9xJpptDnm+pvdbris5whkH3SjlBN9SQO2G7Hddai31Tr0S1+7c1l4LZKxjpzNaaz5wN4EIq
T3Md8ZQpuuW1n8P3fKpMr/z7954jWuWfuf4rzlA/04T02jorTrldIv61+G+exO50coMQuYNH273L
kFV6cHeh2Y51AimvcH8j23N0BhdTkcORi3zr+JSlLJrtVkGVE851iLjxq2KMf3R6dzgFa567xDQH
e4pEC91T6PnkZMfhjwvuaHJx3uSoWcU1P7BjPQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 681248)
`protect data_block
snBc2OkkN8aFdb+mdHkRixB3fRv/n/BcdG/QCv4U9p8c6s+gjA2XdEkm+DtycSJCKYY1pYLR69oM
Wa4bpD98H819x4pH/q8pp7wNJd+Nr1NSWPMla6AZ0khV8NdXksTZuvx+rg5H32t7iB2KnVkMCvZM
UQMuPXttjZ7Y7VxwQe0G26DXyi6dr7tQYkR17gmlzPUL+O2EhdPrM0GsSlnGLyRnuTEGZhrBapq6
ArnHDQvzTtM5NzWJLLnE42hQKE733fZ6b9Ge6AEh3dHC2TUVLpezDZ/qvTHYQoMtZgpBPILkK5X6
UcJIDTFO8Jj9iRQZ3Dj/1a+S02e09ntOugmGpXmt2z6QqTViCP6qmaFDdxUqrWBkTAm38+hDod7X
NHjPnxLB5oKetfRy3gTd34hRHE3qrVqMMz+uKwPgh78eEnGG4+KMhCYDi1V1GHEfUmAB6tELceNd
HhYBScbnUjDfzdYfb8RS0JTujC14Lo2oJo57g09DI9g8ZNBWcHDeMCJZgZzRM1nyYI6J/zCOuuIe
F6hUBf0IQkRlD36JvSihbqZ0GXpQwXwKoyW30vLobGOdjLfQ0MkG9JZImJXBuF+/LWad46+K3bKg
75K/hcdyjCvK9lyhMxdlF15XtfcinXYoFrgt6bLb8x0jRQaESxRtekRj3+6dzuRLKvtE93H4/p+h
R1l+U9L3x6N8uZmFAeHZKeyOV0ME7AAEVOXLhjzFu5/JcDD/q3trDfFuC7KzZrhMVbWueFBzfrOI
ErpX4qbEJzkszkEmRq9z+q5Wyc53zEhMHdyNNKE132PGAoMYbFTlEW0NPn+IaahM/8kszdxT17s9
RzziHCLx941uF5JctFRuhKCCSxPyHukw5LoCXo0znMa2OkjAuBxMX8trrbH0O3Lv2LtZbFJwEBFW
O4T+94tgp1TYcIVZTcKE12RXlmeZ0KdeycaLESm0COgBItzggXrQF3/tuMeO240y5ZEP2XrKjDh0
uODZxhibLDwPE/GXjARM9gks1gPtIbARscbNB8K24ZmrZTbvoCCsMDuUgaegYyEGH/1csD6r7BiO
/8XSsZluN16CjbEATpueK71TI809c/oP5AdXzxHB2ittd05UD8odzy2NCnCfzBY9gm5iB5pl7UWF
f4my+xwAfQjaOxIDh1p4wvjOZftOx/WfPX4DVDfMz3uwraw2q+/QUewbEvcXs+h7mTnv7nKVZ1hG
3HICySfm22yr2AakBAIHwZR8KagaZVUQ2aA0NViEo0C43piHC2plaX2wt1qlMlRU72L8BdLHlLvG
0U7C7ZeLF7NhCJtau1A2ln6VfBQi+vEtXu+D98zDixIgCJAwkjAt1Z84SAUjkTSS+VhcTptreBYO
s7U5pJFSC/dsQRGXExW2LcmVdgbr+GxGL1s3UdjG0P4bZIx15Gu9Uuv5ya7AIhbtniOFXKnHSDEK
cCtiAabMxu1QLfStXyXq2m0TT+AkKvopruXK+PtOqtq2fZppG62PNw0DUYJS0fpB25An0CS0+Oaw
6bEq9nlCutxV/zHpowUPoG+G/Fuvp7rLdtGUJQ8PzxzGnl+kqy8V60IWsFIc9gixKJ0kR764huM/
SD9uOZq3cev7sRbR3NWQsdTF6w29OeFA8LLuUmGWpRsCl8NvEIfuyVsBOn3X1wZse1I94K6l61/m
XJF5FubKvG+rl57bjXXCzjajiAndVCeQinlshobAzyFiA3ro/HLxM2bc5kWKexlNgtCTZ2dC6Jom
xySvHKSvBUKdTlHJcVh5R9vCqnQaljCH2FyjrU1ETZji21BNrS3xqXGrNtClPnrg3+VF//ky4+Bv
44MTDZ26Yws/OLmt33zvKQvBk3nKLqB4jQlewQjshheLRr6umZIWBy6yUGuT6nTo/Txr4HIYPNhk
7Z6SFG0xZIH1vDNgpCPkiaMVLry8siqV5EDmp7OotP90E/Gov2ICU147mlaz04MV9Kmh50Y0IJkL
/7vrhdj1+Qexk0obiuIhIL6aVLrMba5g71D83gSGygI5ApNjO3tL/AN6iyVqs6yaHCLeh8VAuoNK
LPnLop5DTrYgC8hjVElcevdIfnJbH3A5Cb5947k1oohB9c8U04eA9CvZHu6hRO7U1TMGjuRjXPLY
8ptaEWxtEcT1sgXn2NWcmmosYygiLfD9WRtF77sitiUNiB0RDaasN9loWqOiuUm2YZ4ZkPJUrFI/
IdeFZIUgT3uadNdmHZ92xRN5Uh15NS4oakusmpmeCMo4hB+kcUt9X2V22W7KwWX7Hv8eaUZ9dZ9u
AX7ALhZfA5RTXnAZapVz0b/oXGkMjtRXI+9TFfS3brAele5j1qrqoPg0PFdYg3UugKPjXDJnnwAW
DTgJSejNf3FHcmb8Uwy2RaKp2Yg8yMOxMAWGF3KX5z34hkRgardVe/PqVDGvFzWCR7+JTMqg96S5
5+dzigvbwT2kloxAfsmOlvX5FPKgPS+FJncidSo/6Rgj/XL5bLTrsbSLMCM+7OyNOGRyd3kp02JW
ay456GXGq3ezlxX9zyJlti9EZnR4+vcdieCLsRhijc2z3USvKZtuIr5bmeUCwA9uxok9wWB7/2+g
QohJ2oT6JBcNjAm2PKSka97rJ/Xsw1PCXsQEyxgzjRFlMAQZy1vj3EaiQrIKdlameRzUepI1bgg3
w0qJ58u/vt8Xxp7A29PRf2NofDK3FhBWzSxE9rEW/VPyQzOuZ18oH2wRuQOYEqkyfNFrleLDwCVn
0H8sJj+NYwZQzrfXjcFWoD6s3lOjQN0/s7VCY+684YiZ6d7SPDx4riQjxJ3KsRtnDIngaAvYeloX
qJ5P57C3376bw7yTpij+iw2Ow1c8e0T1XmSA72z4S0I0d0IKMHzKyUsQV1MPl6/R+1eG9xS7oXd9
akrXO3Mp1ijXreLcXn/fvkg9QdjEgWRdB6HZwm0YGhM5mzQrEBOCh7gaCb7QdJc8ag0jovxd5GYf
VCWCfxbWsnz3c9+SYEq1hFINp1/0ajBdDEMrSNWszHqzBXPLWvFQLOvj4v7r21i8GHBv5eB1is6w
9degk3gDDlGcZKzhunxzKuR5pwaoJ5Yw1M2EROswoScg1QU9nR8NMU29Cx8Tk+p5v8kNhDqUnGuu
BI+vkrDc+/2rEz+1KZVDKUErnA23G+owRB/PMGgXqddNz7BzRkAs160/hsrrxlZaAngFEtLQDf0S
85EtvvTKTMRTVL7GOh3nd044hcDLfvXDrPKHHVi3rPQ/tV27u1NN4gJeCEL4v5Wpg5E5Y5IZPgvN
VZutsJU6cgK+Iaf9XkbTi/A5XeN4wM+sJalmom9xg2txTSTzfz+6mXlw3FUGqjV98V6UWm19Joc4
9ZlsULVEnQ3uFozi9he/xBUC6mO64JmOqNAljzXhAoaM2/Yvlui50DPDUIWdjIORsNkjneJSpPmc
CWKY2tQFEoHiTaNCh1ZwIlSL/Ah1eIUGy52D+G61cuxfvH7I0ie0t76C61tedEYOc/cAm8TIm7rG
MpY3RaOwLSQ4y02GcekHqTFlFziif2o6SM5fPkRvsKYFgYQWBIwOjoA8v96unD75KoxAYOGB5K/O
+1rGsPg6XXzmrIUYZqRdX3BV00yMa0AGARiB4gfIoULj3R0CriFHEdEhsT21uBPnyVxW9rtr61+F
MS6OEYmhPFiaK1aO4V7p8mQS3uqPzMZobPA6Xdo4fZ8CXRoSVIdP/APuVx63D0ZznHlobWPSJ89+
fNIULVwAmjk91OXb4+3mpNBhk751v0Pob7uR8gBZXaG0TxYJuiizFZMgFH8FRusbwpOwelmzOefW
/Oh5n9pKDuRoRjyQxjXnlG+ww86XUlteWsFkM8HIykgwh/mF6/ZI6Uq/NL1Nr6PwU95o9ni7tieR
zJdX9ew8gbLq3aTQ5syFgRkD8OEhI+BelZnorn2dYU1Vmka0R/cme/95dQszbRKeZqy2yez88Vpu
Q4ce1HRL7s4eLokDjTUKTiYe4dIHEdXrOw9dGIQt4KwnetwbDwIh/g7/PephCxxHoeRbfF/eGU/Z
ZfMEe9/Blw5obD/QSyUZ3uU9aiCezceheF9yAlMZ0evBK23x90U8TI78HrdPjmDQ0tTQoNXd6Rhz
OVxC4+io2v2gvejHTo7X3996NHjF6I0uYOWXgIVs3iGIOp/Zm2sKuZ3HP5XLar0UkevNBK3eTv1q
1+td/dXVXvCrRXB4YtvCyktgBybKP8wnA37shMDG9ahQPSUlXFffe+GYOMAQcynaF1XOllISUkw7
pcpu4+kDn6d/ox15PuTrL5tKBQfhgT1WFx4+TD/5IdqSW+Zs9/EbYf6OaF+G2CrrZhAXAoi0k1ht
YBIK7jz4oLhJdPCpDPiPA4qtx5c48+9kVRi+PalBwMfx+zAFcjJHGyIDjEAHF30iWTdzagK4MxMu
Fje3FTa/4iHGGZ6PhbER0CQ5pqB4guE6p6z6CbmNiYMvke1WjB5ENFXYA+7U9Em4Ce4qC3TiN5NP
/pCDklYz60HElldrTTA4/NX99KP6cBRESlB+Mmt05zRlPwGHP3GdNWJVDq7uzCAJ6B0GGRGsdM8E
U13VtAwHbXIcDW7VdRQN5pFGQmpuUYyxvRsUAd2UAXc/McdccfjjNxUAJNZoFo80QYRe6IT7wxrt
/LwglR3zmg07Lh/yyjASea//3cfWtPJlM5RU4RWIV5IaEtM4KcRBWIjzH0Y5SIzCFSNK7DTYnrPV
ir3UpoHMdOYWm1TPqhJthZnlZJO7vYuXrpOj7AhNOT3moG+3fO6G1XHblr8iOWfqneCl79iGVVNR
BInfPs5wnw2euKm4ZLwZNMWuMVd/zk0DuXvhoUnS3opZrazkT3EsiM2Ut5U50DIXGCVDvzEWwBhU
WC+VgJCbsyi5soNOrzknDqPzO0PsYh2L3qf+5XKuQ5PIpIh7RsSV+Ot8OJRhs2BYgGbxAothxgqQ
eFa/Fy4D0QM/BBdPD9U5Cl7WsK/OsulM6cCIMKW0umoJxnVhwvSy20FIUUDy8Nh19qWghsGET9p2
LaKUBsiuj1q8tgqK1zXIZN7vAp842r0HYtaTPZ96fVRpNgAD/FkZDEFC2q1UHlXkAnNxyEMMSTh9
vaIyAnmAi6baJg2aQNu9aVawPSdtimnhNIEKAYnRjunZB5X9xNNtagsnvSfscfYxg5yUnhgHlpNA
Y/aQIIoO7mzU05SfJaX4SZcoUz+qcTCnz4oG+wYiXrOuWUpEgmunoroHsFXLkViSj450sAZlut2q
Rur4XBrSox6nf2j2sf92APaBWHGKIOUZMuq0rgo2HXLnCPnBezwwQgMf1lTf+DuK9ms/SHrqVI0m
IE5BqqRQsH/3qRcspPPRSHDKHhEX+uO1TsgMoq3IsqKoVwFdDedBj1zVjAsxHiYZyYAFuX8kA2eW
LuDGc7f/mVPHEFkAbrxXyqfduhLcQcbRe3ZSk434KgZqPnxxyT37Zl3Y+yYRFKjf5le5iXIIlNwo
YJMtc5CgDz4FNZMv9F31+doJf0ZWxZhNgyZfqY9i/6n7hqLHO53GHtQOuqWE88xoBiIOZ9jzFDso
paopQ9r49sIkzzDpaMYhwKOyQHcou9wZN0ElsnO+iX7KbLZPR/kcvNFhpLDw2zgZyRE9F1b7wSy9
G3FoP3nncQX1mvNr/VEUNQERTgrqaWjPD44httrboEKqk+DdXPGc4ZMfnu+Kh/b/sdhSQ3QVfDRn
Thdm/4SmhJ9UOKXY2LbPh8G6tKXR6NbOrhZ5IBan6oKv5CI8El9JgBHmVGoMqnNepQ9czIHddYJE
gPIKbnLxfhpuNtzviqQrviVWJvU/ob7zPitxjKW4olNlKauoFy8YfL7uUBVYak1IW8qpceQbVnCD
/ocw2YH1D0V9NXAP4TUP1NJBDHKkjOeXloYLFf5EIV9cT2z4PtwO6DWwTDUhsiXy4h8JGfTiUSOY
/sSU98g/vK0JjRTjrQZyccBgiCckYNc4ch2Ly6cxuajLwnnxLfm7pK3MPijNB+xILRFXxt9f4psq
wOwEMNj98g0eT9KHJKMpMKfqFo37e2MPY5Ct+xKqoptvbIKieX4C5M9Hp8xuOIEgQHyb3xmeZNDZ
e0bN/3KsOwy7g0MapALPIvB+HCMoREBbuWiGM33xWbHcDpSg/tb1qdAvDvNx9PiJxtiILzTeHj8A
m2UVwPfnuEoBISu9qHogkSvnIuf/ViRvBlZ7UX9r0ZWJHlUrKanS0xEgmqWFgFwFCTcyko1V6tLs
4fmYE3JuORjTJA0VwZqsniSyDWmH8J8tE+QF1WXV1Ibm4Hj+sRj2nCML5X9FsP5GgBy50Rr90V5M
MNkqzdMpKgSRutaNCPQw44ntsdS0j0W3/WyAoTiNDZEX3g2h0lZ4/Ozx0XUuhGL2B1jepVdVearP
FGEPjac/JDhqglW3dQ4XWyDQceI9kitVgOZ3mcCxqRkFS1E92mQ+oRzSVnotpJoX54MuDyPRNDjD
/UvURzCuqweUAP5tvgo8IbC2UWKbwDcdoBDvZDUb+211yXSJNtZajm2CTeAxvjtSozBzag03/+H2
6DvnUMcfc/qymTbXEqOzBf+FHsdSFATcjKu4dsrfr6PY9NedTH1owu6x+GXRzYOyeqNW2LGSPitK
E2cIy0/awckX7/Skp0ql4V5IkWRZsIMg520mbbKqK2kqz3RtojA1HbxD0VctmY+O35+fe40zVQa6
gtp0/TfTiU0mmWb9MKaeZiGGyUaJSuH2JBEDXaXflrIux2M4wgd6A9EFow8TIoyxu9HyR3Llbc5A
ktUWSiYm2XaMtmLQMEKJ85at5d0oINR1m9Y+xUoFwWgwODYIelUZKdQDzcvdwP5J1BzOBEiHTX9f
NDcifSaAf5n0NG1ukf82XGC/7Ofg8XOqJitAgF/BpzDyLOwzgG2RRAGiJgzo7jZBd+2BkEqkPCul
0NRPUO36WSIOMuZdiO7yjqGm8SDE9OBj18ztsSM1hsCtMcqsnE9Fg+LMbuAhwZuWS0Vv2Rm0PwbX
F62jJFZykusQJWRk5gVIzYqeVcZZoSo+4aBYHeLK0U4Lxq7ADPddmSWN5ycu91kFIoCkZc/bz0ve
bBhphuyf6mqUxx06s0DEoVEZ2yxrlT9Z0r97mVhqJT4/vBJbVGaygEJ1EC12DlGzi9Pu50qx2yEE
gMtlqDzP0NAiG50k67MEyKY/xdn/U2tRzXTu0paEQMUFykenqciyz4HX2gsRs7QZrBXPlOY8Da/a
FTK/YjFE8radxEv0qDbkH62TGweF3AcyqVned1TJOfIz0xbSr4ZIp4Scoui8YBHwfrv2ekM9bVb/
r18gM9+ZczBQ9gq/9XsdlzJZFu12hzhd36qHxUb0LtRR99HmN0DWhO6hldWV/9gFilFl6W0Ox0qK
PKBrNOPcNwQqsGroyJMGLWXlY+TXNGP8YRGicZqXR3Tu1pxISq/aARiZnlqwibADPsunnH42M2Qt
WqmgLwRMsd1lpaQXBoqrLQCMgsK8DB0lgAWdOZ4tHFagSVnXSAZ2bLq+qH1nRQraeUYwfjgs08yp
m0lITCWxDGuXw1CjSidjSb2lUI8MLFaR1Pi65jMSIW4B3SpJfXunx0ISFSjgTAPDUudqDHRK1vm3
2VsKW4tGD8no1v7jjNHqxgY9JxFRTbYX0wKelsIxrVTWRWxBWoJiPEVpqmGfM0++tyI9QMMQfnFu
ez2yAu3ZoonZpeB23Nuf/TEctzT0jUAKiSs4YCZcjc/+5fA7AoO12kikyXWu1oXtlqqNuJvqCxcR
uDl+79etbzlCnnnA/ULd7pnxWosNrAxDV7gr6NYEi7aW2AiCidnYapSzGPRexnxNDuD31/3sn1Rw
XdP9OqMBNUoN9UHRGqpRZy6gw0b4uH9xF1U05gbapbkp9fbNo21Rt62u/S74v930k5xua2naoE1i
nXSmfFQhpEjySkAkCplL+q8+p/IYGsDNR+lq7vDm5hpQcoCWdTadAmj0KD7h5PEiC2fq1Xm+FkL0
Xgh9ildfZRi8AetvYL116ksTc7vXE/dAj5amUNElWc+6i6+17bQMN2F6Yw1C5Bf3YzNWHsdEG5hX
K+ILszGdhoV6ahoFQYcQ8fI/50jjcmPwTxi50iF641BhG1Y+mJspwbUx/pncwAvE8w1WqMzgrn8w
mdj8/iriMBZHv+MsCF+pD1B4HaBUU2LWAwBRj6xuuEC2irvRQYScbmZfFDIksG+ArUPL/cYvCugU
L4+xdatrKzIc+E+K5b0oM4Fjdn0FuxX+X/VnOV8tOmK9hlzx9YD2n6Bn5pBUqdyhQTxLDTLanQRN
2ILp8VMN80lq34P/VWvITOUbJ3Iq0DENrBqPRjSxMgT4qIeRD2cXwLg10ommdjqECV6Fj3h0ZpqZ
J6mLPek7LBbNvYtYm52cKGJ+SszQ0ALz+KkTcIKz+IQqxOrqbiYcLVwqIjVxAMcpHniTmBe6AqMt
wrMyI8E5DTUOi2VQ6UA0utYo93utAXnkw7tbiBMGLvMVJZGYwW48evJPrCAwkX9A9RykVy8dEyT0
FWt+zFVMXsHEAclgMHXhsGG/Bn9mqBdDNyESIZlnY+BtCRVw47BFPdFLNDfiUWmKNuQZgdu5KmMb
selrT9FOUWALh7ON+NRi1giJBUtyeq32pn+K0ZuAfFk+vQhLVNJ+U6JG1gmgxGR/GJceR6/TRRkI
0DbXN3/pBr+o02VVqfqSYYSiyOw8DKR4EQRs0Pg+dsif8xRd9URkzD0Uu62wQTUNnBONRUZb4d3s
wJRGywdbFMGRkuBvt9e/Q+JbtP6ViViE4rK+jJjBc+utER/44q5OvyxKgRZuTWrvgfJXynYSQjzf
S9kUg+2OTzixts4gEpi4q/UvysU39eb6mNGpfZPp2BpY39zOMo71qk5VdGmmows8dFxgvayIZ/ti
Lco/nv3u5PuOX9mDVOwu/SWQrJfqomEAZIQbuOsm7c4OJITXmLAxvIGFMPVR+GZnuQrs25ynRdOH
skqNuaAGDmNLq+K1WYevwAMaxMxmoN9IckTuItCLrFsqtwDdwaupCQwEnvaSjdldwaw129VaMDCM
fIMNtqZHrI+L0NKOnf9wT56MYrZgs5AhXew3tBGs+jNJW73a+CrmbQ5MTi5YkKY+XjeEjlC+HPOW
TLZTtQdWIQI+yJkwm3RM7RKOvdVELb5Q2Cxp9l+1qyQB+Lsz/GrEKWUj9tWr073UUpqcmsDPu92i
RyNN/QB/71lOIi4p4f8HFMpao0xpqqbPgZv5rquOQ0AAWP04QVYDBe9lfKY9SrdEMglFZTd98uwu
GYaDWRE0+0Da1fTW7cdj5JX+qKygyZmjiOpf7xfx7JyXKZDZYmVWMFlRPA6EMCZQDb7VEkYbkYDy
MeuKV2dvts2VTw1GaNhMyblpZWKAny7ign/L9xxIUqvD/8xUuKrni/S6B/KaW/VYmgQM0XK5XSpQ
qMy5Q/IGM0ZjWKdvNshLNi0zah4QMrqietKO3qLfWDlpw6xLBk7+V4eO95PrAyaSMEsoM6dldiOm
PhpqehUVeB1qXVQd3Iohh/r9HH719nmIsCZYrj+XRqsMyVUpleEjuQDOphcuSLBcXa28Zjh2kdY+
A/g/d7yP0AXPpCkbR4kUeq+dCa96EYR6ore4Javd8dYVY9vebUhQUbXMY7Mq1jvr5FUl9t7094uh
Dbx7NKK4WYhvv5Dpjd4q2imspuMAOXneX/W/LW+wNsPJBuCo97tz8HMaD8rpoc7pvVGQF1ZkSDYi
u6uc9x/tyVftXX+HBjJXpqKHB74+yckbqhTuzatxJIvkWH2QBDNoS6IshSUOe81WtOcm2g17Fe4a
z3K8y3ipV6z4E2eit5SYtMko7eNUoiTQ+Ef8YGoEr4CLeVxQcWFxj30YZPUSg7hnZXScr1kAJ58J
+6TgHYl0alNHI+wp7tZnndWPKJWHv0jEZe8s+1iKVG0G1aPc9gcR+Gx+EQmHJfcgtJ8NLdK8Hpys
VEcXfl2RMm36pfEVFIj4xRDHq30meXQOgZlf4PYStjMngrvyKXy//vVgxwVR98eka6OIFx1tFk/9
TvYpar7XAeVrLSX+UWgxbmAAzsMtKI5ZOQepBhYzNTzRX/RscI9NnyPHTvWztf/6MRPnGFQUBK5R
3DzTMbpMMlNXg6pVSRlVeHUknCrnntLkLIHWcG0jh3ucmmt0kYhFW8ZiQZ0JaVTbdHURoN8dL/15
Sng6+s6mt8mjOhfG2H/LtOQrZ/YPq+RQZL5icFTf254UdDLg4IP+2G9ldtzOCcIgIDU2D1Eq4lbB
i0e6VrQ6tXAdy/thfArJbsZ0EmHYr1Y2gws+kqTkg7lb5kgelcAh34Cj6kcAhxkwGIxsb/EC/yj5
702OCNffLnjZbXd4B5fju/z+knlRG5Qiozq9O3Ld4Zpa3eZbPrFeQCsymRZ65lVprGbU1eSIAURg
e2zxmZXADuI59Y7VKoXobtfR7VOId1ywknFYmAD8CqjejgsAePq1MN3kp1CWJ9Cg2UtZZIkz77vs
LPaM1pHjxYswcaMV5TGf1Jdz9J09fTs1Gjkjsc9uj2vO6vfZz+ZR7KeMGNBiID2cBA0kABlrijIJ
c+ousnzktxAck2lttxndVdkV79r1mBDoWq/DQrcG82n5v3G4Mcm8iNk2yer1FsqtL1fDh0OrG6wV
Wgd4AKJAb9LKaJ/6h4mTRJUN7XtBDwvAo07f/LV5L017qJNSt1welX+UH2Tbqdm+D0pXxoqiIHph
LTZ0sDW0MSI5mzWoid7rxsT6jaiCNJAob6WylOV4nJpiYFNq62GyDJ+rkR5PccqYujVujJVZhspp
PKZmiTEAm8EoPdRfSPJT9yR/SDDwhDhQhhLl7BBaTO/d8nu7+RKFDrpUp8MKjlhG2IvMEa0GLnCW
pJyX4OQlvdjIdk+4ta6/qXW7Q8wUr6OhnIMtpXYMVP5DItbrUb+Jn/Lpcmzvi0sPLJoYqCx9SAQl
KNQbnCEBLlTf6byBbzz48PENKVnoGox/FcW8HKfBG0SeSmPffMQ18AXRncJRFxSJT8cmbi2Iqc3b
ZY4pMjvJzFzMT8T2I8taBzPv33Pe9LLB1ha34H8bf1T2ERZqTJmniDLD0DWic/BohIZJInQsMRIe
Ft4HZ+NkkQkTYOWZNarCSEwE0bLr6YYXr24IzsLWvQX7R9ss2E83TPxzATTgj+KeWZoaGhD91YWs
tkwgZ4DMBFLFoa+ZIJ8w8xK4IE7AVn7oEYklR61rJ1GnUOveJs4+slT5eSx3+hkUyxIK/hzsabkp
BHw+Mla5w38jOqx8PAdF4RcAlNQ2vX0dyDZR65YEjSk7dhwq6UgJybfGCJZoZQMci8zKla0OERf2
MrSuQNzvV75nF8OXNbV5SIGVJ8HEeybp69MLVNK3tg1yyvBvJ+ZwfDPcteeB1ktJ6tno0yTRizHw
9VbWH3iNOnuxoNJdRu5rRkVoWhQaFnztwLm/tcCrp3LWzNPzqu9nAPr5gH3eozrbJZX/2Ppg1Uc2
ILn4mVIzNvpISD7YLAfEIwrQwT/AzBEYbiVWgkT9Vize3YpPaj0asmmTDACc+TnfwASG+Dh4uXwP
t48HyYYdQHAboNdi4dG3DV/zvCfSpzsiRS1k4lSLjVhqF/z6cY7JfN6fgObQXlCJ8n1s6QKIYeTx
7OBj2A0yGyVHLgSvF2t09ucOZO8/FYCfCc9K+dW2kUQQkOJiTmn8wsoMSpbP/YTrMVDKgH07Q14p
GfHDfIKl6SNcUZfqQHlTDbcLrB57a9j737+G+4oWDsYy2aCQ04YzalC94aF0yIUpSLBpEuFe/EOm
AVKFP6GjAbJuwBWoRAq7P+2n0RE99IjseNmvEA2bQ/BHE92z74JMm0BQIRQLb0zU+BoeNWS+7avc
RxMC+nWB5y4PPRCOIyI9vwfTxh6rOIy7WFrPc2kU723R9tDDTVhxTDTdxFMubaKma4oWo4BAVNhV
EnwdmJWltkRceJ6DCZvI8B2nZXhPW4kKOLdn9Yo2YAXn3VawwcJjw7SH+hfY2w/RJmjIgd0Esme4
NZikxpURZT9/uormOmElDVJzfE3cZUscJf4poY0uJoRuXoGH4JfX6iA6da5Cr1kujoRqPt78wzmN
T2BiXzErktdvvFLUw7tg/WFhvJUC+7lnKkFKZquyciQwYv68GyYxo00G25bQRXvMOhOww6J6faTZ
5/3NfIzPqJ+Ceq/r7+GisXw8vzAT2wd2w8WUjAHCgu3ZaxkHamWf0AoW/Xne5PQ+fx5BtEeoJbnb
DHhlsnocPFZ+DVre8ttBZ4vfRmpvAGuM5s8upm/8/HzB5vnjNCT8D8g0DTEbnjifP71zzx0u3P1P
+R7zTDqsWpert/G/bFjyKUEsXn8+VASGzlpsPQyeZCcy725aT0XeefS2bVcXNfcI8wc8Q85Q/El4
MaCXwQBHYjtT6CPcp/TsLJeCLPeFBdBLouHQxDqRzGGnijilel72g9cCO8ehTZv/sBaPbhbj8wgw
wbDiTTp59TymlILVM4rXbGbbtyxKPdLP4YH2SihUMC2BDQHjXGIG/ZGR9Ikq4eDETvh2fPL88U7x
BCIBrbHBs36lKBdIxiovlYCeqinJS4hX0aH+jdV3fGWwXscfFqOe8vcwz0n6OyA0+/ufaGEMurwv
bWpEw7QSZXt8UC0AwOq2XOiMdOc406W+EtsRuHA661IGSGUMwtDc44oUwfTM+6kS7by7oXB0vWME
27bGnT4Oqok5HrWlLOwgKNObNd6pMX4Jpk/9bYDcXBvxid3AT/3AfZiuVg8u5VAJz63ZD/WwiktR
psTNYp9qNub1DufXygLWcOKKyPCSRDEZCxp6NFRmtEebTNbLW9ZskOuGPpVYBN8MGX+MpkLjk3Mc
oxEv50R+6aTIngOBQ7xcczJu9zWXVFkWzkQi8UgZNRKzWoHXYoLLuk/0J2vDqpG+OASeYCpUrfq+
dRz2qwIyygfYHxhsEBokJelXG+ZiF2EVrKxNznde++xL7tFfCOmkAaWf6CXe1dwWOWLg29dEzzQ0
yjiAJ9b9kAOAHKVxZO5JGPMwBZDyH5tPa0Oo/nOjQ0o+wQT6eTr9ktxpTJ5qFArsSEs3CyHum+8F
w/Pdtane4mkBhJn5pD1UrxpWhufhC0l4UMQoOwQRupa6CmVbJvh/Xbq+n3uxyhRCT0pfPBPtL9Oo
sX2Bl+K1kB3CDofzyvqpDXVscziP9/4pSNiZEfeHffW2PsFVyBud4QAOMeugC4UwEmQFquOkiQmd
7G5o/KY5UGqxoaYK5WFYCc1m/0uvzNlCU0//288FUWKkV5ifhvpCWrX38/HGeKB38iy/mF+ExAZc
8/B23Axy4Rg1SLIagsgyvYYS6ZCMJSCXr5TYfUNTg2gu11+PIBKNYoanXnZSt5ZTadTR8k2oOHrs
hZ4v0q2XFERuew76DFiFgf3P7j57et+easPGAvV15RQmAHUvcsya6F0clpavJUSV7K5ZvGhjtjLF
xTM+1qhH44S3KfrItQSuysfxZeZ/XBAgdJhb0J3xPjEMtiB/JiW/ztfqg0iQNkFNzMkRuF1jVyOd
pfWDddU3kU/gSLJBylVG5rDO1tACO8lmhFKoDdaTbtkc+LY9+dNzZWQv43xuXU3U7i9oNvi4m/8A
Rr+vQ7QRdV6Ax+QTnmvTXeFTjhkGR1/xFc7Bk4pkkyg/xG8g4WcMAP01OLkwx445f3g6AGr2ApUo
nOr8we0tFWafybJv+iLk83JhcBA6jtLXGk5hK/tBeHKMQ+FR8ySryXj2ymFX33GjBlH9N35cx7CE
4ADyT/Gj2Ei4WY4YVCYdykITZFWdwBiXr7A+heMyyQM+KzQhAdjc9+ulkkG6FmGSCUmzTB7UTXVb
7Z9VLeZumbOdAsJe9vkRyEKBs7FxA8C9pcsxq5s/KkSGo0bfrc9rbY7GqDHoP1MfSc2q2yAeErCS
YfrqrbvV0djbU0Kfcienf0cmwJ0NxXQBgPck2WsqcV5ByRR3WYLvDVC8+EHN8XLIJJ2klDAUEFO8
quLzCXD3W1ww5XUQ0Y9xPY9KTwILvO/MEI2EQi0evh96tL7ZqYT6jHuwfDeB8XrGaxT5ccvKGPxJ
UO7KmQIU6rpBlcyHA0nv4GlaOY/n4GVyM+5Y1SCc8ZuVray/53IrGlWAY/m9vEQefiTpGJ1lnC1w
pwqTbRtKjJO9IztGHBTWZs/DXsgPeZQoCYbnRK+XAf5d/dJ0Cm8WwOe3saClwlfzVDS91QYYfsZ9
6YytKJmUrqcS2se31KcmXupoUbuTYofWi/vCrzgnwCz7izbUW7OplwsudHgWuy+Hj9Tq2nSo5OTl
0v9gd6SbovUXKWULo8Ycp0FbeaWMhLSrbtZyoyi8+yGSopuVyugsGRDVPfgIig/pJL6PWBktb/a3
dyVB6+z/+DTaehzzUDq5QdUyCUBj0hy4GrOaUiTLcbRDFhFkh3UffPLfkZRgidvBtHSrLiIW77AG
hxbEvDPMy7tv9AOLxX7SrlYLx0yxt2UaQtL/uHtx3n1wqDF5UOHv3Cbnf5O2KQ7Gn9WyXzJI/e7/
MKE2OL2ncFIxGXd7mH2xEW6jLmgeIdjzA5m6kQkwyl0S9Bm0wrP/7mUWNI3uESa4l/bSCgVOAUZu
MMJNq2JHfHu+ar0XCo+R+qrXUk3a7xE4pDURIKMPO2Aamu4kcefG15W1gmlAOs+Ia6pN2FiiRUZV
EotpITPvOc1hHCV/p1ta0t4T4DmZKVIWLMkhFl0jEJjJAoFf0enepGBxF0rPoizWOUwmZAYEd+nU
ckERi3GrHIx/bo/XvpmmS5s7cu/EmKbk551LwLXlsFBeVvHlBuqhrniGSGLa15cLKvVHSr6xSnSW
QxRVY9/c9LHtZv+1Ieokjx0A3DdsUqOWZ5PJQcV0qWwf6jIAwSXAz5QL9BfqXDVxpKTpvmrnoU6b
FVkXfzulrOHSx2DfevlUE4Yng747WUzFGYr3CiZYNBLVDMVnxQpkm8N3mFlMIJp+dvlEVPnAYyoT
1KGjUJF+7sNfva4FiI36W3Y2xWhB9uCSdnqloAtAVBxsz06N+KBfd9nBfbTjpJ/ZXWNrYzSxC+Mg
tnytauoMozUTcWyGTeOC3a8UIsN0KSxd/yWBT0veUa2XZCd3ut0+EipOandZNiyKZmWnr8ToZLF8
SVTjJh5rDeMhqi35WxQVzOvP5fzj7qPKijACwK5zd+MQ0jN7IB0aooMxcqU2bSkJMuQ/fRDUuevZ
D1F4w+EkJvyZdLi0tFW3K9JxFd6IFe+6rNrUKCCBYX5EmXOBmlaLF2dcqNSZxVVA4zt0mO7bdjsS
+BZfIFuJD8UqrvA867SCeRO7g0nkwS2FsnWVawcNuJ/mGzMwd6v7o1k4No1oqRngb6zlXY9hUfRj
LieAuL+CpGMeVKK1qFuJrZBDbSRQDni7G2YYG1parYB1Q7HW1XIn1WVK1c2riqrtTutyKhSc0tjh
m4B7/jX/5Atcj1BUWHSclZbMCs1xUh2mfK7oHkLY4mgCq1WtL0R0gIIsAFT8j/z4w0Wbw1fSgoin
mDVPqzKbJq/bRv1KZiolPgaOvntD6B10XVHyu/uVS17s6gaICPjG9kgVmhPhNHFY59Bsq6S3R0O8
yxabWGBexKtTfqqnaah6luKNbd0LBrGrnFCQjttXu+mu0NIQj6eWmadluadWXPHoS30hSB5AYgjI
nLi8yDOoN760YIL5tZ5GNVgTezer1ewRNW2uJrZ1T/AH8EJ7qvfhmv2mIJjeio+tuu1zlPlj9wX1
YOlkWqSyWe/v//UeVI9stSKQdzXFr8Ff1x4u6PHDzrdU1bMqCXddm2697PFMc2EV7aB+zd9w+DLi
1eDkxGRNq7LARuFYcPNpf24tZjjqlns21HP3tHvVzo3zstKQ7I9/0uTIjWRhd1CpqNAgDC+Uf2bh
DJaZwjA9CO71HM+ODtua/A/HFRKbhm41DjGEFagNc/28K6nBqptw8TqFW/MkLPOqqqb1mDsh/yDN
Jtrast/KfSIb0S6ZjiaGAM9aVzaCU/sX2e6dO9gr/R15BA5hKtb2Dovr7ndHdmjFQPlBbVTZeGK9
ff2URe9w3B8+blWXy96QpfVahK8AS3zSlYlN5SVv42CrmGqAzVFiqG2Kr6kU0Zm/CxL/P6DnLMdW
eY+i/QNH3/h0F0TSiFOu3tBtUjyQGJ7xw9CK7Vz+HVvi60Gv91rL1he0muAvy0GLTrNLbi5d8swN
E1ZLZBI/gASNz9ndnoRGWy4axk/6i5XY027z6oxQXELoehU7sSlTn/DDvmdmoYYusUv+KWQ/JeJb
UuY2PsYSLD5g7/gRhnslXLZxIguZd/mNTenagN0qF3iv+oV1+Vc/NCAhQ0axvj/CCBIm01czqM+f
m3IovHi/MbLA6t8c8EB7rKmo0UVrFpNPFvYHt+TarlgrLEnoPBbZ2xAwvVhVMfy3ieq4lPDQQAXj
EbKVOaqQIYD6+lg6MFR78yjo/PyUM/oytrnW2Tk0KYpVLJ2qkyxunUqKxBmy6VxI68StLo7MlGuN
/0ejXJsEOZ2Q/baDhz+G8aJo1ghbTc+dPshiybHjjiCSJ/VujaqWfhBhPeo1MHsszhfgYwP8Ri83
Oi7H+CVdlhbS8uym/Ja18ZnCoA6aG5N1eKUXMbo2P3cXX1CFwKl6aQAPJ/96fd/xllDJPFH/6muz
8IKOVm2ZiV9P1J7TJNXzIDaKgHgQcs1mIuLMJHlmUya9I9uUNp7ZZsJrjskeJtLMtEg4fRCYouAT
giUMWzgGgu7qyJ8ieRGg8CgSpaBVzuLyPEhF/QEI8bpjumtfq9VgWjFNMY0HK9Hxec/WAuACbbir
K4DDHf+7RLQaFODTq7xoH1QnJx9dnUOs4grcg13rCTt9nRFwOGl4Tf6zpgEHZg4p1kiAH9U4hkVf
bL27fEyUj98uiEUuDo2LJrh9414KO9D/ALB658OLxM8acPCNrNvtpjdYXRLviowYe7vNABomS67X
wbP/oHPsKxe+0jXZlz9D28yJ78l2Ow7G0DTfRT+Eq/LgW6bIiwsOzhDEH72TmgPpmH+LjqbkC6bp
KXpyP1wK5IOE21WagGoZeLd8o4XhA02hdAt2RnL/FOJhxHFDu8D0ecBSPsJLz6THa/nZu8HoIPP3
vrcQ9986msSoD8c94Ag66V+2p9vKZyikXA/jVCk9evjH/YUO0DaBhrTm89lX/9F9U2Okpe/qEGFS
1hTVIQdK8WW/0UzYK49+y2WxQqQ6mVf8d65FjlcwY2vz7Swnkz6Hdh5wEBAuY2wNkOBoTVUUXT6t
YmjQr66wlsS4SXxdTGEIkBdo3jStcLa8wgTRPklOQcEmtEeygHNIfbopJNSrbnbpMpZfF76fdEIT
H7IxssXIY+Rf2vh7O+gUryp3mxp8x1oRGI9czV8AjWXVWU05rTJD0LsxFmEIOf8CcplUYJI0X4nH
omDDyCtFwksiEr6M64IExweLXxCAo//UPoqW+nW+TrBh35e7jx468jEmPRnwQIHSPzoO+yrKVDZQ
XsqJC5nOdAwRQf1Exlix7Bfg6rqn6KqCSfIStyU/I9zCCJK/NTJOcu3X8ArkwLXb9V7GRBqMiCSf
/x6sYBJPzupnZdGEv0Ouo/9PpCMHPo6fRYs85VLVMJs2OAT8nzLWRSnXXLyWk5Gaje2Ycnvm6XLy
Mil6nbYZaAxafFIwhIseHUk6d5cNqGdrRfWF+ajnnBCrz9FPo4WdUD0rOGDzTHpe357QZW06PfR+
neUpO+p4SQDpeLH79w2kHHxSdGGMxCH8DfsAylacTL6pzUI5G+hBRxSsUua9vzexArKwTcR90i1u
MB7Qs7OHELiDzl1vIsUH55yNGG76SrUrCT8r3UMIGTlYs0pPOC+/j1otmpoShxCBvw4b7lw7Zfla
DS/9FWjdHIg6D+Q5Z9qePlkgEVuDVHxIm0T0nH6qzaCl/oITBprBrmxqanKTG/34SioLUuoGmanu
5Y351d3QJQcRbOejG8zrlaVoo3cOq6EtWoOYhjx5gvmS85/BMIJcqx6d0xvrnQr0/ebhpcZUG7ny
8g73dDBo84KgFYXIs04BT8BNetSl5v/kMTZJ+zpXIhsVgNm9k6PX6cf0V6idJtLp6MCGn40C5wPm
T6ZsWrKR25ISUI64JNnYfKtwTVTvTvsB+zijizNR7XonPlEsqLhkS8LXANt5zEMHgcgEh/UCYxxc
Z+OvQMKnqRw4xDC2EJI8H7MXv4QnpsPBRayDPaNNAFRWQ1k2OXmd+qQJcBTedovYh+NmJxYUoM1A
PSx/Xjcq7ia/R7QLczCpBvJenIUdUY8wbPnuGXioiVBxl9YJJstCRRmokCokDEs5ZHOirbwmhMa9
joa3BQ50t/HNSdAqWA5taICmSTpY+fJ2W7AzcHNf/XdSGereQdZEr9r3duvk5l7THdYVlHiutQbG
+YTcwLMT96bYFaykkhpqr+JzY2bexgSUtquKTbGZH7pjiH2d2MlTJhHEZnKOP3+L1oDulR3Kbup6
mu3ZWQyGvrMwgsk2jki4a10Qs7J67nJY70Dgeaq2MtYKbZs3gdSfMxS/KnVYzWBP/GSufpYnAWf4
TBww+1K3K1PcMT8LkoD3NuUQGNKhZnbk/fQ06Lij1kyFnBphpSjJauR3xgEzIluHIZTVtL9YIeq8
K1634ZHzcZrujvNypAGH55ZQRzSnIL7LAx6YlqySwPE3aMxhZrwwx1u6MO6H9BgBP11+v5/oEoaw
kd829+O3L+IOM3kQalsYWut6mtEZcmMKsA+WjAAzv9HmcrJxeyVpeup/Gubcjz5uGYnL5ZqCArN6
UCLMO8HxJiOJnCfG5IhzP/GLMy+GOfI18Jjpp8+/42cDEIPcRfamkstZnj1L5LSDoMi/Maz/pHIe
S0fx/p6TaMdcF1KkegnpMdzu+e3v7+T5ctH+KMz5yts517tjmc9C24u+gpMBaMP1JXaEsN5rl4GT
Df1CehCs+RTZL+WUQMR4NiRKWVdUIjeetSOcCKWfiXdanPvMNZV9gUrPDn9zl+SdDS2BwdIT42DG
k4WLYzOxqIkCT6uGKkVvl0FWciniTzjpsxKeyvBr3kTktFqH03ZRnpUFxKiGlZ/mXlIfqlq5B1Nn
jSaND7F4qtch11/rbbC7xbqr0wwFGcSN3xV7PeVCFyh48rrkGdv/eW6JVKIWXrbzZ8vPjfGO9GWX
c0aI6ppq3LuQQAzg+AxMKU1vBhGBJaIEbdXtphy7eC79y6jtwU0xQbZWaRaor3mekYYEdNW+e2ZP
awbNKUiKs55HSWvwp18B9mJp+kvOq6pl+t2WuhugmpNlas/9sXjh3Z+FpzdvocPZci6+tbt7aFl8
JSw4EtE04OvYzNVnOO7pIGJuKXh87cpp/mCifJK4rr/aHHcmXoNaJztdEWnHCSVCtqdMTt2X/umO
4z0JW6CLCWq/6q259/zqa0itoVsktT1cPXI/E1uiXgU0kUZtkU/oyboY3rXu0CTU//tZ6r+PRGws
myPLnXjNiQlMEz9d8nMVdQ6/4vkTPqjDprayFLvMxxdarxcwgpVs2xZ88hjJe1S2YVmQOi8EEiyO
XQN130lXvutKpT0j8v+a7WJNvE0y4YL75OQivSWvvqnoO/ipe3XoF7mpa4FyUZi6tP/D7HsofEXl
zkvb3SomIiBG0w72PCZJ7menRUJQWjA6rwvHgHu5/bRHEolDhKg4Gsr1ny1wP1UJ80KQPBg6AKZK
4PsoMIqKrci66Cw7+Esnb5JFzwxbRb5i/XeXsO+RbaB1OirANj+d6GuBaFujOamfWWV09BIpcgV0
bhZnuXCKDqE5nUaAMqGAub4/5agZ2tZPNuE42JUfSJzhEf/5IQvKRr+gJogu7k9UD6jjQkOqC8BZ
J4kNh+gn5yFf1NhOkQxlbAX1juMsFn0OIYg9MKgGyOvApqsb/3GVwVDUY2Q/+wdydHn33J2+YS4k
iyIzgRF/+lOhzYtG3szaTJt1Dq+lNKbmz6AF2GtECfMquEjYWYFYfRqiBfhBT+TihiA9BIOq/10z
/1zcKapMwdlq7oP1Z3ZNJfV90VjOS0u4WUOwRzn+S9C5FtLjXp1UanJJPU9gJX4OE/yvTUF6mghu
vbPxz3N3yAA8qrIhj3c67rSxewzIvSuZBCkq5BIkXZusHoYVKgyNiWJKD69+q/hO0BNYmdB3VOY9
MTl3jzO8GXLxJWwo3vJzUnIb1mOF7mFR9KizyjOHkb2nAt9lcbncxrt3a3K8to7nOwHQv0gb48SS
zd1eBSRPxgJQpl8b8gH+GRJ3MPYqT7Ah+TbYQOb/KTzRtgU49LDR5dyvbv1oPIryitwpU7vC+0HJ
CO9FMYFphuvsPU9nIxow5jAKqlpxWvZJ+GVp/nJwdRiD5jCdC2GXf0bn6Q1uTOmLOH0GQMlpT6Ha
38j7Xu472QtJFjt3Vg4jESLJyiqc4bGuFGNxsMQIMdOobGXjvgb8IYObGUBtfnAP2D1IpyA3lbx1
g82mJ+WNlnoPU8yd8kIOc9mKTGGlwoPcRQ2p75gpK/iHeXGSb9zIsg66ccGDZTMXnYvb17GkKhFg
VQwJ9XnBgabzxqdVDdqLduqpegeVYRrF2svR9AqMyUFA9X6CMmJJXvj1iqFqMc0bNH5B8lKVvkcl
mRn1jmkO2g8vUM9efVGWxEau17hviSznrXjXBnvz/5cUnQKaDMCdajaVvn7VruHs+E+ED+gDj8ZR
30dvwJr1tPECEljQnVQRUl/fejN/lgyfFswIzr3ZTUUDwPIl6un3fTKFCz2qdafJnRmZHzJRoe/R
0M8k3kaQoky710REphAIkAtJhiSwg5q4/zhI1QhvLxxgP8MlGNNO3+vDKWNnc/XBqXSEXaN5sw7E
qsEOc+cbi0QZ1pF9hXV3X6epEHDa8ftLzSXY8ZUsdR51zYcuYHmIrqO85FiowR3S14yz9wlrHkma
rgHCUAJG24NdZAS40JOdyXpt4QUNSdv2jFFoIPUhQA/bjlV3WW55MRkxE+VO3aLl9ZOwCZGFI2x7
MsuG0seDtyFxS3Yba69640yXIqiOyUtOSZrVY0ifGGo4F1JMVAuqfZKnBBPhgBLff8uZM/qjxrWF
oX4S4TLXrxJE/8ClbRD+Jo0B/R4B3t3nMIqG37oZNOczuODijDsUlI2I2arU946ZY4VYGaqKfrCr
vie82VXO4akilacUKcyFmr0skdneOcmcmTVrFDiKkDUVSXjFUyAeWQlie+NIzAexOMHpqvWaKB5L
wOcRcPCuZHhnkKlIDkXsIKZUYLhN8bd/SfzvsAqKmNuMYwyyh7UJi1USZpBtD7YaIydOvHZu7d0T
VxLuAAx8hqtXapZvXHwwMLhTh5ZIl6+46FXWtZkA+i79Lvctcw+9KwoX6fINg1wAx5qKnuiwkY4g
bqqjscMcn9p4OdLMoYNuMwUVMIn77S4wcN43sNezcfb9Pgj603m8sZNTGFyHWaojTev9pOmdqO58
9rAWQodEm3HaixlvRJc2cNKQOGpu2T1NxnrrRrGTrxonabS2hCRcFSDC1vX8GN1S7s5As6qu6Wpy
CZ7b7F3sCU/eIxFqTlETmdjPK0uJXA/iHAQZMHhUVgwWt6/URzD4MrJXf9XiypLdhQUTYztflf59
lz+sHwNqKxS2nIsJ2kFfcIfbv9pjBTNGWVDFo3nRRzbrLVXBirZ1Ywlx6plsaEZGZLUP4p0JHY8q
WWJd1nXHHTNj1+noak6Hj6EbvlgknUcvkTsjYEfWfPupQABl9bsavSW75tWA74zEjXVA/i/ONU4m
GAyDD0HKIWxlzhTXP2sX7hNn3QJ1gkpnQAeB+Ni2UMOT0qAhX8hAP3nAWa9MqjD2J4VwCM3XnQzn
HKhjSaiaWyhKFx7tUHZ8cfzzjPeb5RmlLQ+gF3OOMKm/8BCSZnGZUMAzXbSvZBPJijVMr7CsPQ5a
fx99CQSiN+/0dJIzv8kzBTqwALaINzXJ2enlAkpDZihHj3ft+LI+s41ADe8xi9hiugUHms8obuJD
1LOBec4xF0ff18k7yOp1DMnCyewZY/kijxkfOceJrs2sK9Wxf7ud2N/sivnjF0sNtwpqXhMK8D8T
KWA3RWdNSm/0sUJHbRHuitqLPZZGDOnYK7fI6AJQg1y3nU28x8k1bBBUSoVEm2qmkXz7DXuUUqqL
zZauPoCjQRQ1KOcVaQDJRnmrc6dDSwJ4P0k98SHItjiUVDaOlg88NyuetSSVqCuhReeEGuVR7Yky
B9ivx0gaigY9t2SlLRPaBTbZ1SIgcO55iGv4x95fi0aGzoAH7PHLteRcqGgw9YfFPMYGMPJZgXbQ
7ongl5pnLLxPTmyIu/QAKlzz0PFs7rfWx4pFk5rVCyh7j9Y/UQoI2ul5Veq1Pcx+C0fYTzf913Wy
AuPioP6S1Uz1a8CzD/yrHFGglksfhqT4K/S8li5/HGgSBYkomgIZY6GBHsjsEN/Zm9+ItGSOSnDt
FuoOU1OnGu2kI70qfdaWp5B6rD3Ke3M6Y7HQxE4XNNtNJW3ck5wxtfedundWer0eg9tE7nFxCbE/
EGakLZyt/W3Nav6xrhFD6weaNMN3I7YXCCvrL3S/BECSKhuA/WpYY6qQ5MBR5jCM4nf6DN/or5Ao
OatuSDlNjwsyy6CIyetZhC87+GAS1Z//Ni0HwL5+yNuI+yzumxGrAyri8RyGGfNn61igxEoNSjSX
WkUpaFF3cDYTEba0LSJJIHjuvlhaVxiHznXqMJJZj7yNV532hZmAwXqFYGYxXeebD2Jrft3MfLNs
wbZ1ZQAfR1CiqDgv/Q7V/c9CoKJl+5HnFeII7iAJ6g5CtG4jJu/efjitOxxBDJIbA8gt46vw6jZb
/DdFHcCJnNWe1DjnZErNKm0P4iFCMEsoNwzxQp70EwKT8lLbdg51ykbxeY/SP1KaUi4S4WUyNvJF
CKMaWz4GTnN6pgGqCIX5Zz30L8oGNFwUkt1bbVixprBRojUgbULBEm2pdaHcdANTT4HhTdjhHRH2
iJjY/MrU6JxNHKT6XuVWD4AyZfnRdwEkTfB3sjO2ypNF89ITGOJsH8ZWMqOIXvL82Mip1jEHuyek
NFeQcUD1vAeV61/FKw+Vjv9KoBnBhgSzCNx9Pf3Sm2QQR8PxAzgvVePjLb21rFD2YxwjjHBrljGS
AJ+Q1jD87mo4DA5m6kUA3tORoYkW70EiZH01gXe6k7HYXP1fql8fPiGk/blFPaXVdpkyCcLxtD/e
kd55SYdP4ajJgz3mYfcG1DMgy9HdUeUs0qF+G2p/p1kZ2zFI9UHstP+4MkrhKsi2pbBet8n5+uT6
msn+lCtfw2MaRaB54/gCKzmpjbZGgVoB8V/mgQKKu6ZeD3DAX+JpHtAaKsz2LkE2pTXnVWrm8Bi7
v+unHT0sq64kjJxGNi0fRewaCsl/RhLwmyCnvUyJdsp7YzOThI1YvC4jRzEIWe5uxnadOdmxIzNB
KMv/jpyvezZ2imbh4VYcS+aHL+XnRVhIpTPPqkx+1X6MkPF0imy8Yo2Mq6+q/HigjCwKdmwp7AAh
j5jfZcVREWpCAUhrPkl+puWBm3HwDkIcvOJDx6hc/zkQ94dfDhWoxLY3bddXTe+3jb4ozR1wuiOt
V37H8sAkwCQse+OaU/6kJ47GrWZLb1XmBvuR6FYFzPhVj/orGkh1WwapM++9r1iRlHsRZZRYtinm
AKajMj3EbJgWTxyRuE7QfkxGNGcMy7uEEnLyhzWQSl+7SaP/efZVdfXxhbRdARjnszsDbFIaful+
fTLp/DGrY49JTjeHbKZ0BeIunMqEVEobEtkd5+7RSe3p7oyJ1RSpKqTXbqo83p8Ynk2Em3thRX8g
VxkoKs3S5A69MW3qHG75v8MNCFmwbsynfEgdl46p4GfNQ2V8dZQ4dnrRYNUfpJDz/Y9nuanarjQ5
prVrKJ3bp11p3I2mQn5VzPxMdaHEo6o4pxt9V7zABn6rP1KbAfU7ed0TPWxVol/mVnZj8Omly6zs
I6mDxsholyRSpbLBW7Po/qqCTCUT4T4u/kV5SPUFZFt+4WXilOSh3t0Y3xlGSKcIdvkapmSBsN/n
p0iaMBh+skRsjWf5GSEADbc2pejIlSxO1FFSuuN2cVdMrNBQTiV6fC4OwnHS46Q65sBmNvxUkKOg
uGQRTSUdX03GHytQ8xG6V2OcD0cQ+o4gJV0UT3j/1Tp3rbYpTk14bfE1dNWoaxEAqzvfY4GTWhmr
uaP3hj7pvNpzBRex+yrlxddiOiBcqx44JFQ/dQDwkRNUYgRvfTO14VIyaaxkXAfvEqGuxM4qN5KC
ryQtbkWjUcGpUAlR3zhbpHqIAnysrq79r3hB8qxaXOZ2icPBccVXHVwwfgSZI4K0iRTzMLdRo4Fb
i7qB3SjhokShfxU23xFsHv3IPIQLfOrq+T/Ti/Yyk9juDjedGscvt9vvufBDbw0DQoZLsLWr3TBn
ycSqI3IaA9fho+MxzgJXyuSrWApsrwFSZpJ3WX+isVigyV7InSG/uWy4eRvCCEsEEY9pdptkQhsE
R3T1dSKBDFwLZOZzUmcSnb6YRC93Uqjit8S7bl5YDfsJz9uPtHjXzFYXK4avQZzWpvaDdo7k6QJH
I/5hvVMuLaaj5qzg0ETc4UO8LGdjmdFBvLFZW+lsjniJ+yAXn26dvrMcX0v3qD7dXq58MBim9Mf9
mNZPzJET7MWxHkfGrSM1QC+1G8u6m5TPz+lfpRctPGnW4OrpKeOojzWGvZ6+VjeYaQhNwx2092my
zE271sL1lEleCvgwFOBLcGZUolrKYVndhOuyfbw5DknUcwo3sLSeL09uhCPS51TxpO8pBBUPsJeb
hPea1DCxGQBbThz2KCe0cz9WLUG/R7zWX/dY5gM7vwq5KqJpSdVdF0wehHF46PqBWSWmNqmFiTfB
g3xYZ9y2YLJ5vG1Ea6+KRnaf09U96xBGd9dlLxX6v8IiIs6rW87F+4aMlakEbIgG59C6+oaqRkam
33MRZsyt6AotDACLsBNl0dOh1DjlHcxiz9pwUtxamzVY8MjHoZZw1tUmvdZfmhQPyxBVvi4hfGyo
OpFHWEpw7UDrMjF8XbgTDcCupib55mS2jIb3MMGPzV+pgm6TYIEI1thtKpERcj5GtJr0wpujX8UP
4Fr+kVQ2YEHg7ArcDSLnWuH0tigIkoZAxSlKLMGuMNzTtHvex79HuvmVS1ZJT+3lu3zC5vJBKbGm
JataOqAMSkjcedo1UYrRf9eDTP2iacwr3HHmptX23nAtcPkNMJqZUcVxgad2rEeKvN7weC9H3JoW
HwMQmqV6GlkbvDcdNF2O/qMZMSXRWPRxakFJqOPoUpRCOw50xrdIPapxE25JQcuTyqWvRBKZyH9K
J7xyfl7qucrw9LFIgH1z2uIkSlqC57vVVWU1/IbrbEtvXwjECPcovyIPjem3QfWmpxTrvLzpfVWm
qLRScwIXncMxldVo4g95S0ZwRZJLydqf7dpOp8l7TsLYNRKNW5Jccp5Z3gDXJ5HDKM5hxkySauC+
5je0OYmkICYheHgNFfbDaBXy7PAXHA5ruuzTEkHwWapNqPh4MXKxUfOu5jvEuWikeaRCXBNy+4ej
EeZZDAiibgpNA7+CI4VMq3JbmRpe1RS4XEjz8xrgsKNOU0qNqQCaS7YECXNCqIYpKXAUUHel/KX9
45feVpHvxFFxaFkSVW8TEI58eJBQ49yzGPTNdGMjCLmySYyivpq6rUP6c0KacFD+4UQ1YVI+E6O8
rMPyyemYP3uTpA7Hkir7H5nZG9KvC2UyL4cZy6mHas2EHiPxBfT6KxsnUGzG9L95L1QesdwHpn99
sl605hVA0tB2TdjmGRn0QL3CngtJk0hWcztkzeULXzQug4SYE3rNcgYrpRsuXyZMaCXiA34sNagL
UxyG4FLE7CDn+0ZI6CQSh1g3bRY7Yat/5H6aWV7A0EqmKa72YMwjuJ5Ta8sI14tpBGwwnVkpyaSG
eAFNP05TMlV74jbKhSqZPTmNi8vBVPl3kTnf9QOE/4sff8kJUXi9ev6QGU1gkWeRl+nvllrCZK6P
8NYRHAOgCXi83NnRufi7THV6LLQ+64JLsZm2W7tm/7K34rpjV8PncqNYhFICslXoT3tOZn8/ojwD
bsFcqyNupaVFIeUBysbdS5BX2UO8GjW0oGdhKgHPivKya1x4y272sNRSexxnUKSfG7YImDQ+1/WF
samOadeZsLQUv+vob3GrQjJFkyMbt93CDlpz/XDYJpm/qZQ7Zb2Bvq7vpGnw0b5z9FEFB6dLkAyV
DekxMPgGkpsxMDxtijDzbgDVWU1i3Psmd3VYSNdnRpL8cQMFabu6O7P559nSbrEaAMrz9H9CP3gK
hzkleQiw039uMZ19X8dV9m5/zd+wRmZ228lakVRWUtJbQ9Qs/6NLs0VidRc//UUgyk/lrdnBeyc9
IvI6PBnPgub1PcznVLmsAyILPed0MVBPdt8BMTttC4O2xuHKLZ6L5eNKQdAO5QSkys8vYM6kwTz6
g9otuXV0BekC4ZI/09cgRfPhZu6SGIfQaQiK1T0uMwJG9AHZZL/GJXJyeJ9OQlYaZqEeV/Un3U1r
zq84E9Ad+iSOmKMdngI+RgdkpcsRRY32lsV51gjZEhc8Y6mgd1Uku911bH5P04Ais9+0uLNGUi1O
0eT+86sDaJgTJh4lA4/XLtrt6l0jFqqy7AJTXGbm6EMpBZJ6robptcF0cFk6d5dgbZKKeUtiUJ+Y
40QFE9wBkq0ABG64CHiLtsE6W/dU0SUAPh266tOszzkc66y3KCphduYnt+GO6658Mh1Jnudr2KHI
zd1Tplap/476+fN/FSGSwfaHYFtg00+ABYxWewA5sdydYxGH1THjDZV7IutpVOrMHgmy+lwJ6l32
ELrbWvxCej7phU3js72u03WSWIT3UhrjNhXRtvRfvakUr50X3NfoVXyYpnwnTATEU1Tz9TD5FYz/
Q9zqUFsZhjsimwKuR8R0H5RAvm6gTFBYmN2nsZ3bxwPPvrbjo+xOs2TknLnEs9dgPQk+n514NQbZ
D7khr/oViiz2cw4g8sz+reR4nWniSITVVjLnoA0ruIMP03l3KHq1/ZNfATyGpOGPbHLJR7l2NuIV
kd4PYx9NQEoPmMUsWkVNgMJu1Pqd8Y7PUlulPU3K1bTzdTXMmQffEDfKiTOLjRTmDury1yzqnIiQ
WAdI/JVXLPV/4CE7fR9eW0RJcGGTTptQwOkYiMyjO9sdrSIBsbdhqrz9yO73+AxzYtf3dQexiURb
cHKbET8PEhvEJbyeqwrRt3oFrgpdk/5lbn/PkKo59+zBwT3WGM9XgtAUkOP5Fdxc03cGL8ubHJil
o7bX3C00rvnCLudwQDvBFLSRY08Q/4Q3n2VUkeExuai87qMYIsWsVi21+ogUyox9UfXO7D0baQi5
7pW11bc+9TpbzFYn77got6IYc8z5AQV6hdbR37Msu/pzxwzgYSAdrN3y69HTHvrUBonrp/MAoB0t
SzaHdoXIF1k4btTyjP5P4wIH+RSwERP2DUYKIrASSUX79LxvMmahb2o4xxf4CSTiSsWttZYJRlJl
giPsD3o3VkspS8bIqCIgCudWaiXkxDW6//0lAQreX+DBVVp8INO/iowh4G/s+p50WUsY4hXbFIB7
32y+HP2kGJqnHzAMvGce6EdItzuoPLMX7s7qf0WRXnS7s6wUM5nefJdBXUnfS5b5XYXd2Ip6J9He
6ctDbOQISMEOuatUhq226NeqaO62A4uiYFWRz7Kz4QCWF47oOR4+MtAkYnCvtaFvvh3LqGhThw3T
qdBBhIuaOGTFV8RC0hdI0wT3fiJef6KA+wCHyT7vPSgfzjmVYsMeRJkMLdDotPkifJ26HmdUGNpq
LKWZDV8kahKRzuzrKFDYMFhERizR/GW+iwQKrNBoJqD+gqkMlahWY4QEaGJczaUaiqdsU9+zd8KE
7vuR3OA6hhoLzN2ajqBY22U7fqe4H9wTWghWnDk0OOM6Nh0Z2L9YL98Sd0d1Z1tnVVJLgEzt0pfJ
zAyKLcLv5J1BfeU3qhzkksnPDU2kvemxQhmDkKhfAGzxLskW1dN1YjBXry5V1/DLnW17n33yyAB3
7cx2l205zpwrvPoblFsH6y7/X6WaJWnJ7D4ib3ouK4H7KuxmSq/QVOYt+lLXSj6Cvf5CPCg+wJSU
iA8Tiffk7fC0WtLwDMOV7v16vpfgx1VnoIKKTCIeBeCW7YejzjjITaRc8qt8nr3rHXhZV8vEPh5p
XBhMFNlwRd5jXpbjGRPTOBjfhH5x62aRmyCnCE01bXcU3J0r0pnk1QLfQSC7dMz88tfkAQfvtlCg
X7Co7DphhxbwlkhAMmnwILiyZWJps24mZHIIPlW7525lEFOuwBO1uHSprJ8tiXCdLKa04xV42MtL
1fY3zf1cDHtXWam4SV7VzhcFZpaTbMZ0zPKnxsJsaJphi26QxkUQLuThvwEuXi+LNfw/NdSQ1NFK
4YK/5On3cYUpioTJVPBkLpjIF/T5Sptd6tLYnIfXBtNHPttEe721shX5p7R705kLH5HeaKiAvgo6
nz7hpDsTM92tFS2KRYnalbMnZ8JEQPe1v3Mx9TZsnHDIZUvZW/0XBD7QEsU/ubwH9WX6bh/PCaqQ
14SsKbl8n6WCixnTmtmciL0MsmZm4RtNC1gk8HlImCeR+QqSIwbVGcvfthwylc2ysHUlV33Imm93
AAfY24U5qPY9ONx8RIiiDdP4n893AlN8W42y1rBe+J5Ol9igw59luq8cxaIzge+oyHRu+f5q+0Ac
TFe1aBtsVNMOYZIC0E0SGR8dO/y0JZngtzeQ9fsMFzQvh7Rsx+yM2TPyDkiEZ18MKsKNO7FTeDFn
hoYEBpCFnLyVKZ7mRST+Xv3iGGNt1avwoS6BkpAhUEImQ8hNYphQb9F4SjgsHymMZMsV+WaYJtiv
4qosPm7vkM2tOFbLFeBQVducLI/GRAlGLNQL0eCcxRARZXly3Ixq1di7UEmi/SZ80yaACbRGZljH
E7M75PH1YpmTeYJoY13mRr1Oy4jVu0OUpoQ/b4l0roVRcLGjxw50KqGCB+dVK1s1qmkB6XJh7P1s
We/7fYuTaKiQa+wu1UVhG3WIwGHn6PEXD1/rLz+oaGM10FRXFCN7EAiCM8vQfrEiXUcpjVhIzZiD
H97ySX7JtBhyhW4dXG8BfSrbaK+4nKkpeJzrfvHJHmcxhTIPf1Xpwpv7Gu9i+ZYyu6UzjNcv63EG
n1pFJvecbrcBGB8T4KRVNf+T+i4oxlFRo5vPtfqV7vwmYzlhXVCI+B9Gg8X0uOKxe583QLfM2cKw
NlkUUiWZmuAgCSjkDujkxsUpmaS8oxcWa2aNVlJ2LUeii4Hc+4npbeNFOqOxjYLZyOMy7WN0DBe8
iFtRbwBl8Z9M4UFWBMfuDDCZEMOIWo9W+tD5YMioNJZlrduOskUNnIS/PfpuaxCNPAhGt8Cg0VWW
WQunfXWtOztwDSTYUvz+EJQTqN6RfFD8DxjH9kNtyJBmjOnZ8BTeNO4GqDEioSZVTWH2A1KfKjXb
S7897P0Urakuwm50HkhwAEEtpYaxLnEGAccDIuafXNoTZwCDMjRe32nV2wYktlxSWd7dPJvdFbIm
jBjLZ8ihQejMl0oHnyX5PssIc2+HUxDFnE2DkA+WRKw7A/3aBtZTX7PhITUk52BHmvJtad5ziKfd
YJmkw3B3zMIFx5L2R/qW7E3Ftj92OOStuJwoZBiEpQLS8QBLGhn9yX2FyJBZ34Kyr01GWtZQjVNI
PZ6TuX2W/wM4G9tTRSazEaWNybfOobx3t8by858yMGofBBGWOh4SDYMmrMtQZ/SbyLnK+wZNjGoj
NCZt7gxSLXnoNJirMY3VfrhrgwFFjPh7N/337eguQSqFgMS7f8Gl8JECaZLhIjtcCXKbmwCRfuuE
JYHQUbidH669NZ20LbZn5HUO/tA14Z1LK6fsbPqIKJpAqPM/Q3hFlKzLBL1DDpT+pYFmsedhb/uv
KNtQEhuWTVQu4r86nehhXSI56SZ4FMydTOyj4m+KbUg8xWjLPzSzWNEiqHjrVHRudc0Wcv9Oqs0p
dYT/HJ/CFemo3AtrfsBtGslLype1tXe0e4pBra6mUF3jjOMQbPxqzxLJoz9kAX5r1SHeccFpPqnK
ekgNCe1nwFap4ADHeDMX3c62+W27y4vXXIBJbo5umcJeErACeel+PSkmYn0DBkQU9GeOwqrhW7c9
ZkEao+pPBOr6se7qcEx8WLxXRqwcDmOYDuqOFYSJeSrVq7/PYhiEWZpxZiSIdIOr5juGK/g9n9QN
yO7FJ+914ML+OYmaFKmXcxi8TwEhQkHh1AxXfuEASJsIlvWAa2LelkZqLMyhHvfP4W2hNNr4Fb14
CpnxjJ+4I6XxYPVyd+E+SWHC4RN2XfADb0wkx7mUlKOUjb1a3ve+17zTUn3CCI/CrVzOQmGx1tGX
2lLsxZ1kb+TDmpQeuOgF/4LXHnu69+oww60HaC4czWTW4lK90lwr6PNRegoP10RS6Bv4GkmzNxiF
JivKMIFWD7+huD19pC3gNozTyoasD1pwYrxirlpe9JkYIkLG+0kZyg/TlT+O0TK5ayUd4/Reh3B7
G+cQb/D7888Bq0KfvfqvRP+8QCaBt8tD1Aqlz9ae7zhR+1LmWRs362NMFikec4npRtemKVX3Bgi8
KIwRKu/OViIyVGjwglIfVzo9xSucREgN0ksEe6XbRQ/iPbgAPj1f6BhCA2SCwuqTf0Ohin1EG1Vn
Hka+/CPWVckEoa1oNIzJvNM6XsH7SfvjU+OwBl3gE/b8xk2HjMwRqYuwqNMwgizNAAiDGOsH2cLS
V3sldyi//96fNa00mtkDTA8b1PES6sdXB6uzdDKxMfvk7YJHNBdJzKszWpyc4XdhC0d/rawti+De
b6hZb5D6BYaYedMLt+yWweoLdVD2/w8w4NwntPwWoSckiYlzKshPx7ocoUDBY/4SqE6l7f81dYhf
G76Dxl9HarIHRztE+iCUk1uQ74o+6n7cGVtm8XGnLEewIkRGuK/HqR0WwapOn8mhGVyP9t6RfVpU
yCGBlUzcRj1z9djRIWM24Pi/S4+7cvlcZ0EAV/EtFaQiWuJmB4S6zAagCcAYclUtllAmmBB/ZDh1
Y+v7B0RK8H7CMm51HrTW/rUGveOLxm8hD0Ds6ACimKEB2rvNmAWMr+WdySqJlrFUlWtmGg2hYDzY
ke2ctoPK1jHieqPSwtRLZxlmT/YeK+TvSjGGtSDCPIOqvOTTbH7aPz9dTWd8zrx9+2zhGyKxTHl5
0j75zsZY65oqJ2fYCi2X+4AK2LVBWRwm4Jd6Apb+bNGn/zqxRJj+npBe5LjKZKv6aE3CxQoDXXiL
ZeTo2ws8qWVld1u+VlhfsBSuL4T7lFoCpTDD+TeR3t5UiLxUwO5wC/ww/Ndj28pjPtpKt9/Dzz54
+EsFfFFvNRqBWLiuEan6BZEkqCb1cliCgoyzDlLSfLJJgmPHdJZTQSfX8iUcE+Tx4bd9KfwUiMnz
5CqiEPpn05FVWqw3zTvhKhUsS8hX1QTx33o8siPqQimc6G7X812IhTkmjRtyRDp9oZ13HZs08b3T
+aU+wtYv8IkYlri8CdD0gQU8f+aDgRjhTEV8FgaAg3hDo1WzuD/4EGMsEbpfL3zwKxwGjMN5BNKA
kcuylX09IIY83R590horqwbJjYL4F/cABm5Yo5pE+I9lBt9g9qhg9qxWPMDfmSUumeq85kubU1My
4lGW02ksC5aTsQe64uS2k/7FWWtMp7XChdUaJc2195B7uqiOmeDwvaGzn7N7MrPsWSQsdsqDfLMq
28AOoTRd+ZGrU57wgv7YnkR83bC/Dd+6zAidOoOFIXd3Rhz1Bj76izj1Wtr3rbq0LV68HQNCH/dA
Ws8eLfUyWR6euLfF9X2POrfTg0xizmmP5l6ssTV2bMpBJvmu2+KoWBpEn97pS05NWbS+v0t0+2Dw
K2p1hK+A8pFvCJn3dJGIzOGBG/VI08GGI9Ref0Q2HnleFhDR5maYk6GqiiUrowZ2bYL4NS0tRX69
ka5YDMV8L+MAE+Bp6dqncgJBXdadaDXV08eMleRxKNhOV5LL0KphGIr8jZ/XIx3DQH0aLioOExxc
L6pKLXVirp7QKhUiZ4x5T94HNDAnbl3Jc7zDBNJp6zkqFadayP8Aj5j0OJWnfHkbAhMi4Jg6Is4s
cWBTO87Gi3J+1liRtH46f0B8IVSiQsviMwu0eE80TqpFE6iFVmFVGBxUUqVcR+AdIE6B45oCiWVw
sP5CQy0p0NIyzcRm7UpMWKslXWXLSgZCVPySwdfLFXStrtynsok9D8Jq+xIJavTvjlhuti8eBJye
VjP3vA6AMkCtao7CdZv4nooTljxTIWYk5u7TftZd06wZmdd7o25uxtCOAq574/iIr5W25GwPvWIk
q8lLqARDKJLEvMJaEZI7vgNQvGyXA7/E+OIX4twV+oNg31y9JJsezQ6gwXrrc/cf++AqOZFDrI3P
lb+5zgg57kFo33LtiHPw2iwQLLy9FQ+KI3VLkJATWdScZPV06i8iEayb+Cn915xYdtVF5ZVcCp6D
oSgcjbOgwhJpo7erW1nQWgU3ZTjNyEVGO1kdqydxcYWBapVDIoNXTUSqdjxJP2kDzVSSrLEA8zUy
nSJ4aaYXxtcREnjFyWntkDAD+748IFwgBGE4zOUrujoFQxBmn+0uDgHJe3jGV91FNrjIJAvnZK7R
UQQIp7sCBIMCQmyAAAUStwviqwt+vWrcORiKtL3YfdBDKjZ9AoYJvMSas1rq+QH30G6zn6Pt3peX
IK9UBfV4dc2La1XcaKC/xJixUku/GJmQlxUtBHYECvhyTe4Dsm0iIX2TqzmGUu6TXwHPvlNdwQXM
AxmLQQATqrmfLTeSZvbTvaC2oSZTXSbg4NMoD6EKhZjGTeptHPvmwGtUlQZhXfCrXaDj6aNZE0HO
FKQDgCKmFnBwhEs4CZNwKbDgCULlPssmcy3gs7Ltbns/PcJTSEpldiWXJcFE9fsiA+9WXbmBHaHx
CMTDzZqRRoK/jU1620gyaXdF4WG47OtrTlqZrm6K9Sh9+vfyuZ+Bs7TkQOCMYAAujEnqvFoSIt3+
oHuZkoOKcLuoKNw6C4Rjuu+OmStLIqr6yrSBW7kQ7PfL1B1ZFPhdVHk5kpk0CJR+38b+rYXrt5Ex
Dobn811BPg9Mcja7Vk+bSPqfIcU/nKXE0L41N1xE1kiDg5e/S6K3OmZ770HTuWgFit9JRgSm7iL7
MBlG+QjTiFYI+OUhbXWLBT2ws8WEgg6sZ1vthSuCdqbug0hyv+dRQWodGMHUezwU+4vyqnA2gN7l
frcsLgPqy7ab78mlLUedNZF9a0ZqbQj0gW/OaEbq6o2lz46UTX7q/412BBTGELZbrU6nAqo1vmxT
NRUHchgusR8cF/tmmuYEF63LnhcYG32uimlNIxJ4bd9hZ33+pBp22c91hlHEss4IW9USfLlDza4J
BP/1rrXovzkjHoinSkezCFIfPh7DE6gPCMTiGVepUhr+Fe1D/mrelLldiCS+y0GR7MnGk3bGPqVB
Qqg3xbOMGkaFjHZj6OuSna5OJRxY5P1lRvKBEUAldhwtiW9y8xCZPhSwUxLO+yD/GTnUXOGFWz1S
I6Y4e87GansdAgfAfzEQDEHealpF4VaeT8sTl98qYBRFRi+zA94Q6If+KUXxnhAVIeiL7gix6aQf
RCu8KwK59VXMcHiJy0hus+qXNdtHLPsR5EvYnszp1nhZP1qG5PnlY8GFTamLwX49UFT1VzLkkJgn
XgabXd9C+dmJ3R+ERPuW307WzbJj2MiHxzedckp/pBGpS+om3rxkPrtzkvlVnDnLWSy5c+gCFVyA
deob1/El+tItzLhL+pgM92ZnxVg7mFeIMl8f/IWx/QMTDW64DkIm6T2hkWkPBu2s6Bcv0HVwRAYH
135W8xsxDYoq74fl4fsXMIipxJNuXr+3mwWM1F16gLZLd1ZRLe+H0vc9dog3T3zAl7cauKgcCDgD
rBRKwdk560g7lAV5ozzCAzz6wAvWQuvDacth+wiax6SSCDfE5Bx0IkDzSm5j0fxP8GmmnUjUirAd
rmoo37jChJ1K9JVOOTQcObIPz5CbIJbVP/LDLzYbe/FO+1aX38UPXUtzcE5xCFQfeRm1riRyN8jb
1N0DRok6JhSQG5I4TNXVkL1zDo8mqqEFGahjxVVlu3uP3vuY0qV4kNMI3+NieQunxglj1Gmw/Uwf
5pIY/+sPomYEItKFIcAhy8OMOMO5g6OX+QJ246tm/Wg8D1We1Iayv2h8bleeWDvRB1ZYSC5mn/ls
kP7d+2hbNlKDpW7SbCTppEzyIJeal0LcaKXTtd/o+1rQa22wcsmYG4Na3puOOl4B+odayvWrVfZ6
ynOUdQCNjiNUwOX/Xvx7EAfvw8U+MRnsQvfKe02FC4+ULJtZupJEeHqDIA5wvUR0cNfeuqBbbyQX
3xAz5ugeMzT3y0FDTm1HXVBtOApVgYLrKIiiL1qUSQ/sPfa3ClS5jLqa3azHpkptbBGX/e+ieGAk
OoJGP4NV/NdG7yyuEtEIHRM+WyfyuA6sUFjanZUZiOnzE5Sx8OexUkOp+tx5PcimAE/yFI+h4c6h
zO/z6G4ofadELj75C7tDQXDVGv+4NSBCz4OjoNvO1w45M1njRXbLCgm1IV+HsjDO8dWAmSatayDV
b/C0rbr7j1cykhUts1AnSCC7z4pRVttHvxTG0jmNDocXzyMRuhd0j6jtQwPY7jK0TQY1APSmIMXg
yB18WH/o19E7F5jYz31kp+lSl1BhLbvDQTAsF+vfD41/rXfyoKxf/5NLpcG10ZsjievXkjx3XcdS
hyVo+2673HLSuSpQHEcqWjdRJD8iZDHaABlE4Xsl2oTp+wBksPD79UHBzJLakEeg5Diw+OldLQY9
vh9NW/BA2DN3FCIppjs8CXoRVcUsZQTOudqSKNHzmhLbBKR3Xa+8QKVgIQMl2etG3XEeEpnlgZxo
ZFI6CycTaClMPfQJrKGOU3ZeB9EYNssS9Ghr66JOyDl1GtgMiahrVp3mCxGlkN8A22xPLez/3Q8A
NEHv3SQOYaJFZt+AY7L83ER5K78km2CapiV4DI7DZntdzjjR52xyCGjZI8KUkN1mJ5gIwG42FoOV
GU8e/84LL9qvtlu/lyW2bCeGH+UC2prqYmlL8cKQdyO0OSRW8hGN1MPLWefpjhvT4FxILpVHhDL0
+0vB3+Gp3TjqCY2/tvutdd2Q83ZXbzjBmsye9vhFcLV9+nYq0g+pB6tgPnaYOTfre8FD1OafSmDs
z70YEKqXhIg2REBugqFrU4NfMj28RFhCDVm1rNV9Ymx56t9DkesHyXW3g733oMGtsFVPYTiSVmvn
jAQV5i8vtKDPZMm0Hj5DF4tj30BFQypJIxXvjGxTqM1tuUMgqfpyQ8ZRCr8Tr6KZa828u26afyvg
Q75YMF0UUqtHlAyET2WwqKNIE6u4Hf0MA4SnI90VGJK1vhANCht45ebtfXKWF2HYyL2Cb6LsFJww
yZQ82sy2326d4GP0JMxfUCcYisRw7U+KKCsFr5dkeQr5X/i0x2ddhUH5k2AydUfvvLlAsoslJLNA
aF8BoWLQl+LskRKMbpnWsAhDQpQUxgsjX4PHXVda2TUK1goD5HyRm5eT6UIv6qqX8/LF0JFZqjbf
4WrK7cad6f17IiH1bzwlIVbzxnWgpiACMQtuY4qeKWc+gyyy9NXrcKKkkkraQ0PytAsTLu11bvMI
BUOdcR9aR3A0CbGgprwODsQU5m6R1ZH2NAGAgerMzR0yLqOptpH39+XYKLmgCjWnGTfQNt7HHfF8
fNnjGLiF1x3ngBKyrUSUPhVf+aPPWO1oCpGAlqNAmWhOCbiLZGa1Lr6SLN5iuOk/5B+5BQMyVA4k
z50zGWliGwiAFqjTggxvayifIR6zMYHWJ4d63n/jStw/JJ4ZtL561xGo4mI8e7fj+nynvZK3Oqsa
9mYvnXUKSmk8U6bJXmNhRqQI1H/BmQkRcAbAvTtgSYv75zMJ8SZXa+wpyZI9DsFrsYNe0nkSDkoU
rMBS25LaVQbeR/vpcXRTVnv9nrWwvmMFOb/i49k8BnwaSpTtEecDJkV6VJAzuQFR26OGD897C3vO
8JA41MVz+vWRqrOohE0JCr+17Jueio3+jrvC3y/SVRcUBb/EFUgs0oLP+7VVDByKM/Df3jvQPMTC
PfA/NEav54sV9G8LMaPwXnDZw9wvNqYg2xLXIShB18X0q4TKxZZAbOtidFc+4aVR6QzQKBzE3NE7
f2BE22KsJu//kPv7pJcDZ6cTWKNF+YRZomtu/NjcInb+sNgssM+tTZGPOmaF1OgPf9d2Kr6lexYo
3MX81UNUBd8oF1PBohjwhKypoyev8Yzw4Fdri6AxRdP6xebSALPSAzZbP5FRVS1cfLEfPmYVyPQw
8OYLeqY/OT3bVi/1g7sp6t+aVkF0qCZlqRegN17zUdxQEk3EsFW0RowD3DvhOMv/iPTH9s83aj3C
UWEPnSTwcj0nWIfIwa0KbjudK3LRo8idSUf4edkeWoPlQVOQ1o2AZQF7zmshO3gAPKxc9LMIdEAX
DMwMzpAujl7R91C4NG4s9WNu+Tfzcs01T6/ntrnC4XtMO4cv5iA2ilIhrsGjvitHmsLMPqfO28zT
TtZHST55bC8NrIncoqv9lt8al/+pZ2s1fJGkWxPDH+dHEnAuJFOVuMJknHY1i/f8N1BRcoWEvXlX
pbV6Uc/uOX/EqNLYlvHT+QutSj49rj7YfnV3pS/i4+YPL0vZBCPj0nv5C7pcOD36D4+zmjTdpQW7
sVTKEkbufqtKt/PtyujMWYzOUELZm3gJICYvQPgUQWHRgny0v+K4WEazQ2CwG02LodrpDkbIcuj/
1CFZX40LQjUf0Ct8c3at53Rc39xx1O5OGSLjubURdS1dPRV+mnh+/yM0rhN00SN6Ptzm9UtZKlw5
h1buVoJfCqA5n5/nuQ2ANJssAG0yAmLWx3cT36EgcxPUcOZQFUxynKsrl8igRG3FG0WYugd+x72T
CSFIqqVGBhmNBd0Dajr5pSgi580l9QRoy6xerrageq+A2oJND7/UalZNrrZrNihG3NGj/nFctefp
LnTV658lG6DGuCgfcixUt8nzWxxTXnJeXnxKnpuqQYwyhVyj58RLfrDQ9OHdzjwMqOUARiQYOcpV
I2sjhEFEXSJI192Sny1dR0csJ7Crqew50RIRuD2AAvPLBjtRlD0mgb4XWkzrXJQHDz/ZDENwbubl
Oiz7mlShLhqX15oCeDBHf8sQrAqa6gvfJkR9ZepoYMNpHwZQVj/7rjkpbAG5eaK+6syDDlaHjujl
nFI8gliaTnK5rBWSX7MFSLAgZkyaqGpzDCeCc1IlX9UMvvShE6MUlTIBJEwR6zlweGABTpwt5yIX
a/EWC1tJbI2c6GS8aGKDPhSvYgafC2vUwyT1gpIYshMEET9j2qv4Ypj+LVRoMPmqJ8OuyYCsjBNX
OzozsA/+G4he7WZFOKrFHK8halYsUaYXGdkfBIbW5igpITQKQEPzFeoI9vFDyPjUWJbTUpMD9fcD
YzarAL2PFzzWk/OLpakAPcSPO1OMtwLWFntdBKWyqvI6H0xrt41a+nVdu5v/GwpSg57Es6meZWfd
3ODy9+4bMvfykt05gC7sS6tfs1+W4XyArQ4hnUXtrd+a8N5XY8kk18fUHahhFRdeMIvhH5hQ1pCk
bzjSclGAP9ZDN38nlxhMYl2/81gJSKHT/3ub8ysmbKnEczrrbGotw08yxcfm22FsZaFQZk9g7RBP
fGHuued231fsoUUGzsomBhiQ4Nq1JPoTdNy9qU71KSVX+yU3Ljw5JlCMMIjRa1zt9pg51xT+vG+K
eWeg1cUpwJnbkqKOtLIl9zb3pDgN+l6vwXo5dh+Rio+etdh3wtPr1Oa67bF4OXTE1AUBGhruKCwA
ENt0uFe/GvVRRMRUXN5QZZMZWQwPxRI+OWwyxt7lt1742ALgjWPOgj/hWCz1K/Dj3SS/xFtJNfo4
nB0mTEoDqTbEj66Db3Z5ZkNDDzfwAivo05T5MNshRc9w8U4/fj7Kq9kFd1WRQ5iW0RbM4Vt2UIPd
o1/tas2WoWfYbFAnat4Z39BR5NEP5X3yJdvmGkK1xO7bmgd+7xkBVI6O3fJ/LjPs+Zyxgmf5hd2+
ysUER7d8S5SudHuLVz1tNHuzBcfZR4jWee9Sll4sHTA6QZFXHz/khuazd3NbvSHHGgwc/wQ08ZjM
DH34zGiJK2n5ndct/PfjLhxINwho56MxRBBzOcwk+4nLgQbysJbZGnIUoRizflqe5NPkkttuob+b
G29jJEbRoaaImWAj1kds+4Hl7FRpn497JW3RJKMuV6L0LoQsScOIUgfBOZJ4NexaobEeqJVucFZN
xOB/JHpmldlP1RA1/0ikC8zYFArn0IKwdoqsuI8dhk6SRlccmktuQYbX09AzorZduQHznvR3TIEt
gM7vyS05Wd6qNlyANmUC0FemIeyEIq8JuT+U/f6RKaPiqCxlL0EouTai5QxXKL11JF+cePwzeAjr
JnOwddj2Bve7IeOc9n6Cs8eHnr9oamJdJF4uw9c3exZwyv0RdGarjQy9lU2v2DF0PhMg3Pv+YE2q
XUaQU/zjwlhkCEqBY7wLfmT4/H0L293oWJGhJint8WRmbJX18L63QFKPEVvPqSiKdcLiLTkme+Vh
EVb9spAwe2VeikZv4PY2c2yHI0FNe+m5Yi1fmo592unHYaUGMYtVB/UXIBqYeQTp9z3cIuFLPDcc
S0hKQ83D+0r2Xb+/NbkJ+HDqJeorhlv9U9l1NPa9ylTQbZ6VBjxuUyher6YfQsIuRyiJX3AlkU0R
VJon1UMFJFsDescmTtNYVO2lI2BQuFtYiWnBXJWKmeMkMkfeDaIdkedG53Ldm5viuY6a14RjIgNu
jwMX4ELqufvlilKSxiehIf7IZ2fk9KP99b52W8ZARSB17gJ325yM5pfAoKOLOBCK7ucnEChBg8Up
aYaWvB8wbFoHUvsARmf/ppFbQr9QyG5xWiccrdK77zXYEFf/fZduF/gI3em8Wrf8ob5yd9Kj7CQ7
b8rVmEjj9HloD9+z02J87Jt7RIyIUFmbNQimuEG2DkFps2S9yXL9uIigKO9Yp4fdTtdGaleDLPP1
kH7UglffBwEDBJ81nMfywJl/JAaYGxbgWynlsxfLoayPXpDk62I+Yitoe95uQJnUoyj/70AUV0cU
tW9nH1GgXSO6l8yuzR+eHdHoonQjalr7kfPW0du82RH9+k6T6w1WlobMsR8zz4mf8waq9VRJ4kvF
H5r+5UQEYyx4QMXSE1cy24ufrKO+DvtLXERvkXXWrPoCPZIazvoBqj9/8+BpOM2pvb9ynCMXaZaW
Ah4SRuePkr4cpjRnaE1pYPvrT6YUh28y0JqD/O+XUBKChN+VGwjq7FyANl47/ExAFu6BYX6ZFlSW
MfXO3+8QUE5Xao9O58sbJxbGbVn/BjxytpdAS07lZUy49e3ciawshS9ymlt8ZqlPwBu9Dl7m7TUa
JUq59msFy9G6p5/poaBnVIoptNsJYMJBPNtks7OcYe8XWz97+QbzH2+rVtwyDbPdv5qnKJbJUCV+
jeiwM8AX/6PRJIiD4qt3BQ7taQ7Q+W37THrC9yZrXi8T05GNfbjU2sgiciuMDwCU5/HG+Shnf39h
O3TOsfQUeIdXuGC/rajq03FqDiboMvpidEm5PFHuWbd0eaoPqBinjsoAbIZcepriIi99WbSpKofJ
SJZqZQosVeY8MnuxnYmk30KIifDosoEDzej/v2Uitcb8IAifWFCH6WpdWbbTJ6P1JpTv0/mGWRiI
qkShgKk9PLGInvFfo+aHS2MIggMIkIBtKUxH42FL+OPVX6mHeCjBCHyAAfxHgW9U7fgXN8o+CPO0
cr9f8RKEVLNVjA8rNTWXWSP7OtEwF+4519bJuBdmwoiFrHLilsXn/0DbgdLngN3tmsjWtGCNVcBm
CswxADmgIiqNCSG3E3pHhyLVd0WC71ADWEUDTf7CZU5Qa7YgDxRb+nuLdWXX0GM/ZOmi8pOayVR1
8zxNeEGRONSgp/n6JVqAVOFUwIImsv434zb9gcTfBkp7q6wfu02KZx6Ij7p5MnNvYfPRLBQJNfiB
/H9g6i+tv/bqPOMIPz6p5QTyXrUrWNsiByE8xqIycnBX/rnb42tU3t2qdgtVncgy4WTgtWeDo94e
jWaYNQg8BAWt7TLgQZ+RP+wOUrhu+ZE3P+lGHHnvaJQC7TEjugYv6IOQyk8O8DMyux/4+8VcA4YQ
dBCqlqla9FtuWc+uamKmNo81RM0evzn3QMt9CKX4HYNs7Trlb6diSFXqyJC7L4S9O75p2C4cWvqw
EfGze78LEc1rl7mPR5Uvfd26WuOw3F0r/UkT2ODDlJXo0rD9Z3j4c5O/lHlMJpBssWsyuP81wQjW
FA52pNYNA49a2mMboEhFJKZj0I3lAmQLRmeDcHVVZM3HBFXSMDvK4xFBXG1Sp7W2HbLo5zdyid+u
9elpwr07CgA0V1CU5SNn1fJ+bpqCeFpNXQBPtrWDvxe2ANESym1O03x0TQ+FBQ1IAk+9FxTKMvNS
VWIfB/Ks1dL1luP9d/wERiBmd3gqXdaSVyW9I3PERILAMQVX+lrOr/aRUADFLohuR/ZWe6FpSgk4
OLS6EoJ4Ff8e+4ta+EjDRXUZdhRPeMsYqoebeBef4M6PK9EAWaiGTLC7lMTIFAWJYKZQOuIw6YQu
HDqpxACCLkWBygQwTt16xsgIeCdZ/3eVGpD1Lu2kMZbwO2A6LzzjEbt1E8LI5gGB0Ftj0EIN84In
L60zHg/zt+96IaFbFCCqB6B7Koz3BZVHMCi8fbjtn1xkcf1now/j4qdBNRS7MMQs2165jrMhu6HU
P+vdr55wyudQp71zkHk/UJ3jcCki87GXUR/k3lr+HluRRlXglC78TdEmSMkuxuZD+aR9TQeoFDFd
3j2+dgOohuO4/GPY//DtvAzOZWxbIgfu5K8lp79elhwsgMibB3qS7gZG2BLeZMIkpJsoDnU3roO3
Ktq2L8QVkUiSlJeFWC79QhlW03s2TJiTln/N3mNygl5RZTByDjloOjVlO6gJ7dddLX/b/N0QDJf7
VMHdCuiYvK7jET4NTQo3fK9DarQSI0a2ZrN2q2yO9WslcbtULrXhduKFgI9sGPAJ17vfamVTB51p
xhB7FhDM20v1z7mtE6jx5HjLBnVfY7etq7M/UcG9utArqMZSj71AQGr01yeQFQTF+59p4Zs63eIl
LTA0QtYYep3fj1FpJZjOKcaYcPnyWzOdD9HijJP5Y/qVeKKb3xAD78GwaU22cLKPT5/pMI23Me2A
wja6v32Rt61J+APJS1VpGemzB8J5+XnH4tT0qiz//14bwWuyPZA0Pym981Mca/foIBdDeysuj0Y4
TE1ekKSIQOgbDHA6ok1o9bVuoVWi1PNneG9EKmbqLbGISqqfPUKTNAGlM8bdbh5j5e4xSa40V5lt
ar7r11BquouJ0nhqIYWfm/8YprGKiYthIrkNLqturFLoNRSmRHDvYfICrHfbSEHGJtlcbINhDk6Y
fEcE2DcGIq9zlnglvTcqgPKCEPIpo8ck6bPt5oJV+o5D7yS+Y767VIexe7qbuOiXL+F0hrlHWY6+
nN33CnswhXNjJQCRjYG4Wxxzyt4WWVgC/po9sctSKaUEAB33RbobuzYup7+UiGaUz/iATlpJS7xw
pobUXb9qOhhB9a4pKz7Z5Rqw/VFqqiFtun1Xbd9xLS8Sv2SiHO6EgkuQuVNWN16NSumKzhBl8jl1
VzQlZq8qW5e7vXafO9NqY1v7aEWxVB0owHn4zRylUnUNAd9u/7wrOnE/a+Je+G8pw6/L8e7rij5S
5gxAoSrB/sUFJi1kRUXAhaVMx5Ee9Rql+SrUkQfgcwldAkbwK+jQfXeDxQaIzJfbq/tDvJnuRh8z
HxuulIJpvmlbOBhMh4kPNEvUoVJb5hCDPymKZaHbVUFb/zBQk/vJqWD57SX29jBgDDG2fOKFaEWp
ixVB6TrNo0FARxmzmiazWNlv3uA5MfcVyIrd0WmEbZTSGo2TRi2lscTGE0qS8ff6s+ik6h7xMQ7+
u6zAeTQj3x2eSb50jVWXKF1KxhwzUrlYXnyLAGSp5K9tAhMlj3vNqInz/rQfACpBD416bfo4g0u2
OwiuQr6+5VXL+8C1CPSPIxl7VlouZC56QAMAg6vkeSDV67TxbnRxEjUvdrvFtcisUwkqHvwSEpL4
t2COBTgHTOiwsxugPmRgsU6hxI5wPchle4uqBpUuoy/TWRWbx2w6fds5BfNPBaR6x60BpFmeyXGk
44J6QHqW3ia8WruX9sRJz4hxhH1vV/D/DXsq4ud0IMpt9/v7GB6KgplQ5ScRX12fCVndt/YrrzY1
ll6Qc5od1SLNz5ON5n9I9Dni+uGCSCV66orKLAqvA8FZ303uI/lYDK7peqpJDIziQZ1wlNpY2ilX
ErwqHiduDhr0+qEsLVru2jOBAK7UdF+GhFeDEZyVTWkWEdP1F74PPhWuauV4A4LFslLq/2MyGL4r
O2J6X+psmwoXnLZ4wW7iIexdejT85fneGys8nt+/4l65rNVjD8J2jBoqQQJNRdeefFubJw2ENVtS
iKJl17KJrQrp1tKO++9ZCVFC2lK4mmMytrC58/jUYolMGd7K/2FRGdtCaPid7XthGSyXJnHa6VFy
drqXlw1/Bjf2E9h6fWQ4SbjKSjNU5ryJ2bcqfszMEd7+E2+Bcj5kt+b1sF+9idcA1zFkS4NtyKwO
IXvcygDaCh3wfuavX9RDRckcmeOUCF5FX4Pyxb18nsBFohlJmLJnY8Uq9sgeY05h/fHy6637ZTJ0
s2yxMHx6hteF5pvf5/gs/hvEWckv5Dts9MGZzhtPYooJ8FCT4jYLiJ6TSxjfFP9/4ZJekGDF0Rgz
NopKbvn/OA4ih6SPCYD7orFKgx1ssnqVXomBbs3juBVrsgLvDmqaV3w+bekZPBKWeq1lY+6Buod1
Ie0ff1MBs2c7BWnWYJBJB27VBNVwhqLFP9cQI2/VQCmtEniByIWjTGzAjurziOqd/BgF+BAw3Kww
u7QbUqzG4yRjPiTp1B6BVERSZEmCWx69EB9dlDIqF7fOPb4n8CncoduK2c8MLyzpofs/7fI6kBBW
5lujhqSyvydGeewe1IOgha63klepphKxrkpxzAjMnwEx5PbTu2jMgOX+S5SY6YrFjWiYWwXAoL7u
Dgn0YmEFzvVnAcDaaSgtTLl6gYt4P0GHJ8UckBRo4y5V7+pv13lFW5wUyB/zzriPLBiDR3tRuzuJ
xteN9ys/WIt77DplGpO22Qri+LHXZSB939BK9oL5Ux+DVVGjVIRtataxUFYb97dT5/cn45yzvcIU
kKhtIhTdw0AjbZU5VDlKqijOaY6X65aISLk9XtVZ9s/yr6iFtfi2Kx/rYeo59tCcwlwZCjdn5aM8
pdeQ3WuHZ9qu9Ysknp00Kw6swFiqTKToeQ7KvT+ne6GAZY27KBqLCtZbupuIkp2ihPc95LI615GA
hL32BXQ8odPVY25pK3g0hykxomv2XWoTI2UcPqtnv6WHsC1rzWrO0IkYoJSxIzmkM3jRDTW+nGhK
40mnoPaiFDgVDTRcZjZTOJLS+hsoI9i+KM4BClsCGUM9MeX9e6tu8lTU5V9doCwwMe+5VF1gyx/l
D01f2ZsNNQoihI3iXrSTcrnbMHWGepWje8okszx9ZHA1UNIfqMgmwmHdUrCCWb3uriEBiGfGRR7v
zcY12f3gbZ5q8mQnKVjPAExls21uubakvt5mZ6Ya4M0ZYxoWaVCcxlg9mqvTRRWFEs4+C3YKkJLh
TGjIFlvo6zjn6ygo2hJfQA3deSM1CUqNEV4jwfK9TOQsPIMteuFL8+cqWECLD2N2r468adUFO/nT
nQHBIrCEj+e8+JSYCOmw+Ss0YrAaN0+8jqrjQ/Y/KpzlQc9B8wIsIpRnVjVuG1vP+n3zsFSGgiwv
0XPvb7vSiydu+oSrnZoy73+JgGI1rVotx2txLFATZL0O5cGm9CfLOw1P9s/d2+NThdbFxasf67Jk
swmzjhvwcAdFBoJEsFr6Q58Yo0mfwpBLQ7rJS0Q07taMQmmBCaVTU/OsFUpxTf7Tj50dsV+01wOM
0P2E0Ai/eIhnA+snr5dg2hmeVJ0FFMQJyb1gO/0ng7+Gtyj8TY9ZM30URVvOEn1MMEJDOcyj8KGU
2lZwVubKn69wPmgZF9Iq5ClISFVf85hofQ87UxylYkRrvl4FzoUj2H5yMWf7uOOiUbcP6g+ZaBUk
rqiBmjOQy6UcedWc8mJOjiNzzDrtGjyW6oc19kNteP4US2rcyUUdikcFc7quzZmm1BMRhfzONcwo
VBrdWBLj3J6/rqGxxTe8EznrRrIuGMhgdCSgZF+OAA/JW27gVJaeF6wuq/thloH90KdcVf4ww2eE
Q5zJgSfBHXDSuM3TlFE/OYloj2wI2y05Vncnn3Yrg+xWLWQskPKCRMJGHzfbD5RaQO4W7cE0ZgSQ
13k2AbF5pBKjoiV28H5oHPC5209+uIYjDs7CKq0cUv4P9Eu8Z+KJ5Z+3GG0nmZ1XII25YdsmgfOx
Q8BT6wU0BhCV/yKTbdZta3pOZ7BIDyRAwo6EO1LRS4aR3jNI7+AYoytIPaLgXqM4HPOFxNvfd0JX
9FkuJD5Mb2SBl4ONuENRn+X4UWXZrqLBpaUh1i/p+No8xUG74WejOHVUg30zmFTCvL7rFBIhYkWC
jMDMpaEzfa/EEK7vNAKW5fSwWnLJCDYHZufyZ+lfdEbfTtWEePMICLKiJ6oBtM9qMPPL7jwkMsUC
HEna1Ea27LE+7+8QIl2GZNWqogCRgLpb0giC6vHCwUsYHOfpJ7Ao3K9y6rGLSk2JUB/FSvXWykpz
I97JIrqwQ+CRzObfodS4exoXOy/JqFBUvwwv0bc1yj5j9XFk3GSMEYMQO1ily+Mf1nXoqn4NXTHw
qKzI2qkcUaWTkr1aCoopRMGvevoFJcMoL+RnvHpG/t0NcG1TgFG6GoSHiaHiMX6r1I0zWaK3S9Y7
BfrDUWME7eh2gp5QwC/eFKqX8663jB3UNY8p5nrgUhQkacPGmWzQ13JTNTNEKOVoVsKVwYv97hTq
C2M+9+U2QXyPvko6tKZmFEj6Epkh6zbDLTP9onfVOXOjdHa5gqoukBk15v28M2KwKhHcU7PTV9v3
0VYw3tukoduuYsuR3BokCkDqgMkMx9+an1GbDTzuzr/xC95JsgwrfDEz/5VZ3F31n3QEMwZlj3SP
3kaO18YDCD91debQZc2VVupKnEyFBNB7ISDNYCAlBFNmwLfbdOtUHNmpR4FEPBLpw0Xr6zvY7mve
TBRLz9Fb6NQ+l1QtwieK9mzYayvkmpilzvwet6NwXsnp9rZ7EduI/Oo9EBl3+T1fLPPKYGcPsyEe
rsf69xsC8kqhoAOoz7PuI6Lrg2hGyC77hQXjDtsLN/lUCoBSm/1JuESM/uxzWulKlCnQ8Qg+85sd
glxSw9MEQ1u9aQnjdgxzXge972na8Wp/4/6Mhp4rW0lNO74siCpYxcJXLKhp0DA3vn15/yYpCFJf
86FNB4S9tK65Onw5xCfC/DgpiUNKDkiyTNwOfqXsei5B14NknYdASDBVz/tUo5qvsmP6HeNeEwfM
pAPTDHglAUcZJB5tuENEVVvgznVOVs/Cd5OW7LPyrH35MrjDC5GEuGpNVF5e1gVb57Q2zokD+ERQ
h+AYNPornS/mAkzFZyJgbkm8hQPJHJG1/UoVIhqDu+lqohGLFGVDu/fPzDDpJf1irLlgNsbzjUVs
X/sZq0eamo5BbHwLEjE1awagO9XpuZ5fCQmy37IEZSkySSkbFnAeeeQ/lN74Tpfxu1YeNot/EV7n
IW7ON0tU+wlZXCP7IS89XXCwxrGW8PtKOIRh5YjW01Hm87NPR4hJ2WccMbaYE3lfP5dv7nWb6byM
AWq7Jm/u/1T/uiWQzR1M4ORCMes1aweyLRJrF2jv9H8NUS1F1bwdOQhKZUjejLU3UbCCUNavK8pX
Vqj8rSTfWRaOdtO8OcE/bgYdAATAzSi3VviCUY+nj0lLCjscsjMZhwiDl2ODOkxgI28QVH0mgrNn
mwQSRHqsbE33/r3FJMdmcghgIOwntW8skfdybeUfwgxHmRKRi61gJSExI9nSeIuQzrXPbUx0VjL6
7Z1Fl4wAYPVLowtbWUbGlqTZafSq4um2bxWjFSlvtQGkqMMX7ZEeWfD/k8sqFCH7pbfnspKpbIys
bZXA1GqUhQqK6HtsOFFtHdSxIdxkl6wVxEvpXBY1CU2T4ANb9+02VUvjp62N8pKsMgASYHUuRaMf
SP2CtvXFtGG/O9VlCIsUN3hRuQFjx0BKBQSDinDE2g4V6iKm7V0Dv9Vv5td6EfL98amZ9be8LPHI
ucIg1Qp14wza9omvy+rM8GKDEXlp8dN3/ZTslAShhbe1V6p6JyWDLVI8ryf+Bd0a6Rj369nZzLsn
MOX0snr9x9JJaBzfPdYIJkcbMXMqT4B7JlNQ6FzFMjhb/ymDW+3dqKwYEIqSLS/2uY0TgMe+EeIe
2HzWW+WFXsCGXwH6VggwA4GDsx+in6dmP6N/n9ZosLmU2W7wFJtDUY7GyHuYnGpRgyFw0G47la5J
TLFyu7UGQvxq+1AFVUbH3PoJ5eFFyAh4XG9EQ8cEPFfKtLbtucsvUtXykTVJaCzTKcn6EzzCIPhs
kp8QVIc34KuUZu8Qdy//CP38i/7R7c6NBgszR8HdP5lZVIP/56ENylFFdAwA5P/k45/9Bas2QqNM
YlZsj5RrXWOgy58llRFd1HxggD17z05QZP498lAIKbuWS2EqgiyHVlzvm/sX+0Bsg/Y9tTULVRmt
R0hsFs/T7nroBaDZCqvlWG9P3bqfP47z72BsxjcSXUkv3XbIgvrPQjT6XcayLLTjLseatOjfplh2
89qA2aN/sXo/SOD/b45L2qXQkPQtd3W8/AF6YhI84UD41pUfFJ9L9cvW1TkEoXDNBigcFT06Ro06
BUp2xnrPNSPx/PBAHuqCi4vBdZkuBHT+Uf4Ct4h8eaibs3E0J8JV2l8P+cSvfBzyXEQOALnrZ8Ts
PRHJHrop43csf9MVQ95/FgGFoR+RLhx9CqRHNg33VNj2GOvrSEpO4T4GmysKvjBVzcKHPVS9v7np
tK2Qy+eroMenpGm9kbN+LLYJcKmxurKOYLgFYv8sPxFAJIgQC8bg6fLfAMd4qhiSEkgcN9xlwOr/
lttExjyeqadcgJd8PXPXNnrGavtJKxbYRUJl3Lxky0xtCqZS/wZwDkv1S6YZpQPVoZrWDGeiaD3g
0q3WwLnk7fH8XWFI//DIbSw6qF8fa5JTo9ntlDb8d/1FX8HBgAuVaMeMrirdrGpZAmMD1QX6rTAY
gpPqQPsC3p/++bVPj/ZbgMkQ2OlROcgBFZAz15ZGkOv5XXmGtabVwwY5GVOMibGWyiGnVJPWyLf/
Y+ah9iXToIHS+/M3XoxLOZctC0mewe5p7nqg99mIx5SqzBu5jYyjs4u4YwAJpa/EABES9cb2FbG5
B+BA4LZdhT68yoMRiEgaHF0sgFSdWYdEth3PzzZUh42F7Yb0VTpnYBfPgx3xRHjj1vjPkdT1Ifs5
zGRhQuZZxiSHdNDFqCMTs5zWGkgwIu8o9IEOdQB5kpOxBsNTDAAfEWQdznO8ePWdG0JJYrUsOf+l
G4snf4nAVAStNuV54JKZOv8p9VaWqIo/PyPMUCnAePcFQWPzFdPwIqIc4UsDB8oeugGlB/7cCMpK
0KwSiF5297PvmHFkFzCXYF7o1tlD910NZ1oj4meknQex531ODE2H8kr3DthmcyImRBYB2Z/e0tIW
gbKZ3BC+/L5qj/Sx1bhuhRgRguuDmNRB9WsLkGqH/EPpVH9RB8V1u+u5w7onHxWVbQv7MtvtPREP
1zXrGPaU7yUIhJSyGaLlnT2q9pECSTy+lmoHZi3EbepK0hztkOUVifZmXMPS90WzO0YLZMH/lnKZ
mdOysWzQZoJl4+/9a1fr3Pa++bId/zStRBg4EzGWoJp+d45MRBK88UPVTcZ34qdbjIEdvE6hJ/Qk
2vMLn4tHD9BylkMY7It+ox238VURJor+Hw+bEdt1yPQb/NIgwtjil9Ak9rfzqBDfOmFCc46uBMaq
7dWtdrRpAA1AqwZEZmyLCy88SjF09c/THN/MyTLoW/JSzuZuO62dSWbvWj8ljBVbJA+VW4pHvGHA
6NmCH/OjsYTDoAgDOH3GA7qFd6kgA8+LoQdJIh9VsKh3lF3OXGumQC13whEcu31Z50evjAU3nuJm
VJyzSA7MqQfRtOwVLzzqgAC9wcT88LrSnwRhwXxRswZv6WXJg9g9TlbA4kymlR0wZDn3GawyUIwK
Mkj3oTT329pMV2y0cX7E0kekNujrSxOXkPFAcPB59SYXTYqQ/bSN/fniGI7ld4CbcuLvW//C95Nv
n1qcvDgqd6kzEllicRSI5qAcGCgYfHJjXZocJ25n+Z260WJfBV78c0e1zCCfW7qvR6zfXnSRN6Pz
8C9yhm9wAUe7bmKJSqJYb/A0HUSQ5OA60r9jvNNheT3j1tOtOvq+0/ExBaVqtlQzCAomjgNX/Rwy
VG6L5QCOJscyjLSL+TeABW4OsQR9ijanarmL3p5u4H76xF/2qjbNyKzVy+oQ/JcanjbKyej95SEr
9L6mqYmYYxzrTyNdBUXaxSNnvfCZ23xujUBzdlHvsnwWhmPgbBhxnQgtgo2mStZiy14rihCQB91B
ehi6Jrn7q+TPunu4l9p8EnQBZYOFcGnW2iv6wtRYaq9O3/AEK10p4bqH9XZIYanzALpDFCIYb6Sy
o7WDd2KGoC6oQjYt1WAYoeZplZGgS6LGH43AqNRsJ0DwuegK9FRpRpqM3nIMmW4DxOOoHkMuYTgs
bFPU9rqg5Z56c5PUYzXz6hIRvGR+qBRndICIjqiAYyZuafrRxyayjOpILc88bhVOicviHfYV7ID/
X34qWMQbb63Ojm++phWmWqP2TeqmhiqN111NX/P6hF5FVnEf0nXKmdLicKg/L38Ce5cyXMLiIzqo
YRmYelfe6OyYNRiLr5WCeAZj8GzIxiMfc/qWHkWhJWCUn2JOP/3yqURncsZTMZsJ+M1m4qugExNJ
iYTJuFSbRXl4/N+fSRNr1DqcXXKjnnvo6kL5YraeYJf/GNWDWqa2/I6rgyAShog1W/xb3VwWZdIN
QVE2h0TeTp5RIEK0qa4RDgEC0p96sgNiqT+tMY0ZJlePxEqIBebzp/+NaUZ9jt2rhZQxh45+AJ9r
Xq1yIlfcYh9bN459m1KsfvOv8qb4LeAVu5KuTRRUkwiCQEP8rar0VIBtz32/vyzYCSId7neocgOX
w8M0badFIDSMwD5V4hri/lkjgciScKrw5y7h4svveNMI/JcbYlXRk4ZPyVdcldnfafsypXOx98Kn
A73vHKRIHIler63B+ZVgMBIeIMtngDuzBCv9znqSMHQaCeuKPaXqZve3/0jQqIG33sIh6wcid9MH
53WwnfGii2JbnP4Mi4DRDkC6evQMcte9ViE3Eq6q/dAZvnJmCSWHoPtwILH5wxfJduW+/9z6Ggoq
LMT/Cs4uT8Ntcu93mBxAz1IP+pfEDyS4Qw0qe6dGQAlEANiQdXunnA2qNjxefWLlZ6LoBW3F0kMK
/2miVTU2fpZmxaSkkbcPXWvayax+DDWMghW5pcrdjN4ul7TvER5DpOe7oCXf7S5SO/ycMdN700yA
z2ivew5nfZJBqzmPTbyyeE75O12qvwgsm0NOxduri7t5JBNDV/QPIn1aP9lac0XGkj39fj6tOcUG
HpNoEY5Fjy6rqCH3uFtffCdLW3+kn3gzHRtnXB1bDDiB8Lf/bd9M1Oedgq0jCxZo8OfMmRES7FFY
tGfactfDeHzfsZPLkuLvToBQddotwddPdOVOslzmbENR0tkcqAygWQp9rG2cW/tGjsQZiQjecbU/
UqSCZU4t2+ilnuJXX/W+9TeCepRop8pxBQ3kmjXMu2NErcdMWgzv0XeJ4NiuQB+poLElrY0Y1ioS
l9NlOcSpFbpG6xiXQL01cXUSdLKYfrJ59eFGZzq2PNA4yUUydJ7285UxI8lgq1Ut3foKJ2mz+EXz
WJwqZaq2YvPxi/1FNGq7cdZHQf7qwM36Sq03pEn2LobWvrhhGOR6fJLB1/hmywZkzZ02uYkpyue9
DdGeqJVur6makjPBePqxvwF20WuSPaGXKmQyKnGkuEIg60AaaE7iuJlVOquYa1LT7I48TjFcNl46
bBHsKkreOe0enilbtf3QZgaxnQMvNOYfFEx8yXDfVCWo8wP7qXvotn4VvavwLWQcM0XRw1mlRLq0
No7+2EfTWamWJAytc94SOB58uHDFbiylV2CQI+DUULme6+meza5uISGC7L4gG3Tnlbcew/sqWJAa
eeaXMpAGRRucnNpwcoU4+bRTnBHaGwo7wSlRW9kX5xVWmCy03No0pLuFo7dtVipLtKuSGEQZZoSW
omUEjLBOwr0W2RHcDHKMTKNr8HOAiZa4Lk/jSt35knvsKzCuD4Suso21gJGopA/ISU41CGup9Z0T
C2kiXc1Ki7mZVOWXZJTqqyy7ccoUG4gmdxBGMYJr67zu52KeAORRo/O2YJR12ka0VsKm300zhSUI
0wjHBnM+KqDayPzupLdV5NHVnX3TEn2MELygTV2Nup3zGgSdC/czX9iC5xpZR6Oj8rnWVtGxGwYT
3drVzl/yOIuJ2JPGZTx+eCnNs3Km/rSBXxR5e9RFdabCNdJNBYyWW/xVc7Rq+3e4TDG8Iu5Dw9bl
p3NIiTARZqVRYZMx4DxG1D/ii/w7f3N0gHWSQvP4o/ZLcIeCWOo8+TX7y36GnEtevLB0MPw+5sVp
QE6gJnWYIVltz3tbKVS/JBM4/Hk209cvFV972UsVCvUPNf2hZZnAus/HZ9gXpcvDVMFzaHZOuM29
LkeAAoCYva0ydzShOS7bA8FgIHqMP43rIVCQogXIRTvbJFOh0WGVMaMVrMT18PmHezZLIW4xC1FY
aWoDpX5hu2/qM0MhSOlHgRYcVlO6HBapLR/Ytq+YquiSv5zqgD7EJAohuGzME69YoYac9+woSLSA
CgF/6X54n1jCTaKZfpKwhRp0/g3aRRnJTsdm8tJfqw5xOuTsju0QnDfQf4wNURhup33FYGVInvPo
/Y+xZSVg60hYGIRBD7lUZCcxO1wKjgZpxmx6v0OOR9hx4j/Z+uYbcL2ZTqe4AKLaiXXkcOB8CHJe
fxKOFnsF9QxcP/jugl629xXzPQf46YFCmSsoO0kDjpuzLkC5REa0xbHjIjVecFnVqtNYf+qA4tqy
sCMr3ZuV3tzMQMteq47tj04IcbjjnxgAV1mjsmNOACRWgOkahMpPnlfQLg04qDVI/f49bayye1cS
CxzBp6tm/7hBEs5oIubChskaC/PPgDSd5CDdtx03C0jz0f9PdIA7bJHplcSIuYY0vLJTiZxp6PXM
F4ToUrZdPbsVq9msuP0EvIXi4hxCvZhE2EO1/UW2GWBwhEbuXCqLRXyDHkrRV2WRXqrajb3jqQ6P
bkGtjmAdK1pcSkwhEwdPrEEJPucI+5253f+wkJkXIOPdES3idy7/+V9GPWifjqA5X94UehDTROpC
9/sSBJjtJAQGMk6gDR5N64N+EnvyZI0aXrRv+pO1u7MoA9QYvJqBD3XuePDLlH/jwT7OjYb+dFPU
zyih9lJEcv5017K3EqUQDZ2xZyMtEIV+TRzIUDQ9YWoKFJV4dHSZoxaaVHG8Ya03ZdMdnAXEp54e
37d1SBo6WVGjGrP9s5AB/JSlp4b64gKqLBLe9x13SVQ+8RVT6/kh8EUA7gCDrrV04Xw66nr90H6N
DfPIRBdyQeKpTb0m+vN/XiTUVoaW9OWDteC8s3K1YslOgGmnazPQlmjOlfBKp8fw0OtWHVYXbgP9
lN6DpnSAmlKLTwPPUpwz5zwBbWX3mfLTBMZfe3wopo/eFhAecNNOMIvgTMydoPP6FED6zPaHG/+e
0LHoskJ4W/aN6hbTpWE1L1SvY0v/4Uav3Lg4IlJO8NdWSt3/B6uinWo0fKUla/w2OWx+HE88bpT+
lqtr+g/wC3mue2TKDBDIwaDuFuD4JUTxZKcmr4SgyL0Cru/jo2OJ2Rol58XWqiULAkac4H9NT8X7
/lXygLxB3K21n7w+R42UZe6fNPYidCW9NfDtC/SokmWbn6IC7HlaOaIo0PJHoGwcaxgo7jSxD0Gm
c1L1vUNwxx8aRvg+6CCBrg0IjY3/j04/vYxKaU//9oC618zoQ7Av6xIhRj9OTJ8KXSDIrA69gIW9
E/j4BG4aj1MrO9eIXqnHLv92RAYTuLmiqmyz877Ogxzb1zPms7Ltil8JaBMbWUJcZppCdg3Fo7WN
X32u3Z8WsCVkn0DGs0J2gScy60W9GlSKCWEt45xEEzgwXlx3SYC3RPqGxa8zAkIePNeWB41RXw4y
O+ucVnnFmWlODmCPyHtnCUL3TsweGDNFW59MvTq9c/zUkUqvtT1xdiYBDiuL06WhwfZAqixHJgK8
TzFj8sawOetzaWRZdinCDSBEQYX2eSTXCmoY8Dw76PJgnKl59TwWAHQzb3a/kOTurwsSBu8X7WJ8
FUuRoh+YagB2ELFEnU4vVwBOThVqd0v5jCmhK9O6/bzPJu7/1wAxx2l/Yyd6Dk/Q5riOoXQnLhqP
oheqBe8f4nsGQEOj7Cz50I17rzm7V6OhsR38GdOCtA9aJ/i+EGgk5m/z3dqDF0gjH3Z7mmLE0dAJ
swSr1DSyMIUTAtDW1Q6Hy1wSLJ7W9MulVG4i8oJFULHtOCjL2cbUF0/u4IqdTJjIxlPzqVse/Gvo
AT8TmFF1ubYcCrsTNaVeIsZg0WRwnxrglAE3FG+OKez2Sq7ugUVFnweY6iIEKJIGU2l5jkbcpJ8s
Ch0nEB2fHqATsZppM/1+cIfD6Uf61A9fwnLztPHhoAuIiJehhzX9pH3R5P8vsDkfN9E2fysLQ1BZ
Gu/1GUegJmbsBml+1wEaWTrKIQwCftIz8/LXHPxbnw0h4cQ33ouTr5SgWwK904JppDdq6Q+BwYoj
YlzwdSBsQcTN0fhIgGnyNJhLQc3hSnbcwS8JtaIqCiILitv76KpFcmJTjTWGsVlqvj5Ld9jCgWE1
ZTwE9eE08FayppfNP8p3uTLqiU9wu2ln574T2EbYHmP+MSlmD1ch6XIO2jlPKhDflbaRPCr+39/a
OH7nEY6B/eugu6gz2JVnekbHKKsjO+5/Bd4rBACjsvqlcRYHqsEaJEZDw1g8cXpM45jEbQqqUS4m
mM3kNMUol6Xb7XdZjYIvUmQ4tARAzHsbSNWeUuDVjbXBzPCt8LSVQQLO99DOjBSQxmIGQ/XkNf0o
y3rMN4rFAE3ksMDDvxqyFXF90t6madsfnmeB/fQOr9ZaNJpET5ef40c6yYW3EwVzgqyuhhzwIg13
A7C7W1zEe4qDHOC3IiN6Ni6Lx1O6wQ74f+0l0JQbOtwFkN1SXP8vcjpPqch4YKsrGVucx9PJL96h
B1kdX4hmkQyjUnv4Ko/QDwBNrA0Pt7gAFxDrfEuWd98NymwQN28BDuaf2MH2kzyl4qbNEBdWWjie
0u32S7A61GPjjnrt1sf1jfAOexwaR9EeRGtH8uiqNsMzwEvAfIYaoCHqPE0gPxEnm5wAAQOkAKYX
sgoKXeHz8hTDMQ4tHxzyEL18RwP/QEJLxOAf4PEClSFcPirKCtdUGBAp++FJDFmOqxkwV8n9MbUu
+BYG6TP0ioXhDgigj6DEvK/KeOPZnQ0Lhh/GNFzG9bJZZQHV9O788tno0yjyD0/m+sdmX/M35X4j
8H2QEaVX5r4UO3L2u4WfQsznDUP58CNdX20BjaX7F0NOOGNN+vwbWCtZRLc+CBBdjySguMKisDPe
/LB84mGZpKQmtx7IxWQ6SFKWNla+Vujl2N+jNYtEWXYbc92UYUUuTGIWquGBIslpLOp7YycWJkkx
KmwunkyJmGep8wHTJuCkWt0JEEeFIwzxAPkYnBoZSEdat/Swg+JUwMlrO3BymuV/qxXfTlWuVlo5
dQ52APU7nOgwkj86Akj3qjBWqNhQGXiZfmGIQC4qml6I9zYXJiaOrnV343O9SoO+zDNpiuYX7A3s
RQSEZQ32AXyzAz2k+mJVu0grPPElKixtc6MrdpJ6QxU8kk7svzgwApVRA30jsq0xvqrOa6maAqbm
aXLh6en1F+Xn7wlzYrRRp2xR7RnkbdyZQ+wdHdBssfrRDHa3wHf2tHguKQAjTL7aRxNjPhCROiGO
7C+7zinxIfxpjeLBNEJnidYCriUsZw5TdCeKkrGttV5KsFDuntq+nn2Z5bvkxlRCXAi+FF6rj6pe
gDrIcjcmuC9TO3dHZX4vFCQx28lO2aR9YSy/H3eWlO7SVebiwTgpGp02OHxYUuqpRd3ZkoyitmTP
d1MVd44AlWVyQhg3XNm+ZmQiqBHM9000fV839YSkFaCaKPJCNwbQb0kJu9tqTbH63GkqwuOm8jDW
UI2aVdT3Pd9R58xgIToOusixOVBjov+hsDlae1T6bQgQQTrFxLnV/dJBunZkhSNx4tVluQgMdeYw
3vzZUHgSmfEsST6XJqsHQg6VHhPG8DEGsYMNKgxVXRraLagDo5hCSHqBCWa073KKZFaAQbFASVQF
xWeDLZ6iUkWMKxFyiKSzh8t1NKYnaPQP5tmke7vGVVXzM0q+X7UyAIIy4nkgFwQ3/77AKXGRX+K5
+ywXV7qP7Zf150b8LN+4tu/DHnnyWCNggN3XK1+R00yds/5/eM4YCNiFMINflbdB3pFCnCrYhNnG
f2U4QU52jNYwHeqlQ36TSmWNqqzHqyIVdMdR5QVL4zH4V86diflxxH4ute8qtKQY2HKnnG1Oa8FY
+CL4tJntYgUhYrOu6EhbJ9WXMaLUR+nugwp/mW7wfjUPchO0sdwvJfDB7l0WOU7J8xVbduNgpxmC
6I9iME3cjBoxpU+eWb9S/4MBPezW5TvdGSlua4GAQ/lDU4CL8dMfxnxcdXTka+/2ExLTrjyacP2a
PdUH8POk4uZqejOdulfsq2HCy6cnJl5diLHsFtNjNnpW3LSHmWZci46iQE4IEq1wLcKwjr+9vbtp
FFwiSj24utnyHx/CPBj4wSSBHHybX4qa//no9IXwGM9Q3fAQaAU7m9/0266WJQz+x1L6P0QTS1jA
zaetYiljO0x4nHTpZiW3Z7MsaU7HmVVPO80JzFxh+UhtgGrUsjtvBymZP9FJqaFJ4L55yNyZA5/4
sBETeXz2RimbjbA7hzfsbVXbBBfsFqq2q4vGym+qkIlmDUhg28veKwd3+I/l4QXUgEH100YXuydC
TkmZcJSbgdqLk3ypkI4gpr76RAQO9NjaX6z3fOFzotbeiqMe7ZN9JZLnNXiWB18GRnD/zcpfPUtp
ttjazVp/Pv/UlRaALfZeJh46wUaSR8hPBtOz8PvWCAa3T1R5SV67Cy+xX7jMrwdqjth+BatGZ8sU
aznJty3RHYF5ukxvgAI4R//yYxv2+RIRDhb1ATolcEm9oZnKRAY4axn+6siAW7vHOgA0mMlJibOU
G6jkfJZZyZVpgCxzDA99AZCHqk7k89b5tBdv/0yU3Zuhgj3G13XVRZGalbIJzQN1l7/zNcbsF+B7
lrd8EDSKHfL6TYlHALKPJOTfcf2JY4uoFZ1C/wJNEKjPqP/evmhznV0kH9Ex1msZ85ES08BGpEPG
Ehp333aWAJlQIVynNHzWuF+aMkQIWSKkEkf1HsMULUh7zwaKncc8FKRlPqDGrIiHNloiJa0ITtrk
Emk4HhPAcKPfCCi/Z1Tqk8SoG/7+BFVvhhZtzvl5I+EFa7OjlAXeAtUFu83X83VZGk9YN7zrmwdc
vHkwJm+n9Jp9Ip12maSTVUUFOcIYU7+pbUbo+qgbXj922DodgHYFuhPGLbPIaee7msy2zVDoLn+B
iKEv7cYKlslJd3y1n6Z+yse853QhHUw3ZUkrFDLbaNmMmF+yrJRHx/g45eF6zWt9JD3En+nCLGA6
1/Rm/abkyp0A+ffP0hT8GLHUdtffzNAS0GDZoUXTTEqu9EzTPOQ3UIx7gU8fKPknU7mM4B1jYK3Q
HyjiJdkcHRf5rrUfQeOa3vJwhv/ra3q+NPOafD29MwBGSoN9BUwrQN1Nq9kynKeSr7blAb786wCf
f/UaVqCod6EouJXrcjAq8FGmfC/gsu32BwNR8dk9vdp3Wfw9AlK6spCiRzjX/xviEdzFZyivW8W+
n5WFuZOMAunQ8gK6BVq6OXGfvol/n1fZ2NTgWFjW45iiWhPaCFlE8fKS+SLEVFHO0d+baczMZtue
31Gq/qmU/8rf9Uart+IZCYY4CBpGAZtSEGoV2WHGFWuIaJwkCDwk/xNS3+DF+XVV18D9EOD85jNi
tMYA6ez7CRSpLxDmJeTk0/ar5PUG1/iaZLmLMFGxdLNOfZLu0UItjQIeH915tANGgmqbYmCQnkp8
Z3OWFN0LLaSGPg9BJeIPbx0nsGw5Je6SxW6AsO289phKRI8DJjx0EjiuJuIKLK+Nn5z06NFtdjsL
DVjVKIdSI2yp1CgzpA2x4LQH6IuKITlgCcyHMf/nh/09cveEo7TLmTpB56AB1ZVFGux37sXwV8Nt
R92ed1oo9VnPsWRS0GxEyK3NL9KlskOMSorEKn/AqpjJpAxYsTowhGNuOynQVa7XxSRDNe3xzaBU
WYkIpq8UrYl6HVnhcIcdQ1d5g6mmkQQmWf45ov/IY369AlH8+pVqbgmvS/hL2UGP2nbK4C9vcsc8
/3npHEyyCVLzIUsPHH76djVV2d4dgIfpLY8ovAulbFk1RYgt+YWGi8ehg+3pvLt3uZfFl1Oke5XV
UI0X2NhyvVsdFCEcN07FfEw4SrPny09MJUe8iHIr/fUImh2TMsKHhBJbqeBDmc8+xSji7zA7Jwwp
7P4o6HvxXmD5HeQITKbqPdux29gE0SLSRARQgp0uOAYFICvdNj88tZDENzurp4F2/KklRGiNDBV9
mLUMZodCNmmhvrRAimbipme7nHp6+/DtQ41WjVXlBtBlbv+2SIryoACY7nShJC2o4CwaEEYFkgnF
/2INk7kJjhTF2qGNrkYCaoyASrebGUNa8d3fI110YO2UpP11KzecJkf8EU47MCjtYj+y2ods3OXk
DkWO4iLuvSA704EKfg41w9zGlMHuov5IaQAnCwB+vPZRCvqWuVbKubffR4q9Qj+0wgrW1aUEMjUQ
Vows3uVqNdKwV9m2JmNw/H4TO4d5ZKZKLYOsIgQL+sAxqO38eGzLmnUljHTSHtjtvkHpeNRqb8xX
cQVldD9DZWQRWuwO1xwxArdjCqqawq4LXDKVGOUZELGQQaA3wf5VIkRYvVZ0lwbH7U69qUY4nQRs
W7HML1iJ9ieIpIWYvQgehkB70h2toEpN4CYpJPbt+6dAfw6fRwwn+hpFzkVxsQXlBQhWuXxkKd+s
17XiOFsYr/da2xofU9x9rq1lZjZt8JRkR8aSKaglTq7heHbuzh2p3VWaaawnUtQsePaJkSn7enlx
OJUxnPbWMybM7UjmCa2bLKDQsdOjTaEsq7X4PDFxd4/L2d66RWBbUwq0kfRqOJO52jLribiEoL66
dGEe0U4Yy2OlHxWioSmhJ27RhRYBSrHXvQAMMaFd4DFKWKET6bBu+v115DYtBHx3iV4HarlI/Jx2
H08a5rOltTaXcN9TlwpXMidbS7wFSjEc43cmHF03Ha94JvpneRNl2bu2TkCsrGdVaXl2ahg6CbJF
XoEj8H1xZ7WIIrPYZRarQI+m+23nR6O9gqBTcAlwnuuNcbksvTQYiznQsKUnpkO6Oofi5+NmxltJ
vd3yqRxhsC6aQSaWE9DEM1jl1cGW8F9SwhC3EupajG7DoyT9KpR/dkUjX1CD/2Pq5E5Abh4kFpuk
GwkxNV585RK5yq9BU5ryBRiBRuengbcrtp/l+CG8jjvlP8MsUEAreULsLcxBQifH1lJLldQXeq9M
+LL0BXFrqFgg6/rqFx33SgiT5sPFFvYVmiL/LeE8eMdDCatQVlKBNex1IAPLZL04z1szagWEhBqN
FiZuvSEwYLw5MQS/hMIfkt9GoAVBbspoJGQLWgmoLZqhmLZLecB1gDxkDdZDBQEcWXL4lK01n3yF
3Xf0vUHec0sDilu0vfVEPU27lje0FGuBdy48IYQxbpEmFBiHXusE1WfIAfr58jgwKyWj6il8IVPW
0y0MGOCbr4mifBH4Lxuawg5p/HtdrwcYUhoocWOYnIiBalhgjRAFebjM++PVnZf5Fh24YVwHgVc5
EBv6qiSFRCQ5wjJYlrSKu3NJtwR8FcgHoiA9qIAeAEYL7x7046T0reNFs1+PaPVitSuE3eJbUszZ
TvLcsIYVrYWHxy7YE6neTi7+pAhnbKoJ6EMmkEvxAqvB95BeD4DgOP0BxSqrjzLmJBxdIKZhYxq7
hJGqM2CXTpV9t77qsdWkiyaSbKtdAnikXUpVtlepFySqS2ud3iM3uFs5yTQ+vgUg7Bof8MirbKko
xLp82Es5alETdTlPvEaV8IRc1TEiX6a6Yo0JjRVyuQ0+0Kg5JLb6DtDHHHuQZC+GjBuVPC6nQuKJ
h4iIq0SwMQDZkBAeDdwwO/jiTc9Lp7bJ/JhMbDir+Ysp6Ofohi+SN4vHRb6/oqTYrkzIDxNOHVqc
mxE7IQeDBxf+1QD1oZ8GveL7Cid1r8vPLKd9SustG8P+22+lux9zndfCcn7fClAcJ0FyAXNxwEu5
cFAE8X0m2bVgpO3Th3zTyITz04eIDyJ5calDryozB7WvTIJwcXMed0LtXarye7qRqbo6mbTfAidu
2erobpYvcEzM2JwDwbg8oe3k62W1ZQC0Tp4X/nXwiRtrpy7UNZQQTjRrD2jU3MamtZNYMETOnR6S
9YXs+h6Z/WzrMbK9iGqTnmjXh48DmePx+YcHlr+gR+Z2oZpk7LUmd6EnCbvko6ED6zHgTREICxGX
BSCdAgiQPiP3eHTggks01hv4m772NRZoedI8qkxoMMMimu7EcGRuYyf8vzf2cyuDRoH8zXouri6/
/QHggBQsD/DqyoEQeW4DY+JXQ9MAWQJ+a+Ja1AlBTPv7bbC7AuZyk1I7SZQ0RYrmu700xSoQfEL2
lC2TWb6g4iLcyHVTTovZiYjsDuA6JAHvisu9V6wNP537hFo7U9Ng8w5xlirpSaexzXwUysP+RDod
UojN915+C1/p85CHKJMgRI2G5Yr9Qagv1Mznm12gtOZxVFDKpR7wIxRu9pq9hrqffA3FHIIpReQM
A2kP53iatObSpvEk/Nlz5bXQuLS9DIh/3OrRFLj2ZFQCcAvlgJpm9rcbG4n6ELmQQq4djZ0GvyBR
CS3r/f70ZwVF+097icPx/etWzfNYa2ABj7OlC6hL4F49nuU4LGvNpZI75TAGRnySE5KFvtDw3x1T
N15xwjSnSW2+VNXTy9XbZZJfjEQJtjiq1CM3FjhDRykiZbNJC+16FgI6u8A+zH7eIgxUSYQTdMw0
sgClbsABm+s4hy7k7K1iSnsUspZKej5Bpb20NwRI3KPcpAbqrzXlRxhKI1ScezC6ZV95nQfb9xg2
5rH+laSiqQ+LduMc1bx6CID7cqeb92rFlpRISD1IVTzBpDOSVFk1XM6A1S6MSjsSrR3/65saqlHa
uh86tnT9Wx7WWUQEPGJfkKMta1+IOcAdHKovecQob1VrALp1WVaR3taNibT3rkhvu2HVXRUvB4lT
iWADVoao5W7NqfW6g/2yxGNKp0rXpyJKVOfnivdaUMJeG5EVlE43wzXuwSqStPBsXue+1Yj7Se8G
PmfsrYe7Ldkxa9AG/idxTsCr1MvIxImQvGRYcuagcktDUv0J66CcYbu4iTFSlaW4cq2ZH9CWaT8X
sHIqy/W11KzvgRte31Tr2gvDdE4SVTV1r1tV/G/wl/WtE1ZQXHJNgW1iYAH24kPcr/Y4Sidhv6YX
r68i2k4mYWm6TPQgjWhuthwUlgBTbKZyi9pYnCi1gihgtStVauI1uZZYzlm6ylDZ6Zzze8XoNz3s
RClga4iUNeVS6pzZ3GYEASiXNYwjGEUYqxcN+JkZVqs0PnC54ljjYsMDJZMc3N0er+Ds6XT4n44w
+eG6Yihf1HygWQ1vREtPHTHup9vn/CI7tkEC1KUXXVQUEWkTnxQQsZzFVT/CA/jhJPrDxcDdN5n9
NnilUR/CYfj9wb2xHih+JbEl634dZtstrd04CN9cw1QQFXUMTV4wIyKBm/WCzH/8/CPNFoVpDivH
dvfC6o0DnTghbAKAPutIPbgjTzio+53MH/QeKmJI/zrvvc6UVHZ49VxHoybJkMBcjjCsOryz3bRb
k9lHbnkcWcbGzVnWaNlbpPKif0YFBBK7CCzlV/8kb2N1XZGVwgUp2rEHo5ghGsamrGArdJcRMqcn
i6NtnPqBpbc+paiq6kfoceiMFHMOa+TfAZbTWkDql9GItUPsG3BQxRyuAQNk0wC1Y1v3dr5sTOZb
DSWOGmOJei/cPROEhuKNE0gfL86Ils2DXP6sQ+3s7AY8fhdlQo7Am098KOKO5cMC54aJ6RodQGJx
k31gF+tpnGZPqkxL0EjtnCX1BjuUK01U9C9K12pB1dVBRTockr3mpU0dWiyLFboEtkt7jZeloUAU
G+h3G6noJxFankO9SxjILqh1vwRhQ9jleokIQlmhlcDHRfqFvj3bonhWSFzvf+oFxuJ8ttcLE5O9
2gjpfwcGxaf8kb9jTu897PDKdCFNQGEzDCYKZpk8w3TjboKcQwFMPpjoP0kL8Grwtb59AJI6sutF
NR5II6YmIExIb6Wa7aLVWxtBeuSzAegNm3b0CapNJdLJezsfilAMLOyXEhs6bljpsfBqsveML1Fp
k9gBb4sKkb59hRslSQtNd72HH7QIBHNePxAU2UjayxW/m1FptadWtw5ZEU6Uwqn/9C+3pyoxgmLa
+SUH0fZBlKcDqASeU0P5TV38Nh3FtTvrypC1c+q4ibVJ+fFKPjPiBzCwLAoo1Z7oB9rm+/dCXgBY
5nG0B5Tr3IxleYx1UWGurBA2oHdzvkorBGWMwPIgcet5orga+0VluFft3nyZTBOYTGBHQprxYNXo
JVji2A44c9k7E6ecBRBRjJWeoSJ+/Te5cAVM6LTCos0XXrPy48GRRMlsvNkKYLAUx3FfHwbx1HuO
U2T5BiIGv5vFo8P5sqwtsmqa0EbWo46bOnO7GzRy0tuRvixM6LQPAK7Y5V94z1WUixemJPUxHKLy
03VQcSSc29rbgVh/B/dNGXsXRVo7xfPJfMbUFPZkdnp5UE37mUDNeceMwSLfRLmJXcDbm+PdF+PD
bcGR2f6kHsjUf4NRu+7uwypoPKNA+R43QaAqCojQzydSgbpRKkUYT9rKPO0GhaSu3L8q28TmsYUB
6i2BttG4/xtnsnwgmXxi/CyEyt/NCqgc2rXxZ0admelmyw2QdPGMP3819BDO9G2OKzMBuyxAC1sa
N9NoWVhk7rYTF3cayNcXJVl2rtOdbCtXt6UWhzpI/Pv3fs8y8WWR7Fbbq5dxPWn1x5fUKHsSaBBD
9Fg6XrGclLP/On12HYqzerPeQUyASeSwdzwJ1nrJk9WX+uQc0uMh5urk9C70NFQxAFtuut7LfMQr
J6UPkHDS3e/YO7NgqViMNyM51+vAibityuEqh4Yk67XOwqudW23FwMWyQBKEjZBoGR6wDIxVCJgq
diSVbVVHM1NP88BPIyQI/79JtDXq/Rm2Ha+/Z1/NBMYuUilcXcBYEUle7TTSQ9Zauh9xWYfgCzKb
nHydO7wz+wzS3Cfu/x5knmA/LeL9uel8ArfxjwlXd3+C/ok4LtQLWUbVBTmgLu9UvZDHgappqH27
4dOZ0xtK7NnyvYz6Emm1ivg8CPc6Gvw4PX4GtahoWUGYxr6anF3kLQKagfd5K8lSQame+2R8df2N
sLSj8q/ieJv1VceblVrXf+UCvI/hedRTS/Lf8p+rDER5BaVG274OrPuogDkSbCVV8QTwwNTL4pMY
lYBcro7SfyF1z6ek1V/BjR+n6QK1EO+xFJ3ZMkc8iR1tFKIQPzu05WPNlf75dYQb6l6I+zk5tvgr
tLfDvgjE6kb5TvyEGjy57ZdmDkGH5vPnty3krFtEROdZPGyzCDxksyywrn8LKjUyQWEQoyq+Yp6H
aTFidhH++aVl6CdZcBpfHGwMT05WUkKtTwGKcy1fea1eTyyGXksgyPwJKdtJcB87dJz5zTEBuian
0otnxE7zPZflMi1Z132g4+MxGK5hkZFrqKrD2VF0YxoEsjVZs7dKCMVf3wSXKpdkTzL9QcQWfSoO
CBH5EEvnL7dcYa3gYjA/j0IVV3Bi11NRTrO8DbGwYNLNHgt7HQ/bpCQep+E3dHF3WkQ9rM4P4FHL
S0vfFc4hu1xo9vMyCPYKehwfxQzrH1iK7Wxv8FL4OiFoZdGJ65jZIpZv64dc5TPwaB8+NRT7oLco
WfYBcK6rYIqnbUD0UiUXKqgTrU2yLCx479BY8AI0w7DzMiXYsKKnAki4Xj2J448iXeKzDtxvFmk7
X94UjwzLz9SF80B/KGKuwb1apEXjL0fwkLQ3JudFrOSre6q2W5PocKylWX38aihv6RvVCV+kXmjl
z0mPZMR8DlFmLNFMHmMwz83gQaCPltx0pZKu5YPavmymFVOjehDRNdGUwAhdIzCAiSQqxtua7Raj
k1NiLv7Y+29niCOk4N4iOfA2cx/Sp0/RgNFQ9TmW4v/0N40zureuf/NKlJetNmOTkl7wWFzjKUOa
Sa5cPM4XaKGdxLTXP9CDexO4X88rMUbVCTKZn32A0r4pDOqt1EyGeq/zXN5vywYwaIyKCM97osPC
6VoO28GaWdN1AdK6CVy7UNdibS7ZKaM3RpJjxrBFAvpILPNOda/sCo9y0DKXH7SxnugkPZyKiaRR
2PnBA/vauXtrZhIbprSyeYivZ4JEAvsIMPnjVLmoxqL5b7uT1DtKT5/erQ14MhqyPGzO0EOJLplV
hRPR3Soxy1x67uni6EC1UYSbw6n/uWuyslYI7AMUqPZEN8dmZWPpv5IITKK72ktuFbuR13fzLMzZ
C0lPfgHp9JkQnMvsC/9Amheggu5CCvXw8nKesv6t1zDcbp6RjYLFOZ52s/Uq+hL8Yz0wA5bWG0WD
u48IawyzcNY5ECeRSVJB20GasmCwWiD7/IlRcEMsaxs6PMF9uVryYxDTG7aLxFKgL6xpU3Amz+Ge
SFvqfjASIHRC257ZDpo67k/1nis1sZ+xA9FMRnYo7KPLa3m2EBv1kJ8g2XLMW0g91tT9sYavAXxQ
t5bU7C0/raUB2UTCHufIMW2yYCQSL6tQp2lAF06kTHX8MNIabGebim5hVEgUrSbE1D/i0SyVvelE
q4CdrG1bxukollgbl+IClwwwlDc4neKL4DJ1ZxS//fHWjAbkwf82zkPE/0VV+v/oPb7o7aU+THt3
C4oYA6ACrdWTXl6fCG50i7pM41slYvn1HUilysm236H6kHMSklJR2C1u79b1TsdBIqyknFhy0Ab5
SoEo47fQvD7HX1sJQqvFFc6v9ZtHxEe/XIEihxco/VS2GcCQ6ijxagdlbu+7JSV6g5MdE8/yYXeo
jbcy+koSU1sZcSOcjrsWrAgxKT4FbvoEDdL698SRgubWREYrwanwYS4wRiMw6RziFgjq3zuXSg/K
q+rjKdJpEPsicDfC+DQnlKHl4guD+PSKXjQn5nfArkDrgek+mjB/TN2Y9z3hlqfjgxPlUPBF8NzG
GEHYBBQ1GVJdWgiwdqVcmwJzgP8/h4fFlYItAO9k1pVHuEzrs7ev0orcqeAei80g5isOPLQqMMva
23PIAnVOrRxMQ+DenUXMlytuj4471UhCzjCcUpFc2tF/20YxPwmzrj2+sfh397+ttYBRl/8fQjZy
WJ8wNY5fWvYf5U+tfLzDv+fdFHgymDZ/ZGxDu8eZCqD8U3hJ6VPKJZateEFj+907qquBThU7T/lM
xZRrimL9uCBSlUo+vR4WkLDd8Eo4VNuiZqOI52j9VHGMcXNPuOsz6X86WNf4hgm6otH29UOAhFlq
iIMQQTVCRvagIIAgh/9/JsTCeMZpMfVkkM8d7e1ICNPuJe50baj0DYrI4jtlrfkC2y0pbrchWhYx
Ck7n4uywKb2IvWpuTpqvlLsgru4sVURPtAaqMlajC/S2ysfhp2w4gOQ7vo4Cl2vQ2WXMk05Q/Rj0
8wIbjwYk6js1X1Du/PhBYdc7LmHdC3ODwlrkGlzD5uAQM7DHI495aW9oPnpQdpJ4D/4CdPAD0OVs
SNTlASRTBkl7Qkg9WR7XloV20nED/dtIrbvENdOdOenCEpaLjovzgBbBzI7RjDy35tkuABF4uFxC
Q1+mX2Lzs5ofUjSTQzrpThdRw9csSS2HDiAgvAKXG0Wd/ZA8cYLRnU7mitCeia+CplrkG+ax5Txa
CQkEneAXqEko5IezLk7FbPUIaapcMI8sbvUSbScjQ1Ur7ub0Uxe0TMSyQ2ft3yyzsiu/TkFYoM/Q
dwohk9cSn5ByZjKVHErVYkJpK37yRPHDtyf2osyS1+KaTtCQQOhQx21986akdXWTcTloBaCtZjpH
XS1mQfYwbQF1cnnqLSX0r8vZ+S0TereoDh6/bIEdaGGEOzMk+t0Zh/gCOgcm+3X7bI2heAWYUD1v
g9IX34Q3+M9tyY7iPgQ8y+L2MPJ+nxzJ2ZJ6MaYycQEb8Rc9W/yKzboKOraq9L6xwO+bxIlPxY92
agmFk2l/EOvAaNPumnY61UpP52TH4WKkev9NLyh2Ib4qnavyOEZpvpVeFB6p1pZrPc/JUyRrLnDX
x6veJupdAZqrFjgXzkqmAct9T+P0yIrlV8GdPDvaT/9nqmRC6yr/jgPAGW2oXJO8vp2Eocrc0GrD
U2wqJQqRNiDcE9+PXrc1zt5wE7qNMm7ivZlqVft3tXPbbH4xE9sceEtanMJJm/evGstxmRnSQxTp
cHd75BjtDr1ilHlXnEikWo5WTYGad1bIaF4F/HPimBHMRusQaCV8JUluEkxEVUmfN9WSQ4e36XLo
F2qv99vJWECFd7aizeNmLj7AgC/xPnD24aaAD5b4oNxe2UWgnt4jjISp1LLh9IIy5pErroeQ/6an
xyR7ZPhryT51Vcni7A9xWuXN2aJ4Bz4drib6hJO2kWDrFHqQlx0nbfTtUwvMnVd3gIoncpKVVBZc
A2pBYZdzSz21p1gmgqjQ7tsxcg4+FIL7XhWdPcFaiEboKo4DrBEvkBEzGZgS51+J9Ikm2w2Sv95/
2b6j3k5B9ZadK31k5FCYrHCS03qfPLtZvVINmNCWaUJKH35dCLcrOS2vi4Vw9TCRAB/IrLF6p8ol
kmg4Zxe0PI7v5dZQk/XiVa3YUYyFd2ADPU8A5l44fR6OnNspf9DlIN/guCX4/EyqaZvMLXQzqWHx
HZMnk1BnsZGjKmHYNWLabMnLTGgD/uQTEr94+p5e3kbu91CjHPIAcn8CHkKTWMJAYZ6ZbM1uMh83
EGRJmTjKxFSa/U3DfdX00NruS0WPMLT31zqD+RHgPCQRReJYinibbmn38dnRgSKziYuEUiCFiBL3
NHeX2wH4vzCQjSK+J0LqabAJhXo1SS1+HsWnxsv1spd8D2ptXLbWAhZTyV4BvsbrjLcHjwsUluYL
oa0HscMTqfx3mkaWo+vJqzvsfoHiEqtNTBqfKEu17LKSeG3VdWVAtf6cDeANEzoVeXEE8gumOWjs
CLqTy8SwvXUTNIhlHfhj0+moO0cO78gFwQAmTLp5BQ0VkksINxH/Ofe7o3a+QW5hpDV2lc7XQWjl
Sm4ELoNxtOEMNyhUZqxPl7eYh/baGjxZSV9ZT0/MNgcG2RPvir4+ZhEMyfIFa6eLLaZtu40kUV59
avD3Jt8Mo3BtScjcPjqYFoH0UW8UuT4udEIaUCoazvLyMwHOc0AeDi30fFDsVZrtr2UtlUdj+iw/
FXrW3aTH9wFIm4bUPD309jTV/T0mHg3yFn22lHkuqy2bi+yONdWFOzCTQ01rXUN+6bN/7Lk/MuZk
Svlc4R3qmi1rF+e6qyy+HMp2lVN3+j/Byn7a79nd+h7G1e62urqcuwJwd/lvhaM7aXpaECahbRXe
2xPJHmaXBfDrNMka6l/GuD5ud0C/v4wGXLj7AToGIsWBQZpvC54oCHbRgNJRCdyxNhpAHegXllJr
8hStPjRBMTECGM//slIMq+wd63Xv4m1z3BBIRZcMzdKWHaOnUMp1LrS4NYoQEVBVvY4QHs07dPQO
YPoamb59HKosNmOoSEmwN+A2cdf9P0gbhgyZPg31l26Lvexcv7FSk4yvUj1uwfVrvLhfMAMFpa3w
WIsDXHtjZiG7OohxLSbScAGu9bUUcFswNz0vpXpkCz4XQ8TukdSzIi7cvpHwFjFzt9B3+s+XObwV
GY2tt4cw7jecSGk5nae3vjDa0qVtMvpiMALOjBlqMfEtL5NhrbM8LAOHpWz1h/xQ7cjZY4DX2uyz
u4rsUPnqIF0Ilq6nlIddPcnSeQtZQLvKho0NsyH58NbQ/VqgeHhYifx4nVNNea1I7Z1bvGcsi3e3
Hust+LKcjpJd6/l14QAkzJr4AIOWvBI/GBeqs9Fw4+E+RETkqxuNMCgocKruMivV45zp969p7iDm
cUjgKC42+OUeOqv51mGt7f3dqGEx0cIJiVKLQjIhxGxGQyVV1xaW1LlQ/y1ZORHaFAW+WT2633Dg
3SKg9G4GAC5b8LNgzBbeM1iohHBjalTVHU/KRDRx9gjRlp0Y5I6OM1VbRLD1kBHFLRW0FbvBTUSR
Pm0IL7Hk8qDD3767kxIxXnWoqpJcukUflsSzzzRRLb+BYhjb8shI5YgSQFrlJizjc2kX0a2norV1
QumQtRw40ylDexG5VOOA0lOXhc3RF646Ul1Uv7GRayovu8kou9UYySloB8bVoQtxe2gsBT9+rKLM
VinUeNDU4gYZCJ4QdhPt7RyCA8F+4RaAokNtSuspwyDVTzJzwADcpC2MuzDCRyS9vFFY+ghrIpPW
JP9USwGrP0IZd91hjmwlCPxyQPnPEQCwpj8ewUsrk+hGNkZSPfmVXo4K+yAZzZC6dMD1z7zXqKLB
ubMozVGP9ER3FHxbbUnX20skuV6TJVKLh/w9/CxIxzfap/KFRpcgQK6/wUILiB7VSGM6AJ75Szw2
6kplmK1Xw1ZEY/bnVXufChIkVm5Os3TrR9NVPnOqZfOnynJc+PyIyi/bbsCAkyd6de0Ogc08nYgA
fWOHcWKfsEYy60LzLnFjzW9EvKjDp3+HDc5dtvkOIxhdVOFuh/o+3FV0CcwJ34VJeaEUQ+sHONls
HcgPcJmEeGBYhc7YCzBeUx3g+yAGdTgywWyn/90Lb2Ck3oNRDkmc9jMxIG5jxlhnE/zSX3p73C6H
fCQwcVyyF5hy3+SGae1XiuSRF3qK0U3iyg9XYi/UC9DeALI0Ya0kqyQMRjTQf1cRJ/DCIJ9JO6vy
mSdL0C+U6+hKi4IzU+eEd8dEeRGGbf1aEKz9hOfIROcMCYpDab6ddcjMWBfJgGW+cVh8IwcOZZ7H
FptTXLMoP8PMWS/XLs9O7rxSo75CHutrSInaL4PkPcvhxuE7KD8j6s34drQW6zgzRPScHL6YxAfg
FkXPa40ffIgO27tIeRdK+gwdaahOB48Yng2yMeu/rL5qPq+WD64IRiEHjDhXHXfii2Y0qVSGhVJe
+PfAq+gl/Yz7rW1IdegT9NyxpGsPfmbpmSLJeIJd+n3g+s6c+p4lDJMUJAsdpthHi/Oi7o0ur60j
7TnkVnznJaMrXWb0Ub6QfC8JIUCrvbnOnNFhMfwz9/e1biPd3WlD6uMotywJnrWcbf3N+3H1MgaG
iKgDOzbx+tbTfBMjKdQY0e1IyPbIMc8+Y515R2btqHaZ5po5HBwnUH089D0E8Dv6zdzxanpuxMj7
5Tqw94kHaZ6xp7GPFt3sIG8r4VHD65LXYyooYXIsBLI+kPvzVwiN2W8QGK6GFqjM+EdYYIbhTf2R
QNQmwuDknEsaKCjov2pXqIj/mxD8xiNGgjGnKgImFNgGucFqosLhXL35oFazfTq5wAfrc0T61PAR
7nO8V5jFgzc3hHVVIJvdt45krvckNcfB+SKsN/Lf7Bm0Ft0WePC5YXTbGWk4ud8agv8VV1pS00ud
cozUvd+BOicnV7VF3L6+PQhsuLM/XSKaotmGQqf5xoq/pu9WsxdUqdkxixZUtUoVNE+mkF3GCYtX
25DU1az5tiREQKuekWSHyf7g1MPJMuPAV84LuxSzSEx4Wk/kCHETEYT60+PX6uOduV84SHsy4lcu
eKd91OsqsB7PUteo2tagANcEVO7iNPpLWwJLQP2KY3HPhjqJyQf7WPJ8+g825SnN4LY1nELl7xWU
Dm/PpXNr64o+2vA20BYBWFqTj4uxNkfarTnKDQvmBiBFoQ1U3imsIjHrdbWY+bCFXMrdqwgZQD3i
eW/5wydgvI3cmIBip/SfQ9OnMP5YAAp0Y1t3gD19kL6zG1d9eANnxY9wBGX2Dw/4pQflYk8yAytZ
ZQ7Rd6RsGfW8w3gC1Ns06l/JQSMB4Sf8SLUiP2NxM0Gs2RcX4womWqgFYwQe+AvfSrIToz/mu/Z0
gs2yQ/dmlRjiU1PYAx0v78NnzMHAZEBpxIS71IIdDxrs6bS2J6FRWfrQVM4VZqLS0akguJUS5bcH
kvJgXIV+OY90SzIQvRuasoqNJ/zDtGddDjLNUnXvaxLdvy5TJ3evncM11iAg9rbpsjeh7L/3radc
kjhgz4cx4xZ7GjzUb5wtosUG8J2CezEMm/vgfWfNKBuNknR2GxggCsuC8x5v5ok0Yg7RBhFv415u
t/Y1sH1GBDd/6ANQ+ScDw2p0F4F1dkvGwfEMCZvPRf8LiyZ1melC0qMtNExOJ58jCYWRn+wytsNV
ozJhtbixj9bP0Cg4ZS5twQMtEJ+H5zyiRAoWX8ZjCCCidUnL6SDnZepKhNhpnrZ68nFhBJgmxdij
sjWNZ75/1sDXsG5e/2iXFB0TGqqBFT1InS44XJF5PMTJku4rWeUxsyXexmbkTlfZPT2NhLSz0z0V
XOu/9SoyxFt9j0hNTghLxhCiT5Y+mJtudAKzUoqSSVk7v3CBjgfJnEdNKbB4Apb+UJNA/0DR9y5S
7G10+zdA9O5MqGsGDfU+nurIwgHGLDCplmResA/3YQx6FJ+zfsUM9PNYGI9ZHGcz7dK2s0UPYlaQ
Js1QlIuQ7HEGfV9ZEPZ1Yb25xDzZuGGilPVOjIxseZ63h5gr8lAHVxpHH4byR5N33uHylN2+oAIt
2bF3sREkfsNQxgBMAAJVopArr+m+o2yuQmZafJyvHOW7/McfXNN6u8gOKG8lCJ6IJ4AdioMgsmPU
NTGpN962HHLUKgm6L5LwhX6pXc23XycuuD5HRIPe6jwmUXoYtP3miOEdS4GCoZdXiF0lq1px376R
jTKMhqX7Ea0u2wgq/Pnzo9JWKX/rH7GIF1NhpbKtzxJsFL0mrq9fRdGITtiI8oxI0zn7b42d/nMO
pfuJ3GiTA2iAw+bOTpRST16P2HWcQg/v5/+G44EdhN8KHToKNxC2brouHySS2kB0sssjROjxxCES
vnwmfVMgP+aHN9SQkV+1AmVsqoDCZLKwXd6DzmM/6T0mRWREAnwQ0hSO1bnEd73jdJ5lwNTjMj5X
uRV2ChmaR7bhjMBzDR6HzO8lA+a7YEkmOXs6vF/3ZbeZpv45iF8Vj1uG8OuuVuNHk7T0qNVjSRdu
gKMRAegRbgtpsjnKBiD67eu2k62BdFGkNHErBqL/fI7QNIQ7mlKKWDd6IaDk9yNcX5zBD0/OkPs/
Tdc2LKJInm1AIbYTxIAEI4UKPi1bbeTBJhQwbPRG6qjkBkJrlJdROnJE+0RxIfogKJSFgSTb3hxk
994Q/3bEdhZLrPH+lVEZvdUy6iFCxp33AJnDcxhgr1SqRv+/kCl6gcbgzsswzzO5fYhmn4H0Zu+U
/CmILgPu27ILRcnlTawWksKSnzaWzAw1gYl7jRxjrJGC0T5IboHwiJjRzNkwtqgwtvf6bzdBEKuw
lhb9q06byJFhpDOsWFq/ttnME4buYtO8uj3mZD5/HnXSi/HxPJplYucXLPAMJVTfxStfgyenJqXO
9vxmK2RYweJc3GXwjG0JZcYXaSkLVKqu3sO4iaNaIwhnHSkE1EqTFERhdYYS+brQ7dQ03pQyhf4b
l04hKFEwibgJU3bPFx9VYrR1pDZt7x7CuUdL0QECFy/qgDp5Dr1+l0TTTu4SFby9jvQ8HtZWa1xN
JR3ffuz6TRvcCZq1SL+XPwgEBdVM9f4yTYewP3CqRejCmKsR9Xa6vIqNIA4wkI3M1/zTH0qij1co
pJOEn/mYwu3el+B72aj5/fChY8BwiHM8PzrUdR9yi3LgzVJlTqX1DZGDvzJCFjNok3Eb44bJEN1U
B1TGSNvxNf5X/gxnh72jyMYJko/lD/2fO9mMbwT/0OoW+qcUOLAA87qhC+DSYYUEKm7t76hcM/O6
A59wlFATVZ+osfyer70/SVo9jmDMMEDKTdJfHzK9Epuvbdz0NTqt09KLy4ufIORidyrTw1mCsAXj
T1XSItb08er2x5QPtPTCKkyDO0tC8C8e70xIkPiIvmCHDUfKtbgssW9mJ030FP/DHtVpe+zvkYqg
D9ZhnKfMLOSTCSH1XqV4XlG9lTQ4hf8rqAo87z6dnD7frqewCw7NEtkKSdgseBmaH+hre4h+WvrI
Il4VOvFQmb/hYGowcf/EoHmtPxLww7HjiYVDYtroL6fTw6PjdTrWm1LQ83GtiY8KPckizmaSmaHO
DNyMw27Gv2kAAA2XQCXURPW9+FI6L0JbLCZ0XXv1o/vY9kLKjBcRZnszSAPk3hKq+IcuLreXs/mb
HOVveGM6WoTvKGqrbKvRzQqEosZJ/8mkONyiVeNyp3cPvFyk30oiVIDMUf1xOIOnJ8hngGZapfM0
AtODEtmc+2GY4725Mwrjm+QmRCAOgxCwAESib75zZjNCpg5BgcLM49yBv4VziA34CxUTSUcZKO+c
am6T5z3cWakNY1nrPqpqFZ1ZUdCbbVM1u448msqvGb7HEFSTgKGzDrsgSD3kXUXSvyfTHcznUB/h
Xsklhu6V+BUUGbxfBZSHJgQZVhTzaYy94XQKurvlM2k1hshuAJproRoRf3HNJbi+YBr6lDKFy4PL
FhdckGRyyaN30NcrwtJkO5CTLiEZ7XxNaHXWY3xHTFgFDey46AJP3sieOB0WJie1Mq917ljGuZIn
MVgCeYbd3Kg5Aq1XSCR4s6zF2B5INgiP8Gl8kZrCONIWqqgSaunFNBVlHNBk65k4Ox7z4Scl0HZk
pVnunmvksRNLpJvTuQbK1FvNmxOnOaP/YSRYMTDEBg8mukti3wCYfqLTtK91ZaLp8hHfrniWEd8G
815xzFLOvI9I2jpn6eW+qX/BvJ8/WmgLNmPGka2zPx7SdvLRaNpA9Y2AskSr8083fVA5iMJImZH7
C5bJ5dvSnBnd4U2SYt5yTFw6lClskA1Bw1gG8EsNMdlGGN4KTTRJU47xX4lRvEjf8PyAP2LQkE3L
9VITQe0Gu9x3UYKRY2gbLvkfBsHDsg90m1Ez5BI2C+5ka1YKYQfovfEStNMGvLKSu8awQTnGViKD
kKKCsH8Wud7lMZcpqV6eQHqto13sZ+i17s3wq6r9YWJTrbb7q4z+qR5xhPhpd8CIoFrErl4Q9Z+u
e9TwS0LLyOIYwMkhjwBziALbRTY2GMYDHTROUD904sUxCaDSrfkZqTwF1SCaijaOq74R73RUpzP0
PXxXY79zjrerKKfbe9ZI+MKHsR+M8v+Ls9hQsXXiy3+mYrsju9uaP18BgOevkQaclWkPRI/LNphr
p1gbeGcI8DqztGA7aKKV0mCSz/LbgLkdQ01SJ3FfqygdUoWAhd3UYEEk0jF8RDbmwaDeag4SY95j
zL9Bi4VZ5Bjt6tMWPq6ftGMdsB0iWD19cNSq+DhWXSHoIenvIulCcrk2PDYZecIuBWmexcYYNC67
j8xpA5pqa8MSGf0e+vJQS/lETzSyiPuVkwC8RRIqjAE1nsdVQovgVTrsDbhecu7E578FU477v30T
Sf3cPsjX1RhHK4p3plhqURGw+5MlHXAHFEm7dsYo7/rL4XsqFbQ86YGH3UVG4N1KWEN5vgIZxDY5
lsUAk4z4fMUo8SUHyTZvgJnV9U+apdyUa2JhS+fSh3eDXrHAs6D2p45fnMBSjwENlL3F5RDDAc1Y
bHGKAlMY12oIx9nbtK+K7+SDWNy8LKne5mlp3tYfApq7Cjsnd/Ja2wzHGdPIFfyGs0al5UHneXTs
QtzB+EJvr73wCj64TpNa9gOYvqHPBZM53jRNwlJwg74hkwKKqdaexLVyFVGw/d9pIu9YECM0EDvs
i9aNZgSx/aFdGj7UzjoqHRvg3Bvx6MaZkNFliQ/gUnAyqNaMeX+C+Q2CpYmiOH7L5+AfjUU2aEmT
Oxyug3ksyMwugLI0pshhePpIoVNWV3dzDxbQx8Z5qnWogAVRuywREF9Uaa6Ifd3FP0qWFTnL2IuZ
76dw5Jfhw0HjYsomdFRZQ3FXnguKcf3Ng4mYAbsooaIh4DHAACLKB/sEmYmQ29mXeiI6T/nuC2I6
DLtsp//KNqWosiP/VMwHq2ibKKYEgAcfPygKHd1xA7xYzbnXlfg9qirYc/AlNEtzcRU8GJMX4CL/
wTj9h94zsQjrrQCMxluiygUKkaUJiN2zbCaDMNt74bUr2O7zU62fO+JxVmxga0keZI97XptpI9DA
IKJjt823lLFXuVu35VU15RwKuqENRJ8y7DSS1KAUE9SS1tBZ7nGq40fsIO3IhcID0gp0cdQflDTm
j10BftfTvCRT9vGBm0wkt42y9pzxAQl5fvEhicdEU4BfKgWYvAjKT7tJom4RNnh012G+kXVGFqF9
eIzOx1kSxFHNta20U2hcRZe6C2JmV0apjNIp6toKNIl86r9qPcr235dk7ZwqM0jhLIYHWQryqr9U
6XIC8I0mE+0tjtPM+9+uX8ufyh1HzEcP6tcO357edkFCJYDuA/xcxqrEukV5oArJg4B4ol9s/FZM
TA2eNHiaFgouqEt8hm2BNmzkFjyVd3xeK3xfMZX9/QFT7XqdEnGzm8xmJWqIqfTPKxxLxRDpZz8c
N5EzVX/xebwLPNABtoZKYaIvZ1Ko6s18qC1AkLoP7B9ma58254+o3402PXkZhCk5tcKnMnL3RRrz
jlEqLbu3IEMcePPU4XBqhIzWT+ejsvcG5hueDCnnXwmEIef9zPDrMRihAhwgfpjCNIjWnwUh6vhX
/lK/OMDTMpfR1552T3Gz7135iE8qEVnbj6i/6RPCZGIPKONZTss/N0Sj2/nKG8fdVlXMqlFzXtfT
evs1+FUK1MFZ69aTHQy1mb03OdkSThm9WCYEYETlzVHeLVz20Zw/3LA5K0EG6+vMnjXwhd7LuNIw
1kZ3MV9wVvGgzAefeC1xaRdj7B8mD+BodeunSJ5z/X9hZSV16tJg+M5y5oC9ifLLvZU3SVpF6v0Q
nOUeONynVrrrOdyrGjtpm1PLFpH/nzQe4TmJpHsla9jk6qDn57rGTkB6L6fi7GxrWXA6N+reNiwC
DqrxJo0pSbGd0QGZX/8MziTydt0ab51Rjz9z18uQVezB4NwgF4pvlr0yhEnR9KKVGv8iccBh2kF9
rYxyPPvbETUJect9d/7EWS1/N+hJ1wRIQoiFo3XkvUnWsk/9E4kAA6Ca/G3SefU5JMrPLNVJlUj1
zuF+lMwI+JnYmOs8wbIz1xL+dMlueoeoeT9LI+WgUkEE+OKviyCt2tU85Qn/7MrmN3wWMUDfhRGV
rWDsNexn57e/h3U3W4eQTAZ7X8A9VA4QUzO0PGOHBXpJt+WIjt5PWg9BqfYGc/pERpdtqxXIbuqT
KjUw/bdprBox9PLfIpZjKM10et1o4TDLuRVFRQKfJ9xw0RAud44YU+0jVaoWFR84Ogs7YVctffJk
8ChK85SIrknTQdlZBBJUikYhKI6qXA9opetcop4oFI4tS5pwoyoB9v7n2OyF4YXM0y3Kakd+n6Hc
gfDWszl38b2qPzyudr+cKk+AKeKiYmG3XVcVPYCqDxnbXZz3cKl/JonpHeXO/QVIdqK6PcN+PQyV
2Y9RNzKj7cab+SOW0pAR6eOXt3T5zb8nZzYDxBQdXTmnHqUjidZPPC5xhgcxbLK4Uv5i3Yw2YIvO
13hVis428WAuDpi3HsiS7uYNiINvfEbNONCxnJ95J54ouzAlMDE1fDlM1P4SFmvw//r3PrMUBhTV
vBeijD0iYuEQ+kN58XV5OMx0E23IOhPch34cfFNl2cHKbIcsbPRv+iwaChvOD6WbIASKHIG69i21
bplPSGyMfjFIHl61IMK282VqMAQzngYmdRccWKsCXueiwnPNzWL5tlOh9sDQEt/e77nBkXGhyd7+
pDvn4dAvI7GU6dKEAlexvpsQxLzB1U4cOnhZHksYje/QjFGogYhg+Cgn6QcXFEjvYcQDZC4Q3veX
NVa3hzs6jAmbFtz9YE9JtdN3J7IuAHyl08N7+Y7rWouZjy5A7jyoGGMrq05uvQQe4zoQCcyM6Ka6
XLTAD7yff6HaCebKm6JLTtMoiFpGVNondJpnqdO8gG1JH67eJfHeXraGf1MJPz4bZltp4rHB2lxF
mOVMWtTj6qkM/gY6xIRSElkijUIfLNquHaUkymzrZ2Ku6Oev7TDy5EUF7y8xU/0WIGOp6rd7OLxT
gKUGLsW0wtrOQ6/txvtj4lZ7ddxE8L/vsRrvGqN8fCgws7MdX11u+Jmm/0IA7fsXr0dDb+dKqxy3
XSIBSPNapmg0SY12OTivYX+Y6VJ0jONDgg4iyCdY61/MkCQHhs6FuA4DwEQbX5x4S4mcvvCmip9X
cBFYxDfXi1pF7otnwFdVIbfnWGn48zDeeInmw3mI0VbyxPVsBLCPVDQKt0OCW2BH/xpbgtAICHmI
MfVZmR2RNhL/OHHpt0tC3p8TGHrbT//wk/jyr9bm8KUKn3xJozTIVTTzB3S6uSQbaKpA/GYGm9Ly
jDWzjkDXAIVAZ2a3T942ERlTy/v7Es6JtNCcbCRvaE8wA653r/NkunCMbyH+6FExgQGLwEiu7TEQ
DzQnslv3dO/aTHEuN7plgQ27hlUIrQC0mGHCB3D76pb8L1eNSq3kRK88LWbGGwsQ4LWkPqDr9+Lo
KMgr0MuoQLFR8CvzrUwq/yWTFvyYKDETV/OaqI5o58Ig9EzULJEoarfxLYcDak1cGvp7hx3/HBIA
Y8KHEKdy4JJMGkIrDtFTknV9HjhFBlHYae/bzK6QuCWWF4SdiN5uPVydjMwZVwSG8SX72O2HA/4i
n8padpmrgAg9LuLqQFQFF4f9nb+6ote63HDQzdVixK2rhGUYC3yA0f9kwMLOh/wZ5B1D+GtY5d/5
1GR17FkQU/xg1DMNiOzni/TQ0AkNyDhHSfvFiJVn5h41a57Wlp5HShtcttGV2lpdI+aJ+r/VBvZU
OTl4I4yJz/BfKGVZOS+vHXj7hbuAIQIcosrdOqJwr6Ybopl8MY1/iECrhMkL4IzCe4HOTnuekhAJ
74/vNh7Esrn/YOaunBNal8w7rWgAzZgO3OC69vz5CvX1HX926iKl5zB/qVhrwehwIMrvVAPHaQBz
MH6IpHPqeyMYcrh88YhnhUIHB3XGk2D+o1NQKu72kGXUcAT+UW6YQyGgDgINQtPtfWZVmYkGS/TR
MiuK7kN3NFF3qoOF3syWY95sQS4tz5j+AnGAD80dreu+SE3oY5sAJTaXeeNWN5aXtOSbq/CyYBHb
sUCI1MApNCV9jfbostNNq2y5960yp6CCQJzhqVkiV3uGHddKlSfNf69Alj2l7zyd1TbtK5IHYdjP
tXmKZq8W1iKde60gj1qe/sc+MOxUlsngqs7m9E6JFjlfpJ+SHvc8S187JYzdRhCBhndMqfm3kCd1
/sDi7PnGPiVKR2LW5RV/H8LEc5NK6J7iBjshs4dcHfiDcDcyVY23vIBVNpg3qybAo4C3X8Thn3Eh
8wONibmMbmA8R+Uij/157haOPmLVJmVGQzgpOw84HefcdaDV2SCrRiJaiOkSakc7wnVraKHKg+yV
tIMG4KPkp/iNInm38lsEB2yRTWSCrQ1IQ92NV5+p6zi0IH5u0oqtUNZpqkG8gZZN15yDTl1aLJym
JL3PAcfARyerjWHFchsyrYlkSNKKGxvLkezyDbkteOzcez5h4QMLqkJFbcNxUO3bldRV69nhLYfa
y6SNhCxxg1xd8rnVMkMePfbpzNBO/rRG56lgcjdfjK1qekF2GC4GTcMJBZqIQtPPwmoTi8/VijVe
eoR51AOP1KvLg0NQFIvgvSO4NDieYX5+BkZ7oQKL/nJ/25Nwzx0qna7Wp9fafXbIGsQz+oE7k921
4f608sJYf7ckYbcMARoA2HsMOQcdXVbyyROAJgXda+DZsukH95Ko5szp5HO2BKZcO8e9yuj5sAAF
U6X4zhzBTq/GB9Q4MhUoZgscw3sqNWgebLHxqXXg3TsgtajtjDv2aW733t1PSfkyP3Nvx/QLipd2
v7BzmLhprTW0CPRhsVUFamfICl3OlbQIwtZYMueB+D9zImGIhzxkfSSLT5gULqNPW+eKk0I8S5mj
rsuAAL7hRWbuNjpmQrDHkCe8DvGwsEE5InaXSP2yAgMkvjVlXA47EB9ZIPP4eOd9jkCd7PzODOix
ONJrbDGoGT0/UWl+na25PabwvTe3I6BphicuaZmpRAkAPEV+8268EPfWfCVWopbP7uQve9OVZEl+
rIcWrP2NADO4MxKCUF/1N34+nSe7U6vbibIwk0WFNc+d6pBht34VAn4b3AhbTi4KP102MjkW8ZYm
HsPiwcvBODrwwcL3D6ryPiBsQqlcINXokPSknml1CXjlxI4z9CKvE+E1RYLYxas1f2XlYXkgk0gV
ETqS0cHcIPDSPd46gzdQe7QEBdZ3TasumrOHM5b+kHSMrTsBFKzr/N5stOPNXX+803v/zKHwmd7F
1GqQhZLIbR44S5PsMaEdkzX3asGfYanMZFdVUp0S46y9fyrXHk6Fiv7ZVFZcPbX4O87d2v7eaBQk
JGlr78FJhAAI/K64rNfbubWHfgiHZtdkVyLcwaOEIqTiKNPRXak1tM/jWdiv05aEeZt65KoRgjo4
VUJdUGGmINDVL/slmNy6PI3h/BGKomNW9X70jbmjoRG3Cy+fOKoWPS0e2vsQrdYUUsUUFP7EDFbZ
KjlCvfOEqyC44Mm/bSgKBVQpykE465VpUJ+WfKgY72XCXqtT+FcbvWpuqYsWBGTOTzpZ8NJhKhkg
SctXfyDVppGuDKD+MfQB9cMiNmlP5H6aoOY+InOddIbR9Dun8pOPRLmjoCxt9qsc5Yb3lX0BgEyk
m+j+uMGdY6VPVJNt3TGxsGfD0wPGCF7ZuOTdhWlXGlG2hlSFg/gFPnlI19EgVxmQp9NpaiQ2fzUu
4oi03J/V+lbVaWA2/71mkpMXz9J0gkIcDVp3umwQOlRYxV39ER4izXi4GTdxcTi855tDVkmkjZvB
gykAhiQgAU5hMQqIcEbyfNScOeB/asiOux4VQGt7fGdrUDpkasB5NYTOL2IDvK8P5/cnSSIvLb+L
f9a0XRa5a7PKTp45n0NXDaLVo2myVEkeEaOa3aw6eAH2B+XaKlru2mjSKzTfUEKLa/Xbxgo6OxKZ
jFjZX45hoUQQk9p7vTUYwaOvoEMdLkcgcCmeWG8rhfG5NeVGduwe+bqoKZdv/LxhtfB9fRvKmkaI
hbSLRqWZ7/eEZ1YFVlFmnpnr3EGYoFqpK6y8p1UTzmEcEM3Goda2WYhORK/GogW8OX3YR0mATBk6
EB17suF1BGpKZri4/vrfqNrmHxe+RjwbnALhnF42qdjEM0W18mWYhq1QhZ5Bd8LDO0qtVRPpR5nS
xJKbnuYXa5qO984C9dnDk9OSyc8n/bAvNbf37p5BU0uYS7VmXb3ocehVmw/XJavN7pYhw57Hs/pZ
7nFDZCYUy+R/yNH1uxNPRSQJvQa8i4vgZb0+Y9DMgniFZWaTvIgvpm6ctw6hI34rxJNg71Xn4e9W
Whi3wJEWFOlxVzy4QkCe3gyH9hD+tthCwxszmI1TS1FBO3ZGkb6qr+kNWIPXr3OEgeNX5o4iFWpG
RcELz4U8rjqeNv7TbYc4l1gLdVZKepRNq6bMfnYcY3gypS1sURsxwKybMfNQphOnNP+uk/OPpao1
qR/SRpEZytKLRXryuVkHYkPfint6udqbbmuUV52VGfKkeMioV6NAw8eW6tSOH4BTADCO5ekMrwtH
r56iSMtvx2XnMBFbUHiQWXUJSRvJWX+t//PcDqDZyibFHNu/GUiCGjqxw1kkZIPbr5Rt4nmsDZEQ
5RWsrfDRi/wA4cSEaNPmZfgpfzIL/gdPi2oZ/ygxhWYEMYb+D5tDO5WyzQBnNWimSu80eMwKWosV
pxI8MKPBpfRbrJzzBElq9+zEBnJ6Jc575GR+/Kf1Dm3Gd6G/yDAkYagbSTxcbUE1zmdUNvwXR82I
4h1wQyu3JDI/FVtiafA8v+P5IXU1vouCK76ciyUzWvfbCaukxdRBoYg237oBMdQD1DMhdr9KMwU7
JVNFydIxEOmcMAa/C2nhhIkI7JsKm8ow5WOE2FIh/KlsS2e+rBpI4LtvTAQYHwmLgykkUxpKOgga
vEIzxkvu0SirwaMnFBUBMU37/aTQ0WnFyFB+O/rgHoI63mxP0kFhJqCmU3/ae9acD020oOfhgANP
Pi5xbxCheZzFyEBvwYV2AHadcqx2mAIrOnIobr8k4RQQvLrFwNO/WFsyueTndtFQNrJcHuHUppOL
mksv3aovnS9sXV3BVzP1dUNRl+5SyQgDBFwq8igbwF8unZyffUcDLHCuCaT01YbZIpl6fKXFtBla
fal5Ta+bQJ49cSd8S8OPyFM8rLKSTQlr/nTRjYkKZpjwc1e1kbPbaaSwPayNfR9FU6ugcu1v4WvM
UWLqSDgLAVDb5VqLT/D5Y1MaY/0EFO+gpCwOkby4ScUWGwsa75NdVUoHdeWVgjA1fqQL7WMa/qrB
mxx7V4ep8skgvs1xum2yeQMJYHgLSB9OH7xg0N1P3/XO55FqreGj5H2al9VUkVdW2CCWcbbfDlan
vcn0c14wPLgHlib5M99fRwXyXDKOEKJT74OuC29rI8u1fiHjI/Ao4h9mi6wM798+pOgbUwhNqSnw
TQzWUugaGb3DWui7l4t+drz7ydRS2wyRR1flIZZP42kMT2hoHPLfb6pm98MmLwWkEogQod1wes7M
Lj8Qo/wh4NSgK2cI1zxfUKjHrPJey/4s7Y9jnDefxhEqlfDsHOUQrvXo47tBBDUV2ZqY8nqVUhGt
KrMyEycMi7KhF/IFo5LmFYHoF0R+4W+cPMaoVYl/4lr6RWM5ue6uBM9E2Mb+F2weAhiMUVR9QmIi
Yc7DoUgTHqa/sIVsFyuAau7JUYeBvHszZ4+RitC0cq5CT5PL/e3U+MOD4s2vJRBfh81RODXe/Qp+
8CBe0qYczp1s31KQFHFNE8Qz1ZIb4RDSrmMrh9TRBTCzhSeNOUZlyCHJRlQNamghR66NpreXXKXP
jZMio7tXsIYHrxxU2BfpgIEpTS2rSgzH+/MECT0fqqWG1Ws65LmLOUbubvQ9pCdf++6xo5WZpWiw
sR5O0B/ROfvnfE4zpM9n0iZ1KEnG+qgFgQaccYnKDzq7kvI/A1TY9OkGjQ5ba6UQ62iIJJWIc6+y
PY5mkEyqgRJ3IVmHZKz0qdAwc/VmCeSGSPoOgiV2IV56ceMdbOTg+18K7F3YFCL5yQUahj2fsHPQ
BwN7mYlL85zSIR4tpBgjOFi68jzEo6ig+XJLHDemnxqz/vKbkDYyqUc6iHXKmhZQQvmaDxSX4iKA
sX4FvOsaezze7cFxxySPTFXOdl2JQk26iA/Ho2YzFxJxGbFZSXQUk+ZDn0hRtc34KfzLFYlnKkFs
S/4OZA61jW0G7QQO8xF3dhMjVXSelydZ3ElS/wEgpH7UXt5qQFENpgZAJCruC/WJ9sCSFz1rGxMH
NP1RgJUCoXQGlebZI3mVLFEGMR6sN7XxVqbiRuAJL5/QRj4jH7psXJwolen68HdQwaBq1RGf3iVX
DpQQmjLR2HB1sIYBXEmkHors90AkIrNbnsO9IScf5AA5xnFkA2Dk7Fr+veEdNXdAZsu87G3AbBc9
/dzzWClbknS4sFSC20ir4cI04R5g1Bj7eFwscumuFn5agD/LTMWrNRuzY8gjTcfSQnMFCwAUwlCZ
RpLqNl6Es9Wx8/PihjDnEhXlcX2M1eA723PT0dn7z0W458UxvKvEWCVnfp6dFKm+4kdFt2CzBJ6l
cgRNG7MYMarsdmSUxtVA1jy6gAoiGCeJ5GMFN9cWsENfSNJWyYguOPnFRuBTUBiEKRsPNmdjBy6p
IiEatqdpmS9ItVZi+M9p2ZBhJ1P+5zBi7a55rFlSHsBTNPM2R3mppWvNq88NVohSvrVIa6mXFrSD
rgb/VoRzM8NnuZVR++yFiYO6hGC/StsUBeXPut+YCknGsTglBLFnq8qaBnIrH8YxEuIiEyzJY3UD
50USNa3pNTW+JHpBvsGVsEpxcFd24coLOvitTEOazTmLYtZeWhbI5r32L2xzUONahuzPoFYzlYp8
e+IRYTh6c9QwtmK1Rg/xG4l0cG+0cTR+5TAv7Im7ruRAoV02xT3eDHL2Feyfp6OhaC5DbxPwA3eE
GOVHbCsnT9SyRSRyifXkd2vYVvtK/DudN78rd0/S5sOsyR//3TZLcVpTrg5mLcIn3QmYtHzmixpJ
uqibhBuTD+vGgi8NojnvPCKVT7v17lHCBk4YW7yALpSlr/C/BkI+hX82kCqUg65FGxAMVRs82iQT
xIbJgZuOfQxYbU7XxAHYkxPz6swJI74Qp7zMmOOB67Zq5V70dNLdvmi1LBkwIKsjwWSMFelUsUuw
uGNqav+uBy1WPapyGe+kyQdNlsp4/gvKxSX0nxnO5CgVbjJOCaS8I+q/O9InfrU0D+/nrYgAgLcm
enRo6wOoAqsjVGjDwtbZ3ZnzLac35W7G/rJKfIqC236p0HtCkLGeoEGIVSljUQp+5E9bbrM5i+ql
0MJyrCQ1eVlx10TeGGV7JPAWRVUGJlqxUgEvj0Fa4DZOwRfFF4bt64e30IHRd6PmzDb6RQ/lggpm
zdpaZy//jFUpFhHfTITtMNslMBvnjtVTAHP60k7k1tnBzKlZu5YemCoAoXOdGsBRR2AFOREhm6VU
ZCI58yPRJfjvO8hpw4t8LOKPPz01S2XLGT5c/Kt68lD9b2mR30p5YOusWd4UGboew661lTWfMsWj
G1SlUwkZ0xjGlRZJCdtsk4cRvawNTgxwabfz/4YCDGrzYKuXUdLGAB0BpC0iBg6vivZuJ3kBpNOm
36IT9bIowp93V5mpSo312AL2ZNbhcEfKI9jFAdi1ZUDYz5niYy5F7uAh3yV/yvMyblX0LX5C9LIK
o/v034HjNDXgYLaQJ238niFkhvpjhEJR6njLRmIKtq3MyfGOAN72NvW1FHkj4u1/NkLs7iH+Mud4
psX/r5ctnIHL0yrlqQ1v0vrjh329AoNdVzDOlJVzLtTlhkD7uerUA7RVvKCMx1+RFwh0lLBw+MUj
YCFpgou11VeGdDk5moHqDqjY6WaTmLAbmkZSYZgX9/EAYZNWQnXdcS0uUNRfLrFcSTypIS4uDO54
CAcE+nNEHnIxFh1wFC10YK7LmSFAUBkvE2o5hc+xQX0Up6YEBfFbTBl9sqB7F5qmtHQHHMBsSEq1
+yLy9oRhmzgvz1ZIWk+r81iulW/atvVwUv4sfd3cXgeFEna2Vvxaz3rirHZiLKp+72uorTuakwb9
mUeYIQkxHXC70Qrl68qlauh9ZFjNRe+1gzoYqc7ob2yrf/HGXHxtkryoH/F2bX7T4bBinRjNCNfX
D2xvlb679s7Ee49ef17do03/UpMTtSHt2zZKc5wYRsPyli/65deWZbtF4/hS3IAz9IJOd/c61AiG
HqIi1hwXkBjXFfwTvPmKm6Dx6kYHyklIlfgvFznx9axOrWL8C/abyqvQ8JZ40nEpDXcUDMjBqbDW
4sq4bM+Xo11ZuHyThwHv/yeTKtie6SJLnGwlZb4PdsTMQHQf3gbBvfHdXly0AvkjFsGfsFAWH+T0
vuMUeHP4Pw1sp0DwIK7k/cXAcvcsAI42e7rMAEe1dPBiX6GT9IaE1BJBjTUNHwS2Qn4VZPdrs1Wg
lNfcQ8tFaBHsGh0DeBv9fDjnZopQakQRsL3ina4NqT/MPt29QyvhhYp1L1INNhiRUrTo1j5nKKD5
nKdlkV8ft8QAYHPqp5OAhwJTrmGhBwTG5HgpTJHe5FnDS4LbvjCxz5pWZJ+OeVYpiDKZi4fK5c7c
YEZQ6t7WFZf181UBqjNkGRjxirlPj+777F6g07ZXwPjFK3vzpNJurSid75Q0Kw3AzHl+zUrLAXql
OjZqM7FuYsHO7H5OJMCzTL5lu9WDAQmEnkIXtPZABiakHTtWB54JGOdswV2x1ZWwm3CS3dc5oGg0
CzM21Eg46GhdF2tbZHNQuI+a02DuXbwhITkqE11zbKuvc3tQb3w/ZoCECAun9EfDbEXiwj1q/lzo
mLApkthyRWqQMZnITCmFanqjGkEhQUrlivpZ4leJ3Df9CUw/0GHDQroUQG3Wp2EqvO+/0gnmes30
xlwO9P8BEL4Ow4SnbU91VzttQad4xd3SmdYn+75noT4cJUYYtj+WI7BkI1htgehR7/eXfZJmALlQ
mYMZdb4YARDJbt6l8V+buZWrCzY86zBbxfCW6oSrWIzFrhzrBRyjyB4aydhiWyWhsUTEfNwgxLsW
UvbKbBa4PnC5VZj2JmCyP6QYdrBRBwv13Lu+MbTg2XuGYK+/DdUXbZPGJuFnZwx0AUrELSPktlL5
KuoGzVqMwMF5plQp1utRJMeqqOt2XuNjKXKWYWth8w2JphCcOpNmokrXp+B7QBj6fUqFxKpS4tx8
5uaaxWrclXkPNyVrcqcv73HveB9eB+HpxWE9u1HmCfXWot/bPL+EvbkHneHQJasLyCrmzyASgn/V
ry9cUiv0ynxI8U04w4KWi3eSaOnoELZTjvH/RjP14iX0K726ZyM8jaZbK06eUijeMqQgWJL1O8eT
cVzHRKyIwpO9EWL51RrlBSXliYYNvjuMGyecFQvK6l434vCeomhducoazVcuYUZ3ob4vl8ZX+p9b
gKmTIkXDuUMA4DYA1QlJ7Lah3biyg0B7kA1yvfjaNKf70ihT3ID31waJF4E4hfr7GfnFLErN4cgL
CZHG5V07Gbq1tiONf2lhvICSpTb/QnnB1vKBVD/RrGvXi4+qLD8ZBXkVPaYIazENJsxXgb6uCRTa
SPNCDkJJruBuGs1iUTnn0iF83imJFg+lEF5UNhI4u/6U7pSDx+vCtgRpf6fy3zHr5HzhtJ/yp+hH
Dc6BL/JgAsNG1DC0evr6tcRSypZuevv2RkBRcAhf+na6dYCnQzKfJOMO7hq7CTwi4xHaXIpdpW0x
m8ELC5JzCMomTf8bQOJpyyyOHNSIGGAWDZBHeU71bcA5RTfzgsLU975Xox3448HUMbJH4AtZaHFH
g49jUUWAlCYo3/MnypKQLsQAMPNdyt9Kr50HPTd3y59Nb7CalIUFVAWkAZawMFK6wHlIxoPuivRM
CY8jOZ08EMrlyiEvxb3Sj8B7KROkeuKaouqUo1IcdZKbouSbKel+hAWG8NmwMFyTbDH0lyhrtp0m
enna7Td1VZaiygr2g2Cj0GmCz3BrrnLq8FcPdd3EH8ua366IHggBNDCK2rLKrCNy8nUuel+mKjQ5
TPEXzmKIVYSTrOId10gLBL0eflZuMPGjkn42TZMT+BoNRiEGPJ5ABC2rBbPizSCggOCvqwnBZX6l
MDSQj+pj4rvV1i3dsiKBw+C9lsDfJ5KC3xzAY8eJhqvaCJoAYARA2t3h8qhFEcfHsAxlifGmMmBH
gY42OPmJEiL6S0/i61BQ4RZ4IicCXj75ioWIrzTpvOZv/Y6asTaP8B0DAWrC7N0iowA7deLv8Ghu
A3tHjkRvaez1e3H8UxdUjUQHDTB3LlASI+nrKdR5eIRz3gB3WClwpESIlQGAbngJR+tYJoD7yjaQ
LDkeNulfqj+zlIS+nDdwj7GaQm6wdGF1eNLSmW+5YiLv+pCknrlmJSgf8gG0I2T10srGx0eT2fC5
smIdXMDNRjS8wf1ZnD3ZVn8lw3m9QAS/1nQayMCf0r7wg0UcnBZzpqPH/+KRFxH69SNEo1S7iFaO
/+K3PSjqjCBeX1hJr6sp4kXxGTkaKv2etwYONwRcIwWghhrgAUVqX2nnLGDFVGmBGsoCiDDviWEv
PgFko4ky+XFMU0n91HYnPZHI5HB15z3B3xgtBsmg70c+iYdTbRS2lUABFBvgAOiayzpMCnQaCJmh
teWJeQoK5g+nu7a5iy0E0kpG/ZQgc3HDhaMJFKGSwrR+GCG+7j2tNPq8H2k4nv+lFs7Y8i8sMOCz
xGF/mqOkKt2njqMY/grWnSDnFHG0HwpVKMpSTzlk52c3MUQZThCtsX2mm015q3gtlmB+v9Y94ujY
UTn0+rk8k9dJYKWSWKPsOz91wPvpJMPOUntogjO9BiENaAyGMCpsGfSE4dcLIHbNm10mVHMDEmor
7WYu21YJDGIabHvRyJDoc12F/UabU5Xey76x3GuljVqLXYuAAMVdcUxz2F76HUXgH3hri6Q1yoDU
r1g9r13aObkT13csTKu+bBnN7j1rcjgOgymebd5ylnyfEr+BO8QnHF8IGWlaVO5O5Cxgvofn1ZMN
9jZ70PQ/TPQYxPmI3OjPLY1dAq4kSz5briT1QMdBc0Wk5NXFtEaFI0yvX9i4bgAwctnMxW3YU08Z
1pQ8jpFcd15JdOB2Xj1CFhmkoTwk8WcckN+a0FIud8hAZMVlglVf7r9iLCQjBBnHg0CwOfPLY718
tUdR4lQI7FwOjHX/309Tq+JSZxzocADhxb1ojiK1+uFRTg3A7KWuqka0hIDzBadDUK0qOFxRJuZv
u9F5DvyNi3fIEvzzQ2hy1UzZCZV1XibIxAzeqNI/KFug9EsIyXIa1KxvqkMcry8m8/UdwQRSCXco
NjM68cHB/dkm4FjCDXxNX6bzVQ52E87tyzKRtp0I2R808v8XlIQkQhHQqfJleCEOxk2JCIFCc0H0
KlGslWqHFzHBYVk8LLK5XMYG8i408yyNm8/D6k9V6jLJTi/RSxsCLuEwk1vhgnhzaqv7GZ86Izin
iDTW/FK+GxjQidhPMnG9mIq5LjpbZSMgJ/X/fQSjKzeAVC2SP9tpzpeeE6UUJhfPVe/Ea5a+zmX7
giFCz9wxsHlvRBfLxxk2A5V+VpSZK/RdbWNztmhx5g6hLdCl5yUK92ndFE95pkGg/Cmw4bn1MuT5
WHyewN0IHtscdyHr0ssXfScxWreIOWmnq1Uwxxi5ysXWrwvP8OP5NZx31heL6WmUOKtIGDslL+5s
BfWYks6NcRIppyQcnGfb8QdnJyF5HtiaRX5NDQty3PlFBkwdxcLHrsIWe9gLAZaBh4fW5sjGrdsJ
8hXmJRGMD+ggjvK1gimK4HyTNNSB/l454A0Z3vsMVdMtvsphb2wO/T3hPWoFww3CRyoUnJfvtmZU
hrxJUIzxOwB9rwEpf9F3x+zYVNs41rdA+Tgva0nUei29crRGqjnn0eXTIdI+I+iBpWqhHKzID+SE
KblLDb8Vtve0lnb3eBpehtLCDit3HiThx0qR8fWj0RDHxDisSqhe4gHQT12IBU2TGO2vwB2noGBP
7sRjRMpvk8lbqlwWYE1eQCnBD+SnxE7cZKsT6+Vsz0MUxs8VVCFqhCg9ujBVpx9uhtka6f3SAroD
CQ1ZeQg6kiaHWauKqcMJVshj9p4hN4nAl9L9bFC8Bt9xh92cWRzp8d0MJoOuRVNwBmRK9h1NN9fl
mPO1Vz8SHqZbg1ZIh+wASgBj7FFqI5hmSevSFiroGZ2iCe7f/JUPI2fPYfX554RTCWpoNiAF85nU
nmjhKlSS5vDuTGIljfqheervOdhCCI1LE9M704IB62cNtJubjUzAQKJD3hBOXoV9vj3t/uHokVi+
LYvVPtb4tvXzSrlETbt144ImndPAI8i/TzhRgSQan4/i24kkWFcDxqvXdMwcc5PjFLZOBoFSzWNT
j7r/YhWqus3iBgflytmho68o07WtBY4zuA33rl+PDQQkULW34hnBIR7XfKL37apzXjFz6q2HVysT
VEitXqYjmRUMpxKLJ7o16VRdw6ByHzecp5PLOspYl3X4jCC3Y+F1Zh+xwfsJlfvggHE3dBUxambQ
hA9wkcxS3fPD41c0Wq+pcM0owmHlXnOyyQKl0ZkdGdKOIaDZ6Oyx9CJSv2rBkVTIefgonEdblRT3
QhzpXVRFHub3KHUQeVWUJJPOpXGNqWfvxn2eSXfnObxl2gAYxMh6Dc4a9OvAZHhOwVcxuZrAw2ED
OYZihuHP+MXeJv2Ni+ddUybv3J2vNzpzXtBcyHp0fUblEBfOlN9ASB2UG739tN/lcBfGdP1tXhJP
to3hKU6jM0wWxJ2V51e449LfZHMNix8HQvT2sAeub7fahqX8J3j8m6Qk9fvVS9uVhkUeWfMy9Z3q
N8K3yYMwAKamVRoaEC8MI1yBcUHEhEXMdCWt2oLQPLNjp51PWQtrsQF5/Hu0NodLELeEeNdsomlt
xN4VYXvqBmpBFICLpjlEYhb5eAU63+I4S6frY+9KFxkU9Aqo90XQM3hh/qEOJ0hXMyY1QnxIwrND
Gs6T5qXbKzjMwf98qdlg2+NvnyEgSN3eB0IvMUdAbsJ+3UdDL01jb+qx4GPuo4WooW9nuZ6/Bl6F
mxm0wuorVlmloWKkjwtTHoTi9arC7aEaX7E8qRH3e2TXcis0inc8f3d6E92bUzlda+LVuFeA48pT
4vnK7RZubuVTvs/0t7E+/vUgL8oUKBaiuuyRDz2CLZHFDtuefldPpdilrpahf6Z89CI1wMPuK2U/
0Wbtfs7kmMh1ivy50IgeRmWAiZTk0VXQ3OJiyxBo4Evns/4uAsu5XFGmGWv4pWuxuhvSRUbGO9IN
sqzYKzZq7sjPSzoAOzX+89edRqm4KiT5x1qcNUcZQUV6f1gqBC8xaOIB3kuLv3YVKM//Bl3j5udE
CrDdDdfxCtd+qJGYOmNen/qa5gfQMD38uNqgoY5H53usba44escCNkL4B/vazsfWwGFWosB1p1vA
q8t5wB0xRRY4WDwynzs44lkofY5K9R6fu3AfeQhPVwJeLisl5ZZcHc+S4oJ7C3GQuTmngYrt2qEm
j+fingyeOePpMKyLryzSrWpfVHyB7mQvKJbOrzrEndIOMn2NWlZWMVc/p43MFwuHCOiYgKi88oWa
DDDWjfKXHGnQBdoGpdwzCgfhutlTM194OWo5xyid8zPLhcZzrxIvbL6oyJpXQ1DSVIk0r7HA2x0X
eNSlJXx9/KndaY8AhrqEr7YC+q1hTeb0282ABAyccDOxsLIckBeYv7sIboQLoo6QqJMHCzxleW5Q
y9iONsWugNmCf5W+PPNAwmL4xzTUSWDv/82t52xSGiv/s3aauxIjp6EhR0UVoDwkKM0I/LZgVh24
arXmCIN0VGJuEcy/oCXfXIQiemxnIZNi8k51GKEbcA5TS7Ati3JyatFmMPKcrQoXdXPAuLhcyJWz
qSCUPvyRVG1bQg1KxSZ5dUqT190WTiXGt3YDMu1M5aVVokcK6KCj/zF6EvGSS3vqFTvPZ7u5vtzB
K9nBRXOhxFAntKijT+quq6n5LeJd7Us9UB8kFAoQ5GqtWIHUxkUI/UrfvA/ph6WzsNQKqBmUjc92
+RZBlCI77N86kYs8lDoS3UWwuEsaQiYGPYvsnufBBQYJ2Ezi+viLc1tNl378daisPSPFaTRiHhyU
uNQaEnmAuAB42kTyK5ChD4sgHYAjKONIgqSLjRnRSWMuHJc+G8M0HARzdnoINdcZuI9pV4eiAp7k
JPV8PVt8Q4pB35y0V4mQOd6toEHyqiAZwyW8I6KrIXDW2KiGYG60NMLC9zZGN49WuHKg1o2R7fP7
4DbrUIyBxMkYsALJjx4jG/tviqGdr5oJ+PJfhmuKX0F77xTjhdHRPsidOmE2i1soPgnNtDV4K6lI
dmPH++XTYCmvWgExEphwiSvP5b++WYtpdgS+uB9jfcXrL1B/HH7Go8tlk/mBF1mvgaRjhkQeXAMz
ZoJDhZ+Eied2M/mgYlI2bUuj/CKfg+udz03YJbRn13scSrHii+XxYsspSKou65BOVwmhIV0Lrlzf
65q0lOZUg0eYU85xTgsz/htOSqTlb1IxakAGygSfLDpNyVxzAtFQspz9fXhwQbg0J4R8C/VsYs01
F9Nd9cJo6hVEf7+oedhU/uRqJABq3IHdjddRU8xWp9REbDh6BWJwCpqjGZUtE00tUN1wzvnvdvAs
pZ4Lc/m6AFpr3o0/PKZbCnxj/dmcLDXGXXKsEoVPEajs1xS5G5M686n+QLHCufrOfTkZL3UrzVjs
kr8yK1MwWEVCh6PXpyDAmQtEL4+l9hNvrw4PjPRbN9VQzEDI0Vlp2WUrrz4n0AZhqGde0rfwrFMQ
7HP3qOSpLudGqj3jpAqIY/h9NCbfjg6J0SBNOu9aNLPg2Ed4iq12AcNhsbcbQJnS51k8G+FOAE5e
6vL+MAbUSdxLau3j/i3y2Je12/66H3a4OZWgbv0blliDMqx2J5uKCO/juc3Eu9UAgesr7ksdfQkU
xQbJAX2GgHr4eD+aDke8A2pY1pt7exRqtpCMdvOXxzCyRMnZbDXbljwC+7248UuiuU2VAcjR024i
9XSe9AlSnWKP/Savt+yaCHcRb/Vh7DSTcSZvCQcqdfow1xyW72lQxcw8hzYGcC7ppd8fwr4zs98P
wpebK4896Mlt52A43AL4OzfqfLvL52P9+zlh6Nxr1apwCKVhy2jQxpPjQij+E7+GkYaczercFhPn
UltEluhU8GRAxYsXJe6TlVype6+dq9fhvODib5XWZJIz+m+stBkYTOWJOADfT4OrpQzFYx57bsBS
8CF2ZWLfvYRk20qgqEtk3FZmOCwfjOEQ4865/A/vZyFA2JamucZC5WEB01J51gw4V5gV0M+yZdFG
btYJq/EHK7GzOguflOIZjpkFtEScK112t5pMnhPz4ypK2BeH80PYhZtun6TiFrwip7C2oNYcp+a6
RetjXY818od+dy3DqRHn2EX99311vqXdRwICm9gw/xdZhp/NnvH7jsvghZbL9wvCiNI4cP/6BKL6
uJsVcbHqUxttlBtu/6Fnijd2WbpZuLcVEyz/ASYQ/Db5K7F8MytIdtv/qyz+dspadbMJ6ZqY8Zri
y1KczhBqKHwqMJtPvh7AVjgDguISKJcY8X0ZTLi+xkXT/ByVN3MTBGRTLKnnmHOiZ1qOxCqKAa9c
LuLbZy1Bw1xOl10zLKk8FYboHeV+9AsDtAWAqEin0Xf/SfUhV2Bwib3zZ/hALvmb6oeX5M/YuupH
lUdm60hYuZZHjt77VJy3dR6WoI/iSSJEf3JpoAUpO7JPMyislMC/LEw8NWnE8DiZiwyLCBLMXvqX
xbLkCSN7gHaODiROSG0kYkeEu/Waiu7EKYRvm2nIyz+H0Jch8H3Q/PvljQdcI07oPUB7FcZ11Rbz
sVCsfO9XbSph2xUPh+4SvH9hNPwdqO3SXmjQAncrzM+lR+e3NhZDAY0LXjrigxcH/TAOcYQuOu8x
po0e61OTQ71PnHauNIBKks/61AJ7gZGVQfv43vs/MKqKqXT7VOGUGpNziDGeur+2t4hL8RdxCdwd
wiG4YQYkvniWpq4D1Ycl/kpiErt1LN6HOt6rTEf+iuXWeqrGo9jOGG2XN7+y3cjNqpOXNr1joVxd
0OxoCIq1M5hT5Az4P3kIzA1UDup3euRmJUa9aCVHrUYo77KjQ4RY2D0VBXEE8RkIxN2MKrtrW8xA
ME+ovqiK2QbIB6/kYk/AmapIXRaj+4DtOCA1WJyghhK0x3vPu6D/FrYpveHnj01uydzO10+ypOOX
WqsGgWjZh4ujWChzutkS039xy1m0nQdPnJ4ZlcwJUxMSngTvQJ6buu/uKrdsbdIsWSKuwa6CJGZ3
dWHSiZvX4SPcJOnP5gX6dDeI8sWcEmJ022w3FPwLGXitDyqwIgY+kYjdVYBbqAF3nNlXAezugJgF
+lp23QPHe5/xM9ABhfUd2QbbjjG/aMRIxwwi3SU3GN7et3a48RXhP5z6WwqNI97bitnMPaeJaS2X
5fz685wn7LfnwW3NEXVaXIE7ltV7nHikiMzwEZWdpHs02tpCGJt3MidMYpAkmQZUYrAR03W6PH25
WN7nFOacdCfwqpj2HrsGFf0Xwd5bzzJzSMsvAKSvh+Pl+VBw4VO1qdaDEEsra6F/FN4CNDkxiVmw
pVDPhZtde/UDM3ypx7MBlVXYNP3m/2mJyupL+xy+JXAMu6I7oRAR/XDHtVr4o0Ff3pgSljga1Own
z7wAalUNGm/2kDZVjwa4ARHYcB0yb9bBdyuw7BVqkKiZjx+vYkesYJ9OvqgkiM8ZNPQYC1GVsZRI
mywvdLS4AEYHoaTKb3U6gbei4mScUkQJ6z5TiTHsWOub31RewrqXMjik+Ti/AD6gGUnriEBBOjIT
ZKbDDkXUKRia/nTg8b0XesE9V0GdrzOsfq0alVJC60+sp2Kl3qIu4oXgkEmRNz6N6xvxmOsGRv+e
rpJ+Zfadz146/ojmzGv12Z2sUXlQUzTCQAwh0kXrZustQ865sbk4Lmb+XPE4XSmgwyWVH6REe/j+
95Wv689uzmT2hrTV3EvlAdkL3mqIXfkmt86JAXPJCsamUpUnMO/Vwo29D6RWyxZ+aRqySDaJFh5Z
wuwUpxoNn9cdnE7D3XjC5Nkja9ywYdbApoCRsHauPx+xHfzT5cNf6yy431rdVzyZiHZJTyw9l62Y
VoapruW45ix8OTGy/9GEEHYV+L431ThMRs5PtnVukgZIS3nRTXSiRL4f6WwsrnYuNf9s2Vustdt9
RtaQt6yog33ewGhLe6ucu1rdE8VblhYdvDQRJD280Nwk78qYLjHaAmuZD0Khhpdh6nPKvJEgPmul
Z8pQRlynQG6htqxtlMnYwMcuwN0MuyIS8Bj4XfxPee0Tra8WLqrsgIighSn4FcqyQL2xDhwYnvx4
faxjoNEDZLT9OyrO0efvt3mv6hpX0fThnp/kozEg/UValGcH0PIRAkWJk/fXXO+vqLiu8xfSoPy1
i0v6eJ1tJaHkgnGgXkLruXekYwT1NdjBJTIfy1IX7eAdE0zwqGw+UQCd9R5i0Io4KKS108QWorkJ
ZMX01qD99F00lgKCIaC9HRlgF5sQdbmyFkTnIV6uH9ATqEN8mdhC4a8B/xcgjOdzSr4mmIKGr9tb
kjljDqO/lGuCWg5ZQjCZUW6PvL411SF39dAL6sd1t3x38OPofZDtpwHEKGc5NIbjxCfvRTt3nkkP
yiXPh7TmQwui97Qbyz2FZILqcSDwXeL9y8h9JBb0xgjaIHsg6QnJG4lJuJaXUu0b1QHaFwwpMcZR
TUMXHwfkMqpmsCbyuMKt2uAQpNu4ouj0gJrc53+uVvE0B4LQR3WPTuBYhM9pq/hPRS18YF7E+Mr8
ZWFIUQfXakokZ0d9Rk3jm9IXfap1ThmgP+uZ9CqoTlY9wR9coS3w2C5QwUkuOEfNXxa0rsNV5V7q
S7No4dRgeb3ZxE9K7Ul6NwCViynTip0vjUOlbuYWS1N9M9Ccz9RtLlq6LyWZXdvnQTwvnF7nn3nJ
AzgnBTKYhvyMX6OfB3yhrlJkoknGzPH6V9ISj2ZHDIqD/o2I4Y1p1+hGAHccgK/BYn8YD+kIGiVx
9Tc8jXpHjtO9NxGUi1B+EcAxAIJfjzlD/hkzwcyucnIIwLUGoJHmkiEcL/Yt1uw7GxgqMzBB1d/p
oZfcVEuFp32k8Om/tscbFJmOO3lyVdW1d3laLEjY3HRim+y8aamtIpk+adRhWaoLJq6JM/XRfuFq
jB2qtQKgZTll1qv6T4/SkEGGkl8/j55kBBZgXrayyYWjBuEseyZoREP4wmirYEnYJ8emYhKaTUfu
pcXMVfwpwLmG6+1beluz9AHtXvevipxa1HTrdzqKlAXsmPqOtzi3xMayvTNhVPJid7/EqQlzQrYX
B+e/B5ttaiET4/27AwiQLk6nYjCZmtaohofgQqXvl0X7r+l7tBjUFNBCCq6XSfUqx3UGqJV5pRZb
Ba5LsHz/L/hesI0kgjwoCqPC2/9L8rKKGKnpsnuv5KQGOpmCX6OSr5TWfpufbOe7SxtfpstUTleE
Ycm5vNJzJpcDF9BAsc7H7jqsSj49V6DiJ61Yu9zAErbahC6NhsSqu8xdKIpnLt/qdwe7+G21JniH
RGv7wxZxqZ7M5BqfN5Tfg6rVpA2z5p/NaYsIGhYO2X7KFMQDxAYcvwpB0Hri7VE+6UDRP7sMMUGb
nD2Wrjl/ynTBBKDk4qm12/lNSc3isVdMMhqBO3yr77qaj9o/yxzhgvO0JUz0f3StmuNy65mNIYaJ
h3qzkdc7idw68EC7PbaYmuWhAMtNJBnLM80bQw2HXkD+S00ulijx86LwShrATRPS68xTIQFP16oO
oVm2dypmjC3jri3NCCna11BrJc2suLcTSKHTI0ZxJQanx/lY31XjIsXCsauAMEJN4HMmeBou0TCG
CV1eA4zEUh5jnpn9KDVrzEriYH1U32NAEEl3vF8/xqHiuSpXcz+IATcMeQBFWaB2Wp4NjOTuS5iC
dTqkTU7ndRqOK4o+dP1CprrW47cJo3+KqvEXx+pBFflxIJ5VEDyBAdulZY5s+V1A2HWLhsWnVcjP
5+heEbHv2nRv7XNCxXbzDtS6oPfZesr0Zq9eHbAPFIAvJ/9X9EEpLWIhf+DY/x4oi3424f45wAGK
gIIZouAcvusf8L3QIF6XAdRUavzSkEf5U+hvJ4ktK2ESsbzyffyCcrJJMnUwwJ+iuZPE0I/o5KVD
uz+DfvUlO4ddXohMtJTVk01gXP9uViUzkBPJkN1c6bzuZfvqeFBi/ojGBY+KjXJQI3b2XnSGT6WB
I0RpwMiWxoS0XzIl2IVEslUXZooKjPhYAjXcLje87Pn87h9zjirn+CCiE962ghdRVaYjsJFZ9H7S
/UAuABlPpxkA+nM5U8misY0bbJ/VD3w2AOCiEoWGslu28fy54SHklVfC6mtF69nDLg+Zny1jxgg1
ucaQ/KGP/eyYo3Yh9lSYp1vGvUjpydkQihI6+MBW+RBs/SML81bGHD/a/wq/ri7YM7WCYUmDyOqw
X0nASf4hPD0bEekJxmVC19z4WSGOFoLPsMMbxUfTVZcu38d7Wx6UdYncsPLLdAFdu29a15yt/QDz
vK2vUOsbYJI0d1c04PDQjyHt54vNU8jCRaEApsSgH2QP58ikDnqi+muQxkZ1ixan0csAgrJZ+SNV
bKd6DCgmweMB1ME8vgNRvWThqm60DUetvEn7LLptzQE5Ef1L2Z2nCJZTb1meX4hOgTvc8pIpJl9u
bv0VNYU31DWRtdQMvYepsSJOB+WFDneJor51vCT/QDptiWayVOx4iwkB7jr52GwA8X2EhHZ9C7Qy
9JoWPYf+pfRO/wTxbkPuTQ78iZ4ddADL/uagt5k5ELp5RAmJDFIdHZhtr06Na7k2R7M8e6ZaxOSk
8C6J8DS2IO30aH31qYczG5o1j/0eexj+ZJAuhMxoXYtVGx/PmDke2WVTIKGeu85sLraBP1hoafe0
dv0k/kmXsTXtxBkPumD1KASMYz5F/QpYA2T2msjuKS0z0HkdLhVcvEaTp4dXS+NM9ijSPMED5310
4nldxyZGJMCZkrRqlYXFZlHLkQkTA+87jUVDwbt2dmVJ6nWUTeodJ2+7WaUKJe/v9Qt8Nuxfhww9
rj5EU5njHshGMFuUs49sosUm0sPaAFKNhvGgKODclXYsbYgTRh5rh8eemfyBFiFQ1VtEmmopOCY4
7iIA3nE8yvdZtG34PL26XPIzmZA4FEgkPlX9A1nyJ8Ynu8KsOAoBAU2eGMirxsNu7npF+36Zv08Z
qLUk/4lms1w2ruCbt59z8hfO3boIqQyr1itWuShPvSjb1FxTTY84q5hIMLRPd9geEPcNnhwVzdnZ
DlqH65XIgAJCVDR1z/WDYdbY7ObLN93qzVLBSdflo5zBsahgV6MXqsLp82ZzdrGbCGmCmfMAZIdB
L1m2P/Peh6rrUwAnaAJjZTmvRXLCyMYYGcokqhbdicSOYSWcjqD20qQuq+EaDn+Bnz+ryATFRsOp
7Byrj2uBwWD7+C3NtqecgdGGju7H/TmZsbs+W0zwmGgjU/qOEEv0MM0mkYFkdpy8a8nf4CpUOgXW
WREXpifslKTyH8fumqj3tT0xJIFPz64OOJjQ9NuVIz8GKeCpSEp83wX+JCkj1acHcvjC7IZjMVGk
sACj/ZwoJuc++7TorkWY8S8qd6K1BHSCpmuUMsgGc8w0m/LWpnZG5Q2t3FZOCN3627F+4ogDMXrn
kSZ9s5lx8WqhhXrQlTySwP4xCsukTKGaLk4ZRQZ8Vdsm2fZQm1ASs6EzotN7LNDdkPoVzdJjBpf7
WKEfvsKCvrVMuIRFZJXM7FLKopRGRW/myyISr/8P45BfhuFlimeVudJ+1FCZUBBQMGRtm8qUuJ1n
bbG579EL5fnl3EvLKdb2vXY9tyhMPUSvVHkcdkXSOSQL7ybnG7EtZBbbGpB97K/j9yMOIDiDIMqm
fHnZwrWhA4JOhJ71PUppLGISAJRa48O/gCZHOE2zMAMkarz1Sel3lKNp0WAswWg3VuLpUODtutEP
bq98H7/AM7Ra9LCphdSUYOExItid+C7ssV4r5Xrw5QImd/jHJv2NZ9IEtOP67vHau26UkAuqRSiz
wTWtcCJIVNRpDIaNFfr33WhJn60mwYskMw/YkQ5CalZoGwDT8T4XCP/DO3hr5bWTLWEgQnQpYJQV
QloWVKdclYV4sSBayvul+K5JtURtpLo+oj/RVUc51ORMvqALGzqw1phrgtPEzBUiTTHP8yjZHORr
1On/etQpUXCkWQyiLSPniocmNvaEj9l+Ptgw6iaDpgEywCCTNj+zP9H4D0POi00g/XcOtIG3ubmC
BFMwvX+P24pc74fKDOmDT0ANSneYL22M3WaTFDc8AkUHcJCWqbpd3jncD5+PeLPF+4nLvR08Paha
Si/LZ5oo7FnNoAMe1H7G5cH7jpFv7AHTjpFQCpmfIKLCgJzw2qXdxb1zFJyItSJwLACiqEAjNdPw
g+Vc9N3Wyk3UvvFxRYWLtb9O365L8x6WI/4jB+G/MiPG4fZiA2uIkxwtS7Pyx1ei3Zmt8OjZ4/1Y
vkq3mV5MkAf3Dktm4yLntctVEQgUBAJanZrsylHFehsUagE1UDjo/Bq5JiVYJpZLQZbOjFiCIWKO
11J7yArwDOkCq/Pig1gxe/hfGn+3mkkbL5HVmqOLyh8cUGR0WqPhO2icyfvsteQojZSzanh+5K6E
cSmrk7RlasRJXwQQKIDCmzSvBl9h8V8vM5uz9S9UYdFnhhb7Brb9zUIxiAbac58O8ecq4n51db+m
NWXPERe+vSMAwO7M70mB5NEP2OE5zfjHbR6DRrG6IJOKOELEb5xbOUXCCRPduXF+6Fmcky8DxHJ8
S8c7zkwvJ9NXzM4o2OKMTTDrjs3wmaW9Jyd5BotT3ry4f8JPnC1iMScLB2N2IE6hwArp9iziSZfU
z9GbBhN4mI2Dj5m6hxjL4Gu4+CJ3I8ElOaxvkzCJBpFJ5nViROgnIu1q6FHwmmu9k5Wu4SdPkkwS
5+8y0i09wx6xO874lCvaC7Bq+u+/39eiHF6QNNTnapwy9N8KHnMNu13qqqmsBC0Bj58dmno0Hohk
uoByexN1ghiLDneFSUXxWzjYF6IPG2Ncvqmt36sgtZmxRWhq/1k0GlTsz0fatABqwepIVQONfZXe
EfgrM+UnaT7Gy5EXL3FXkTLoFvTlvTMcpy4p2JZMb+HgRAzrLj2bMYrjYrdfXepmSYmuuxRrq+QE
WWaPB+T9duzpc+jDV+Xw1Vya/GdOKZRwVj4XP6Fo8KPf29nWsZAQ5pF4uc8upwdH8y1bJN1dXjqO
SG++ZwUCfGWCnv15hDHdr63tKUXbmdc+Qb5Ui+ZX7c/Z2dR2fwJdse6gQN0pqp9reG0tgpNIYUdv
gRXdug4W7d00FiwWrJJcMPCdwF0fblPJtJKSl0Nr7PP19cWnkFKKsGsXfKuVNEa8E03tyDoJh437
djVdJFicy8GxCFaIbg/u/nruSt49qQG+ubJsXpmq9RsKU4yoJZQHGwOfmgB+AS6vk8HW/LWJnC9S
9nloCULmBiPvP5qYif8aeUL+h+I/eQZwjzqdEfim8SZhydQ3mpXWc+pxfvO5YduBjHtmOB9fGzIy
E0y2G0/Rw4IfEPoKMR9RIOvF0JXi68MSq9pOvFcQ9X6Y1SvcEIfUOA1Zf59KQeqETVZCX17CD1OJ
fDeW1A7+Yo6v//PY2tMurkDIHST+1AxQal0ttyveptHmMSiHkONRGHQ0MyyQ+L47rZGg90TniDfF
pKu0bkkP7BczolrDnQnH62+GXJfuNmPLXW6s8kcY1leOgIXDcQQAtsVbzkYuYBkEsco+IEifj/F3
CLOPw1TlYS6U0VyMx7mo5yE8Dlavj5a8dxLdpN/0uxlBKeU/qk6Aea0xADj46lQMjj2ikVL7atwr
p9Qa93PgoJ6bKo8D7BaOJx7CW6Ekpr/gl/HyDmk6s8dFssyExDUogyl2gO7dA+GFO75/CH5eEn1p
G/ijjZYZtISZ/zI6FvdSZ4XtiJaXieRrkHgooboRFrS7cu8PEETrD+xCI6HMNQa4MPtwP9+muPYU
yquZJBCAm0iE1ZIs9fH7UmtmBLS7/M4tf6AXUmoKIcp2n/m3KOsDdLT4Ua5q5QAT/vwiM4dc1v3S
BxnD/w4ar3aL0RxYEw4v49z4FeJfFs7xvo1/ltNyIZBqAo7teTX1hrUCVA/TiA7RPkFkEDccit4w
VrbuQHZ6+fVSKTz81v3mK8x2JEdY6WmB+GW9pmUP6651zD5xCQFEgj6FGJA8PePN6JsgvYKiJy77
51zAIf4QJImnfZNm2KUdXgpcrmlCDfJcj225fraQtlVBLD3qooPm6y8qEsU4I5sTHxS/xoiUoeOA
Fn2NFdKvLJvmreoyvYxJFe+VpWcS+MflxBdUPOu20Nj1TwPphh3zu/oAnMW1rTWInKaZJKS5EuXl
BccHlvcnr+h4y8VqOUlrOFcUiXcd8yTVriDb9FS+nh0eXD02aqHUZ1ZpFLUccoPpGUJFERIKbQtb
KvA3BPVXKN8tYcpDA8AulcLRozeX97z+igpa9BRRaUipqPRwu6AGL2GWz+3oLcYYM24PeaYO/ZW2
QU6dpXbfC9xabIuh95Ds0W2VBaJEG4dDUQJ5YbGN5M5Ycd1akvZvWmNKgR13n8LyUz1um/g1inw/
bje4x4HswsDmld4wFYJ1ycADFH/7d7pdqIcEabLsbJzoKaY2rZnvOKqjRXFXJeIBbdNmelYCKyfc
zkOwo2z2vtvcl3jAgDPv57YtCKFvdWLwHpymt7pL4IhvSrWjqgD8uBXrZa+8YwDDoHyhf6XW5ciD
M/o6VNkAafcVdYmzoPoHaxZB4JAv+BsB7XpOUVx/q4neOvXSopnXpp/nrqO1LKF+2er/h2gkFU11
1w3xlY5S+7h7coTuJE4Z+A6/MP/tNNp0ECLPX2Teu57mavpVvAzaZxfUI5XJ+W/RZAou0Y+BZWEN
cJFUfeMwxChTt74o4QWHKZdoupKxb1C4q/m6mIy9SKQFtCk0oc2SQfGu+hpU409QFAxGzIIFTBKA
kKH2b0Rr8Q35g59x2uGOAlXhxv6tu7fhEIT4VlnqSbGMxHkA4LcDetshv9/TcUiyymMYnEjVpabE
oQTZo5NPkzoo1KDWEQNGU2xdYCJSh1cOwszAkAnp+MULeQBb8RgaEoLlt9oA5++wYQF1qSBjI994
w3mckdvvqrT4fp5Vweh6LIugbw2lyP5p89P+MX7rj7xRjxeRgcvBqzrEezqkJsQjpGToKbNWbqUx
qGROPYcX8ussYFJkVvq/Qj3dmlovbxoZyKABV8pRuuzS/9h0vZXN+OEfvnl2O6jPdnqNnPz9vnLp
zMbKfWgjJxtVQl82B1JqwHekNloZTe9/1E1dnpU82hOx+Pv/lT3MOujRNPRovpnVuCkIGXFtMEnJ
YpTnoMR9hQPjcZuz63hrMiSHpcrq0vi39XZXgcBZsbGiIYTcSzec9pkMVssLNfZQve09agHTKqbD
b3ud+glfUQVeDJUK5c1aEj9Wjsa3wC7n3zPSs17zxTL5vHbCac1HJSIawJZFj4a8gQSl0rD/7Thw
JIhbcW33O8RIasTD7XAZWDiFc7wcyWPAFEyawXEe1dlv6dnonbF/S+LdPLSPBUxd/TDJEsJn7arX
81cCp6UN5YZ9xoVLlKQBuVAX9RJDzam1Vt7Ke0d1skwfZPUp6KU38VvEA1nDI0R6QrfQCSJ6yTuc
SKjIMP7dsZOkCv42+OrzqYJOe6aZ2RkyddmnW+qziQ1GMh9m5AEOtKLJbqHeRnhpd/eAVkoc7753
8k8r+qVg9RP1teG+YO7ANU/HK54ztqqb1EsOIYLCdYk3QaxCVxs9k5dyK6UdVfmRu/CWq1buJ8yb
6z6CnuD5MOtO7N5noqERou3p3/0PieN3K0nVoepliApsMuOyLFrs3Oggp81ajzRYf5ZAAY1+299a
vlOXc7xVuaki7T30MupU/xL1M63wsgF4qAdJYzSguB8s/rnDjkWG5WMASFPAa5ESDBRfk66lVtKI
H84+TZ0E+dzoXzeUjcaK/Mh4aUAWCIJlKpGUL2J8FM4dZcbt86Wbdf7madIWkiDbP3/oWt7dzu5S
irZ9dxsw8Lrup3WphyTSR7B12rYxLrB1O1ZF21/TCKgh5a4eBbAdvBne44YKBkQYK1rxT5NbOPoQ
EAgxeJi5lZw0f8Ue6LxDBC1CZCqLY5BSbOrRRnSg4KFSYJostqIOVDCn0eR6B/4ju+ACfkZc8ZP8
j/TwQaCmeZ5CFYmvEp/DZ+Pou5j14+Axyz5oh1P/gp16t4gs3dYf5sYSv2FbWgCNWXU1hhpL1GV5
DJ/oks8v3I/6WGN1kjxfNOyf2mYhTnyIojkWj7qYp015XaoU3YkDHPkAhWoi+YjUl2bC7ImTdlOW
DxQIYq1RZ1E00IsBIRf3flIAjxwwo/Ry3IemNFnlyL9E0e2m6n8L7fo4wFICGPcxzulxniKPMzcc
+Q7i3g7IW1/mNQX/kde3bZs2ALN2GfvlncSa61DRTYVaZbztgLdT3hhcmcttEclzGYxX8i1tn0es
Ah6SHKgY0NVOqOjpvj8641+T1t2PM4O04nfN8+rTwe4FC/zJW4SoiCnF6zgHIFaj3GmjRk4siXWE
NL1guUkX50KgG8Nhf+9IDYRAQ8T9EqazeVuPWvEQgl6fy/+pvrbY4FppvXzJPT87FY6v9riIu+Lt
q4z64aweQ85aw7cgaO/rzryHPt4SFXJZyA8NLStq/808esSminysRa8fGlK0z2lIivIWqCy4a+ZE
D5uuv5ErvjkTd+stgrOFQ3B9wc+NUgNGqWhqexD1XUTqENw7DwOjt5uqyWUqOyf8NfKuiZzafv0M
bu3xWp0Bc8iWAkDmOhTbvo6+3+B5ZbSQ5tmYei0ykMhatZn5YGoLoWoWKu61jR/VIIcZN89jtqvU
DuHHc8/TWZxo09bl4UC81v8HfzUVwNTh1BP8gL1uA7WESrxMOY561gEVHUAEIRraKm/uaTBV1fhr
lr52rFo0jbdEAftZv6PiWH081YqfGonDBXcDQ97eCtHUmzrOUCbvcev4hdMmo8nmaZFK8Eh5r2Ql
wFKbAzPXVD6mrvOwTJRjCyB9gmlMif5RhWDlN/6Jue36bAe80Lh0nwUCIpcLL/yEZlLVVFQsW+FR
EXcvzKwLFs6EQb/ZSkPdoZ4xAlKRPGzdE6IVuKAbvlc19ZcIgnGwb0sHXyClPsiJvbR52K0yvbG7
/1wer2qTjOzzZ5ZfHL38LBk9101ZqcJPn06SS8ija3mmGGJbLuk1I+RtkD81vlahp+imSq7SHu7M
pw8/FItYWnWr6loA23peFmbKZAaiXhpv49NFqecn8cctinFHJWmh0rh3096dHmKQTaC5dPajquux
8mVZn7IMhe2yzeMWLavjTNTUjJwVqHJxhfCMwpJYTe+rqc8eJSREuJKdKN4W2rX8PNnz9rCLsmg8
5um/JMP+VJ/kdgqUJNMUBqF3uMkX5G9sW7ChIbUTipbs29DMXUw3hRYEx3/CBppZJ4cI94cQHp32
WP8tJFMO2JUeSpNqFVxefuFo4AzdMjOP8XVAUpcSGPXZdWhNLrfIPT1Gq0slGbfIsMohP3bvns3u
7GKVzWJc8ZB7Fj3r/RZX/8fb/ZH4e+El8D/+XJlfaZBGqLJW9QCIQfc+BwuJVkDpqbbkPU2sKyCv
1zalRk5gv4q+q9GmGQ6KaST5Aw95F1ZmXRDAZYQxgQTrIEwrE12lTRAtOarX5FxXNqPDcGwBjIfp
41C1KaWTGTgBkC794wKHEWNmGBULk8N5U3zSNlV0d7/S+gzrhKDI5RaEBOsG8jwFqguCXnu3z7Xi
cI9MsOSiSHRaWtmfh95X0DGmEeonlXNDK3a+Ey1KKipt5pd8lofEUbIkbBzwSVhnnwUJf+cAkE+2
BYDsu06EG/zFf41g3n3UknGWspRNwcLOpuibfD/E6L44L5dKMqllvUsf+RVQ6RR9uxzmRxqIIl5h
lARz40aYCjngp7JcyjVmr23hEtTOf46I8I+Dq2mXfAvbA0cZmwsNHmSHB1lgZKxyOz8rTamUksZ5
Z5CUYWYoMin1DaC3h3Mc0AovIqnF91PrTrSPETFW9Ogc0t8yefHvYpBEluc4RKDitNC5qFgJ6ACt
aLqLxORH/tWDpK5eREO2MQBqur+QQjncJBOWD4Zbp2yuXRS/x1PLDQI2cS3yKWecP2bUicM/t+ZE
bp2NHwlwjNABa7kETDRwPzhc6yIqj+auQDviz48KBC/TeljCC/m5Mdrgg8hvJHBsQBrqulpD7s5s
MpTg0Nx8fMYPNmdJCMb0np4mvhjr1gtP/SxLz5Hi2gC7i+f/HU0hgL0/Dot6mpJhe2ynjOkj50np
HiZpxEJC3WW0ujWhADmnJKimtUza4o//e65YecyTCEjmkcZIUAGCO00tSrGlnIpJyY8qcJHjXJim
oQaFNv3mCjA41qHPfySJSubilgFwbJz2Bbqcfogfug5ZvmYmOY0X8HRe7nmzShAGLraMg40IIC6d
IR1Uvh5u+gTTGYjjoDJdkiCDhcAxDLPxApCcbezksIUeG7d41wYATfObGPNjOLICwNTr/xqvunZ5
QQDZIGqxcFRZ0kjg6bFnXE0kBuwrU94TW5c3aGDPwcfVlZPrJuSszV3LiUY5z/R/pohSknt/Qwlb
mkigwZ85yja5CzXHPEit68zD2O7elA/tJXCczLf2aYv4iOTEpeiNAJryx9hlnX8nbyYO3iz0btTh
nCnCB8kqh5wwyU54U2dopNtf6omx6GH/u8AoLxVkGhzinoLSvUpiUSmhwt0AofHUDmjS/w3acfQ8
ofbuQQBFmeAr8DuNiDE/gLd1PfUFEgqVJj67/6MG604JAIxYEfBNdmspK+a3tUP72PaUNzQnRNbI
gwzoAT0p9McS965nH8U7q4GQ3+evyiPz4VblmLNBsXYobbaqUbCHOKvTf6XZZhfAq0I8ITrCqa6b
uwOHmDaoYaDgh2nxri4rcjr4k9po7ln6ddm/oga+aYSDLVCcK/ddMk/LU+6aYAAUdKs3bQF2qUaW
2EWbPw7KasWnwNnPFAA//RLdaTmHw7RxMrOE5GM5IdgU0zakKaRJsr7XnpRyAtBTmOJxxt9S1YG9
ALLhRWuPR1Fv2GyGloIaMafoPanRnrNJglhX7X0LG1fsR5/s9eKEle3j0p5H0oEmU4K23QEXajJ3
eVaql0JD3D44TqE2GJJ88p6jA+ml4w9HtXmwZsDLsQE6ZVEhR8126PG2LWhH0VsXI38PTMUbi6Oq
4wP+qg2vvWCmIEs8wSOfUCIiqFMafveK69r3v8LBxpe4hxaJKrkBLxFBsJIe200uBbD6jaPuUFlR
Z4/y2SNguhLO90LBz8M1o9GIBhcNbqi7qkU+s1r0Zo//xExI5SgdumTAT1ZJgzFu/gUc6N7x4DoE
875KmSy5ROb+KxGBacyLdbwEBBN5ITZyJECXqF65OXYxxBZ/Otb/PtwaMNVGtsqMUG0QtcGcq54b
Z4LHHN2w5LQ6PUjnAcmMRaFa73FrqfXEGyvV8o6HAvDs+IqX0hIWj9K0JXrVdYXSdkUjNJ9g1k6Q
O0/o6CdWF8NbzdwI+2XjzdzYniiEjxV6A5O7ELUDqJ9HUh/zeQGFuziC9WtN0XbQB3bYGASY8+K7
wCypdkysEm+KsofMXVMl/D7UI9DufrBfvpOQUHPbigCdLtf0KBpNec+AWNhhBs72eFBNqz5OfRyW
GcQEwPQLlxobukc6cHNw0TdkiiacK1RUwjNDzXk8B+UZlwz2iLbYkpqxm18X/EdSE6z2PuWQz3O3
LFn14LIpfen6IPvajPPvKAIp9h9w4qEeFDXovFfGBxbsfnIGwpc+urSU6a2WsYOTP57yf1+3KF5H
ekhjWRAp8PUcMpHcLIgOw2lm2Fc3dk+2jN4ocEvWLPQhWATrGmfBoWJvige3/8tDvT1Mkt1Tgw/6
c5pfekk/tjR+xhrlLZsA6H7ji1jkIzvH1uOTZQcv90JE5suSOaPfE6sfkrZ+n6YeE6mI9s4OQoMx
AtjeItPon9fmH9Gh9kJNncZA8EVedxvpcedclD2txVE8zB5tJ4GMVeaJdQIgLrDYfhBmpa3b6PLr
9DcKUgsASoZzZCiIUre/fu3iD3eTX3Ft3eajBrkHbhJiEJiFwCXL3paY/dWY0InBbI/+fcu2yPG5
N0ZICvSkiENmZ57d3hvgYaItBAYVt+8JX6yj0LJDUbdx1wsBBiRd+SaS0e3OGhr40QbnOozTpFjh
IvX2ZOC3q1mgANBQ2l8btm2gs21vfPjgZLtD+pX1U1UbeYbjIyiJwLFO8ScuhR/k2nXHC4Qifnki
GoFPTSwKZewjBpVjwR060JpZAC6zNjDBjfH80IwhJlGko/qfz0Idy2wj6rC35lF7WAK6BzMHoCau
shGuoNkQaSM1dxEIOS1OsDy6WqUbqP3xbmytRwvRKXy44eQERyasLdrf0/785S+WJdi+fx4RDHQ6
Ye+P8Y+4/X5FXNFEtbTc/vHEo2ONCod0LgCeEc6Dl+bwjqSDWm+1vtnlfz8tIMEKj+DVBwr7QMmS
1ZRYkIZUzpTcQat4j5QGbkNsXWUjZlfet/zg6J2woMn2EnyAwJkewn5VUONkng4E+MKe2Pf8yiRR
Gch/OvOtxCxxH41hstGVCe4lxGdf5zDnHXnRurFlS63Q3liVcQb8OYmo33HWkx4bJOzQfIKZNZx+
VN4bmvkEeip6sy/KGk8S74fdYePYa7l8VHIoqf7OZO5f2lYcDahdptOV4h0vJFoUQEcff1QxER39
EqUmC9lV4gZu8Hi6axqcB+wzJrcxivCTo8/bL6audSOBd7POc9Y4aU01ROaCqvJWHAE1vrrOP74E
Y+OBTicdmDh0ElhK/vu73nCCFA8jEMOLJp0wzlkLpqjh/v6/0AtE2/8E+O8Wbv9xFTurj9VYbBML
easx/d+Q13N0J8czdkKYR15hbjhhoReArWGmzahgGjCDEEwzmdiS653rRFMA+ugMTGVnTVoUAYAd
5To6s4MKK8Y8/7UACQVOgpuxMEGW3WwbVZ4H1lqT5UE1eBsFKQLSzOZ4R4jYtBrxHSq7GT0Bm+t2
jphy47Q1EELVDKFPsT4oSTy+zJvb86adRfUgyNNZqwJm7V1JgA+EgcquhVzaDudT211JrPG3S29m
glFzqkYSfDpFnORQi0GsWnC4dTOPa4eQ3vkProBDZpO6Arbr6+bC/NlzeW3saElCbtfTkFuLTrJy
W8hX9LBxD4/Wd0NN8W3d3fhT5aBhdFTHpud9LHDs8jHyW9apJxRaTm/P8vlPUfc7IkdsDa5dU73j
mJPLofmUcBHpEFdrm49j5sDiC+5c0DUlTNLbBTLyujFXGDfHaZ+kxTO5NwuNowXP6Wflc1eTNpTn
u49uvDJeM1m460d2k9CnoMyBvIuFPXevwaK1i/IJ/a7SQSj0cLZ7HMkrv0lzH0mfxaYZgXm8SHaP
lNnkScI4kHYnMGhkjuMKJmWtmh2/xph+++rfluLdPwYLRzEsrA7FxfmvMj26yvMwx3N/qhCdK/64
myvTLkl9bO4oMC8z4kwbewtgTlIS19vfnpjKDr29osZpNPjKrMY8ltgtri8M95C1BtLV6xYo3sTj
TGd6ez+9BwQMYqEcpG/cKz6u+jucM8HOmYsqptlJrTxnq8TKfJqUNCZyNe9qbYbfYv3JMKH7MqwW
3wM9xZgx+X4U0RKCli2fXsBKdnQ0eJopZl0PFSSUr9nhq5BLwHbl8xdVEm665rGfFgFsBp2Rs+Ot
gRuM4EApKfi2knt6V4dg9/AHFcxNzxJwce6xlqRuLWCgoTxdwcpPbdnlibv7J0zRrGXpFghqSOC/
nfKh+M3cyLfQytzYF6PezL0gJIptqc3zgcUVB9QzS/64JY6Itf8QHar5GmJDR9GofQ/D9f2MXhx7
lw1/r8Lx54QNT77XgfNrPpObV/CGgjEQYZW5wHQyRLQAdeWhP4n0x5Ar8hrs5srnwygOmRKeZHsV
FWfGDB0KiyqQ8cQeOwiM8cdPJYjKRBo1Dy2bFLyBa+HUcePyAkrHzp5BFjc4DZ9Y8IT8UFSi3TxO
FLRUYi1M1HgpXf4SsAgwJzwCJBxNgi6RpNvr1kZxPpAtbQE1zOyeXd9GhFeoLQluYzcZClTeJRw5
nLairjxgb5ujJIIHabpqHbWwyfLZa5g4QcCZPfziQvCvXl2x+jxvmVZ/UN+3YpDy0JjzsQPfR9FQ
D4fSpyWC2WZ9EaEqABwQ6Gh8J+E5tYr83luqXil6RMh7HY0wUfBxCvzyEpNA3pJXJ96GO/8T5bUB
XDD0d+pB7cuDr8kRdYEaOg7A2UHxYRBG0bFfvxWXT/UEdhUVLa7NSULrS3FK4TPer7TYfCEjM6oH
8OW+nCdB6KSLr0eoS7DiLSPD9kkVNU/NYy8TDJzni+y7T8V7sTQqNl9T4qQZRkOiuJGVmklG6a4X
MHMcUKFs4sVv4Kr4UcdX68ZsPlhHAzVR8d7KYIlR3cQsj4wcNwc885vQmc3xv0EowWn7wC6KgGIw
wdLt12CqwQ7R3c+nym3ghPEEawkBq4IOrLo7be5dGAO/7s3K0Mz79sMGmn5TT4H8FH3YbvzkKz7D
6Agv46SY5ggCyM4oOydcSqxQWJwXilRbu1Eu3+p5IE8Lj1QG7e8u05mEbei9lUNdA1tcUze8E7MG
yvwd7khqJNT+rlr5d7Shwm9T4D0ISy8M/PvWIDpeeW59T5EyQoxjiicklNfh3tRcDc4dV3eV2YCJ
5QVZhODzZXWvPdDxjXOGEP/Mq5wm2k4eALUzTdCy04FnaCAykoPuDzpSS+ahDlf+w73bra9Hk9da
RdlUneAbhUNC1eKx698QbZELxCVEQXkAR3wYEyCLCyK/Rt/9/YVEJwv36GKyKK/v0iDOjyQK3Z8f
8UXLyNRiaEMRwxJ4fE87kMw2oKO5kD3oOSuFXovtE6JaZn+tG5seUh+uccLjPNWk4tmIUfJbvnB4
7SjCuXSz6Gi5IY0l7KlhBhL92NVFhATQ1b2ih3pnQtyZbqm2ln8jhwc4tybhhmMJoFEzZ+VtMxX8
BoghdJvo/RR1NsMDIAjGF+MZ1m/lxtzLPdq6LIchXhyJyfKfrUDHbhjJ1PZ06w//ZQo/rTmYz5iY
kyYgQQdn9URVqq3lcT2SyecW19PrvsJ0DA/twcQXZUhA3sQA4DHD/0/iisihqmtPplIDI/36h5/d
i8Yx4naGBckmRHyBy1PhDkISOAa2BFUKyJBAGSpZs0CdcLJk7OC4gIo9nS2ejeA8+k++lv4Rj1My
FazykUDEfSSqkcsX6DQJNW5uVnyKvO0KMFPYRtOumYOuKu3abkdVC4/RHSpn+qpP7ubIbIbF5Zmi
77Jcyi9itiFWfbJlawcB0MGb8wd2XlUt3UiGrBZwyuAhFbfhMzEB/5pv2EF+VDJ1HEG11Hbw7u6l
QZv+qoJcHByUyfv2ixfuJk8E6g6O7l1QrI9Hyt/lU0qF99nXGvlKgem4Wue407itHdlc7iJNc6b8
x/HqSpdwSlknWPceKPynOYjurApSZnql9NZMa67tG5/dwWvtE9tTr9tkta8DLM4LVYs58wU4GLdA
bRAWrDY6STv6hPS/NoYPqoDcyJhQL1/cBLivUpQbuv2zzulfdK/VpdGblkaC/ZzB8HvGt+ohq63R
ZQrG/LKJruYMJzKjfnHvqXArC/DJlPQwqGE+r2sRDikYQwadfsSfKLOS2WqLnVJf7FLPll9+gT/y
UruYa51D8glsm5KNsYQ+6bz1kFiYL0ij9EsPYS9O5UlKC/XULqoioLuFtn+WrQV69A7f/58OK3Bl
l4q0yW2xLKOuAAGKLKhs53cQhNNq0jkQm2uu6J07Gxhdo+naub7yQRNfItrOCVg6DXIHXjGT0Ka5
qTRuMo/4JFbu3XVRctowxmsLPZBHdLqOubUzOL9qW1M71MeVir7ZzGvnvCvzlSruCybBd2uO571m
9XWQrIVvvEH4cf1N5LLLQGqlHyrjFs7QYt/sU/UiKyZvj6eclwK3ahs9g8baSY1R3LCzx69wxoW8
2D3rDOSPB4nIms8rs6r5zTqgYJZ4dPxd8x44zMJ5Gv/W+MdzPsrlQMHT6hiU0WdSBylUNBi7QDuM
KIHtEIPmm4LTOiyQCZccnptUYJApquNKJg+WlcdKA49pLsPSFBIq/QxtJBDPxhsSIuMq9vGsuyCi
66nqU57qgCNOOgQca0l3eGH/ugP6fMqXQ8enrq3cdqUuduEV1h/sokUODqaRqnkit6aIPL+hQI3k
M7ijYeY8AlpyM4K0hemipYtc4u3fXmdeelAvTGULkk0rmhXBrs0/eVUrJXP8Q//GVTsQ7w+ibf2l
anKwygbp0LuC9s8IurOOVvfWqFsG9FYzYBb6Wg6kfE1FdVFj5/mX5IbtPMmqOKRyf0NBKl9sxlxv
Z2qEWiDVn0RcRY+36wI9zxKEfiqVDNHs6Fsm34GJvQxlBtcBIdQ5r/pdn5AzAwNAu8WWbDX+j0vt
kE5xcsRkuMSS70OgxzGj9G8hYjQn1mwo/63/zwcMXY0cWCxvTlGZvbLfFS5BNdDkXCPR7sARXsoc
mM8jgCBk9bYkOK2yOQ4Cn4glo/x13HbpaUhub8R3vihrELkU65b9T9zUdrEQUdrPDnMwThSTYtBp
zAkEtEhGnn1P5Al1tJdQ0d3cAhIEqbqVC0HE9hy30pOErk8kiCOwnJWRkxj/KrPkAtNXn9bALvlJ
7s38T/+mVLux+aVrvRgB4j5juJ4k3DN8cfdO5P2lSah9xfM8xMkYIoo1QhQhVfQTedEFNOIiZXg6
0l+QUxSfSadXVtXlVFFO5KygI7Z/sE/lwxncvyc/qaQ0euqD/8RfkjesSgngwad8pE3ayQaxWimo
Mi6gprQXYruIWSqDSFSspmMj4KwLMUO0GQkiOP439oxhXQsup5yR2DSqf2gT0gpDUCnb0TDgNLm4
CWGQAo3q3DorFE9NAS1TmtCVQCbozKo1NbR5VCGbwfCqA7uy/nuC8N+260ojC+B6IaT8ljOaTG2D
92Oo0dW2SHUwmMY1GzisScc7nhs3lNJ1ipLNNtOFxrDjr18e37rPNkGCe0cD+uFc6B/scaQIII37
qngOY1MwnA3LLzkCtj8JyQJ7Cafpb1a9Qw6IyO5Zf8ZhdOjXz2zoeus/ZYwY09haIy4Kx5CIAjO3
pgja7NoGVSRz0gjAFnRE9RvIne8O+h5PYjD9GQ5wN7gLX9fn657u4gtARicmyz78DWmgWCkhsQQ9
NMsaoZESet6CYQvigja2oFyIfMgMEDl5sqdplP2lImCZLT9ZeNk0e+GyBKlIfd4dPZEZHCeNo4c1
NOb64+oCCd+d2gn2BBiRjdApnb/3EpQoCrwCClhV/nM/34JjlZRC1JstJjWoroRRxw04BuHNVb4u
kQ4mrdus4iRe0E2Fz5PB+cRYroqsrBz6CCV00MGvOLbx+F0DmxGZyTMr6l+7tiAKGMzpBv6MtpUs
jYKbxeuT0mxa+PFkNG40VCMWj9QDvhwfhmBIey6ZaxyVUjQkPBA13PPOypVw07iQwCAAEUEFVC3h
7JZjuxHR5lA73y5bbVcF5bb8f7Smkf931LTZS1IsAny+5ieAHLJKHJJnn4GB9IkOmaPWNrlsl9e8
NAVxNFI+VSWAsYVRNhzXri0tLi7bZgWiXJG44bplZcdd+A8goZfYbZetwqJfwgPGvwdcVXnb/Dys
1zAFqgt4GPzLF3xz2c8F+SH0sXFJ/dL2xgxjH0pnLCC7nlVKxbybx58nm3cM5UVzZi9/LuWEnsS7
R+/g0B2p3JlyLZLpi4L8Z9pcC8KN0w+K71NyOX0oiFoPbYTuezp2vh0qanY3DN7z4nFQwoEqGawi
FpXKdbGLNXcJgo11EZNrMVsu6NqzrjaFEMOvG3BMlm9i/EixJT4TCIAS1fpJpbviJ1MLxvGBpMvM
YPzNudbW7jk0IJxNM0xFpnCnv90NJoJTgHe3l93jsaSMJx5OCikS+CCmD7kNcObUKOK46beATloX
8/FkOdxn8Gv3gOz+1XedWwIEB6fv/QHIS1heojpR+A6b8n/KDOuEReKI7Qi/x+qYa9vHgBi7gcDm
nSJospGihrh0/NRf5sdoiNg/XxfDii84Zh5ZQZ7PbjtM/RoKkRa4/xgSkJcLVS8FMluSbsBMLouC
ZI7iry4U54vTkkwqfzbjTEBSJaNwCodiuWPVEymYoJ1+UROrwco84RRgwPKLj6UxrmqO/eBT9VC3
F9gfHULZXEz+3FloZNlwHq/bT42kawjcIMaEgwAdeeFMsieACpUs4wbfstKSOSjq34Kfih0xWGm7
D2yA5TUU/9YXMYZMiw7mrAVRMh3xLp7zuqIl6x0SxhpiEtB0CxFed/GvNvgjfIFsvv2TRwDYDKhR
Kxhowa7EVvxmBT6VFoIt6k16fFoXBhIie29Kjr4PoHeGkgUXhtAxpSQGloxH0tdJeLerAu8SkaNh
rg14GsXLYRNOBOx0DlNV937cIaKwIY2ZaaHS7KhNQcLYPE6l051h5w8A1XKAoKE+49JUw5335i2a
8wvgbaBMcaLbFbpB4p+WYvn7txg7eSWmIQaoIssDkoJG07FXu5z/XVM42hBXYn9auIOspz/dGTfR
Xx75SKHqDFWo7/ulPJaMz7CH9nQqqE6chUyd711CbKK8Zm0AIjPioAJ9lipYpIswLctVQmF3hyrx
14ddvanefqSISMfzz+B2gXDjEuFKlQrOhPp9Onte57GGFnSL9QWmbk/ubGyxaYA1/g/oI9zl4W7I
ZWRcsyR7E1INOAg9zyFoiorsTmThMHgbAdq8So0YfMBaKtOOkVsxttjA0uedKG2QzsVWZJCR6a2N
sV/IIA33LLmAcGmBW29N0tcIJf2puRWYK8wBaQdIiXBMX1Dqf8XBtlou+pwX3UKa6UH1e1OsE4My
kHzLYzYT1hcKfF7FVkgVsu28EOW9OgAvn2L+ilSds732GDMpn+l5C7mzNFSBNO58kmPkBTJsZjcq
o+E0ztv4zteiw5SlWsXvb2hRPvfESZPT4kNvFBxRLk21J34LB1+sqd6TjUy7HvWpusJzUmcd1dSL
LP/KB6ciJmL+XWnAWgooqQ2lLH/C0JzEavrRKBNYp+MuMjXMZwPXX1GxAdl13QM5wR6KYxchXdkk
uswVrC8DERbuJtW4u9SNFj8fOYKWAPOv+tPxDC+BUHBFZ2yqyD9/0S6+FiR/jHi8oOFEvGPj+X1G
dpALQCK/atZZkzTy5LQWBX+BWrgjOdX0VeOQN41Rq9FJIh/8v028encoCDftjTTslZQ7X2xlQN6F
CFaxzceUHuVnFohZAQYpwDusFti15CGPnBZ/rnb9JgxLWXHAO/oECSugEk2by6KZme/QO94o85/C
VsGd+F6LCFzuFFaWlkvPoKw605a3965XuyXzXvg1q32IDnhlCPDYiZBZSsM2AlcpZ3nuVx61/qq6
FjIf4msdNfn/cU2yrK4m3x6xVvLNJDp2i7Q8Prp3zmAoAQOblL6NzcB7t1Fbu8OIqWMV7FVN+foH
8OrwTKcirfm+U1amJ0jE+AH7PIP5VLVXydlt3Ppvye5sdSQ/kkJxmHS3eGHdXI0fAismRwREGIOl
Vs5yGsIoVP2yFz75EkAjIDuIBXyjOjc+qBVpPT4gfe0SOij7CW0AKb4ZviTHmyUmvBQlM0cQ7BNP
cxe9X1pw1OtKrjyQsCqU6rPN735lupCU24+O1gztOCEXU+1A3dV9TiudmWk5iRoySmY9BU5gbJZg
XMMJLnOptC2mBpfRUjC6N9WJ0gjkip8CqmfQPXuBL/7cY8M39h2H3iiH7FWXk9xwflKMtryZ0aWt
d+Ff4mKRcIHHq9/h7jymyIH4eYcvgS4jbkLR1J97M9o4HS72J7FGUg41rZw8mtdanYaJf+1qZv3J
DgJIyeY1P578SDONWuxnkOWUp9vLN7TJ8kpmjiWuw6J5RJ7kRbtuYdDWNXRA87PT9fGeYnvZDVAP
+Z1voFKcVZwchaf9sirWj8WMjsz3bTPsSad3ll567gPSFbgvrTT+H2heetmDDvUfFZFMEo8AuFIv
q7NLgsdAxZ1VAssKGU6LU6lRuygjbHMtHf1dj0Zuq8piUJR1rx2a2EMO9r6z0kECj1FY4Pwj2bXP
Kv+amvH6GE0zEXfEQk7uDm9xJoIt9jJm2TDAdwue2O9KQOlOVxSkDwoNqNHLzfnEujaHZz5XUkMR
u4LhUVY+PEUlgZ5IChJuSU1V6TC5a3l6pghDonJDCLVudx+jZIk5PxJuIpr5wTM9uuV5BBRhhG3W
8xR6BgrZRDCbScUs1WcowUpK1xjWak8nkkNNE1ihB+DnsTAUUN6m3kyop4K2RZDMRtJhqXjPDJqG
+Ud1JA4HME66ay+zy+DiDhEiuJvJ6jeJriwixDzFZo/ycUJ+rTqNJupa4WWPAyI0vtLC2aca+eHq
aJHYfZqYe9iIxZfWCn5BiuBQOeWIhmYpQYBTOT+0++ATf1zYuAZId35jwCVR8VY7sxgrNtQN5QzW
SZcRCHfgqTK4EEl1dbxn2uUROOG6pu6Bz0fQd33UfFyAeR+nn3delS4G5C4/7aa/uUe/HfSziShl
geDWpfnn0YMuAupMexpsQSN6tNfcn9XLfS1FHfo9TV0KdOAzz5fHiI3fIDjdLUzb30Hc06tQfSSG
gwiC82Mf84TaZzFgVDjjVJgFsumBfuoVcX1J6OyDLoR5nXZc9K/WQJ9tlVMoMIDLKHE7LP6Z5LQN
52YzDh7nLl1tUSTVdSDfJCRNyOwKYPjrMzrlk0LQCyyiy0f7A3zfEiz6zKb+AHSqPr82oExLDoLc
ShAkIYAvFYkZgFSTiuoCuChgS8VibmKQXjWJdCAq+7rsYrTlEXzt82Ls7o2TSTj3T02F1j23ay8/
CILR5iPWyqp99HsihkAthFXj4C359HEjMjH94UwqN0HMLSptUfioBXgW6PADHfR263kM/j/0lC9f
a9qPufzYd8DmxJY//8rUojnkQ0WHkPYMxqlkzBQOfScGWgp3PvTeH8trTTonfP7/IIgwfCf6MSTD
r5BNG/CWC5YXyxVyJQ5LXnvbNnYTsID7vshfRtPh2ifId/JqShlOY10vMttFzUVulE05/x6JtjF+
eSOoA4y0F3hwuCw1fCahwGJ1rokeWF43Sb1pHlXgUIjDKHLj9zFnMnKgzQ9FGjoyfEmMzgm7eW2F
cvPnUT2RIv1YLw4tI6D1/LUjym7JRiDG91PbA4lHoKxjdiAtfOM9BW2XOQtdFhzJTYOWFp8d0WNj
/jKvM2cg1XVg9mqCQMJMvu4M9fueKFT6k2YG/Zm0zLkEpvH0AwkOCW7K4mm0VMISMFZ2VO75nwe0
zKgITyIr590OB+hG+gKVjF/89v1egDDMdHLAtVaA+t0ao2kMCH/3JDrMTv+Hgu0FQzPtYpjUvPfG
uVSz33w1SDqcBEY4FDiMMkzV16S4XhMBiPc7eobwRBzmnomFiMlQwYun45Si2T7MrapeCxh5LnCo
jJge+wr8IHMiUNWKjBcJxFniIjqlWBUlwW3YcddF2kcrRvH9EGWn0vyS9rd0PrU4uuCyMbvBleRi
L9KFgJnFLAWVLscgrYFRUc3UuCkSKpA7InZSCQbbiqOV25LucBNVX0MqPPMRHYCRROAKzG4yujtq
oXkRiZQ8QcL/4ZqCK1sbaWVHQeBf6WDbn9awTaGugI7RgvpVXRLWVxn9G/YmA1KpBJHCqewvv4WK
pBlXOU4mtDkJ2JoeVP2mPqxX3DBza2Op2SPj6xayTuWBKZwHxb0y4mQ5Rf1bSX/UEpw9pLtMNXMw
s/yVy70xMrt/0wvm1UUWVozKmYLUBsnPMtoAZ0EljBuPwzrA4E71BpHlgWpjA749zJ0fNUYDC4u9
/W+leh98H/kM6r2G8DxHGZuVuaqEPT85tayQvMiD1nXYac7Uw1rLRA8PE9V2RYci4XKxE7HDIvem
IHlwix0QaGaws3I40NqlrWebeqJNSIyF4w9tc5lbknBWNC/QNI/RQ1Zg0ZQlgQfHgdObDi8up+JR
/0aWZmhA3StSTZjr84sLiJCIDBp+ns79VVl8WPvMdbD7RyvTOPQISo/mgCN1Sg7urVaADTa2Tv7z
UwvKtxpnCf/Wl0yrRJ6lM2r1+QBp5XLooHirVpIoz1Lt3dm8YheTjXLGmR8l6gfm2qTZfnd1TZ0z
SWrVBwgInFclD7+7R6W/TkBynu/CDZDpuK1lb6sysffusGnXwX1PkGDQZFqUxVZCKdu0RMDP+iYJ
1rEZZ87RYoM6mcylcTyb/Dx/CiZt0BesVw6ZfSft03VqeIjY3Cq80NJeTcbTgNt2wCh3r9XkOafX
9kENdzqmU2uMGQhOwxGF8MOX3SkA2YMj3xd0M4AnVIfU+t7+58OSST2zB2PkX2SVmNlb+Z+XleSC
lsgxiTjqebdZ9JSUjRkjhF9QPdNJdWsLBF8T8DZdZjIx93gJw9brJBzRyniqc5mDUYXEvc4xW2Dl
pJzhJhRSlDjPFK72mSQtQ0gENzwSh2sJljbZ1KuEg81U+xRC6yLfWOtkgRAW/4NoVKHDWjfq+SeZ
939jrCQvw8fuJDP63oRnqtvDU+v3jLubIde9h5vO6ctXQuPszeq3PoLhyaGFpPPn2fUR2seJBclG
IEPKQwtEZgb6A8q0PX0f6LP4AkmQJ05dsAXRWuij8aIZxsyuWSdjY+qesv76ESWfl+Y2y7gMw8qH
DzFixzPtuMufR9dENxOMKW7/eqrcShRSYUVlTCrtydU1EheFubTGiPLz/JBvflcv3DnhNPZAkCJA
Y/lqR/XaxsKioSsg/KGpxofD5y6rtIMATwx/52U/wFFbiKroU8kXpA/BxWcN3bzMOydab8LaGoHF
qY2YnZz/33idWJAWxkzcOpSjhKdjH9gZD9hv5ClImSQ26ELxNIS+dUQeN2zsO5IWJJCWye3OOvFe
IcT4bVpJrlk/c59Hk6Fz1+31cSondhJ0tu4Ls0TnX9+/HP5qz/+j+1Xx+n4Ilipo4EUvZbLBhzn/
WJlCPYua7Pq7a5T5+McLxtFBlHxSgSKQ3Y7YnbKXxDopCBkxA3oPeFXPZ92Z2Qjf/facl09vKKJs
YMidlyAumxXqhqgDQ70PH1GKb0J3ZVAV+j/ufzghzapafF+DRlJ85HllF5k/wq4cjF2z50cv3l4H
67hWTChbeTNm/E6iHmUWCgvmMSFB0wxRUwdTe7Inw+3opWr9PE/3D9Oiw8XqRe5bLNhsqDxzk3nC
/9GTUZX3YY5uDGAFLp7EPWrOzdvpLDKaXBCDVLIgjf1nWuw9oEOjLS01Bm4h2LOoDFR+GcEb7wPM
rW5aiecMxXlwqmTz2+5s9pYGsY/IIGV//WIhGNKRhg71tBaxElnbtj25VHv3y47/8fYj3OFloZlw
U9dbeZg1XcZYluFfCavHGE0VW3HDFN3Gh7lNnVmEAYZK0O2x7+kE48ZhYoU7Ls7wrbDoPHXnd+c2
efHr0mSCB71azcdTAdIJ4MytljWW5El0ju2BIhiaQtrwxoTVqfx5J13at5FiYsOeuTRFItBh1k1r
G03LWCtnV8N0A/JaVWq94ZYE3XlwjgOvQ//rwEEa7KHm3BdXvp0sH4RO/3ywVElrxYKoqRnF3KbW
fPpkIhAm3nSsBw+vzQ6SiqHCeVmVOSW6k1tXZQYkFXY/Kd33kHclG6Y1UJ8NcCHww6CcVB8Qt8Js
c5gMsyrbSFPAV5B2JFmPuKXgstgFFbWQXnl6BForzo5Icgavq0dkhciU9/RYWMxMoMqzcAY67JZV
f42rulQnvkze4sIAVfXOucEaHRv1YExo/XUEguMxUL+5HO/WvaqflluwVXoHJFilDKvy8kfcP1jp
I4kCNXIcWQrd8MBEe+HRMFdMMVD65SKjwnUldb/fnHJYNx8yyNSrDRjRmxfQqL4hcbIXwn+nirkQ
s1eW13r8FLPbc1bEt/8WZCDx7jJZWw9xjojp9iwEO7p4vEBQfeBHdiDvW+Pa1dJx560cy+Nf1wQA
fRClra+L5KpNW66daH9PAWWwAiENXUQ9B0/e6UJ2PKWLJywEhbi6i4llAACv4iMgi/bXuhPz38M/
kbGjBs7+cVqkiANMt2gCE0DgnLALNjseuhDy6K23JXH9HrcorWH8iNpW96l/2GgwAgTvBM2s2K8o
nrocDC6SitySpVGe/AAMZYzsSPpMJ1nW2m5mmjUsmTPOTbTILw56KI3oYtjM2GBoo3KKo+aAStAs
7EF5t0UXI0+k5Ex5lz5L0bGrultRLQNuxPMdrXSV1vEh7L8gIgSuCNiyzi4jPZeSR9XKOm/ZwX9W
CifDlvvrXDBl0nU6w0As+98x0vtllfuHCrlTGojXMb0LifHIKhAUQMaKrkG8Y5FiCaaJkuYGtrq+
k9sttszK/cgV20AgLZqRl6UpDnuUy13HDqiVS3cR90BuLUvrMy3j5HF7reCtkukIUTQvaADf36KS
1InhzRSuUCdlzqnzJoHr52eCoPt37dmrQ6ZvAhpmOAt+jAOt9Cv7A3EKGGGY7ueh2GKZE8lz5Zp5
ATEkLkAT5Vho5UM4B5ypGRYziL+e/ms8DOPigrBXDYi6ZNKMcCwq/lXEv7JFuU9NiGNu6lN+/ls7
bJ99yemNAroByfYa2KkdL7VNnj/SejJWH+70Jp8Q3cN1RlW/eLcXp4BduGjTXbAhy2RX2f56JXps
+OXxY3TiY0llBkj7xx92tgXKt5Ts9N4WIiu29T+JIQYZJVtXonbFRPJX8MlS+2cCjCokmS/cKoFy
5nmKZq+0StytqMUouvmY7mycsAQSafPLiuP98sQ+ea2Fi/PFLbF5AfU4UD/LSnQlYoQPTgV1f7f0
TB8FFVGKazV7HNWVJcNhpDhG/s279EYCbM/qyUKXpkCWF6kNnGFpzUnKwrQ2P5kCquoJSurAkyBx
5mGC5k5FYyxfUQn7eHpG7a+QZ3SsM6Fp2GzYa1PsFJ8WqjL7C8UImU4caqRGNn7Cz2f4IrACZ2c0
kQcWnENzonbVrQoVvoUHJsIXSMHYQh0FYpJDUaydwH1S1pHFE0IhzdRpWBhc8tvEvoqyO64+03aV
U6FGfTq1DDZ0M8afigu9I0m2Xoc1DOHzXtBWAabiH5Kk4uaY7aLuyP1XPRFXRKOFGZwjqEliq97m
/tMIvEnqGQbwY+GFA0+RbgGX6UL7+wi6fzdcmLdUAsyME9Tj4SU6J3/HFz5rP65ren7IF/3MvZ5f
n9DSkSzoSQ+B4WvNkyCU9IN72VygMC14tdK+nSeQ+C23AP8OCh/fmi5f8C2ggpSW53S8UWm4QhI/
FwnursjhUtEjORBr0tKpT9oxokdrp7WLSPHeKXfzhxMkWl8CHOnoKUGHuUzEXRY3XPcYNg/OaamH
GQkAVL0ejTXxlKeAU91QoPkOZsqZER4aqV7wzyHzoM+KlpkXC+olIjLU0DI3S744zQb1oPtA+DAx
45ZjlSXMxjxyftxfQF2/ThVs+9KZrzxs4iti0CTBmj3JONmgc5bZOTL6RcgoUoqJ8nxtLJtnys/j
ymMoIxV3RhA846WeJ0JpD5ULCf8+qoYCeWuq512dUofFjDzFTDPmUxHdNsElJTrJS1aHwwHFhn+f
p4yNUXHzqcMxBqpfdSR1tvPuF+KbxNnIIBKMPa1OCevrx8/3PW6mnNcbk9DKmgqFK0yBEZuJEGTA
68n20nzHXmssUjhzIqK2vRksyGMXcJFgBcjBAWqOQ3UB20R3Ok8te8XKXteNK53zjq+cBdAj/rw7
56y2KAhm5kvhBfl9VYhunB89Ibe1uiG4tN/ZFAtp3ZlejtYHAELGMkfX9mu/wbMY8XYBG3dm9R7F
krgcDXuA3ryBCcO6+b44L0jztYGwi2sqtK6vlX2fe9rEZeHcded3mXljoTDbZMG2fLiCryJweT3Y
l+nBtrANqjjvidxC1MAXGYRsGeiNfJmVvLF/5fiITXMZpKRbunWO20tpjA8z2q5vkV0H/XfZ3Qb9
05Vksg4rwbEjc16XW1duSMH2WdzxbI0YbU+n71o0xaT/ng0qvjF8w2fUxaXWXlXjw3FJAXuRurWu
GLrXO7FOP3Grg1KjQjqbOt2H1ssktY7XG6KSu6sjd85I9TVn/IqOlUwedORjsSYCj0NP5DXaW5MI
bSfIJvTHVUzXfphf67M7ZoMu2PmbEiEAIz2mXHLG7vbHBxv+CCAsM1ODlfXVZAHRVNJGTyTo1m7L
ud1vjl03mhQXaUMBVJcToYTO2MY3oywk9fnihB2AslusxvT+JjSKIlz5MFDUYxNGBHLLExCEPAot
50tMZTBB6XKQC5T4B/XfqH2dVr09Fdn4/Dm7RZnS3PUg9OqvFLbs4FBa/qFrrBF29NnQJ/NfC5TX
Y9m7NBgqsi3xK4S1wqJEFFD4NSCLSisKAfOxzKO/Hsr9ZeURLWO1Ii1tlm192hHBPF60EeizZ5+/
J/IV2d26tx70YpbLRbu6nn1LGA/4ng9mWLPFdB6nOgzpvFrFWP5agtEJ5jSswl3GkOE9J/axei/9
g9o7nfizG0Cmdi4BSMSNGYW3kE4l7aYCNLkTilAfQeIhN5BXQeikXjyKmMgXHdgKrJf3J8DQal4K
hYHgkSngi4iq63/TIZI0TIQpbvvuvhwo2XLLtZgkACwKyFEsoZzduADtvsJ/OTfqf8703Z97MZ6N
0C/qs5TM18XihG7e97/p6pXlMBNB5dSyy4VGzxh/QuFevr7uDcIiiN/vdfWD98Z8A2Yd1Fzpy4W/
UdIhwL89GXAqmZ1NtmVQh2u51/+uXUOUdy7Ge/RFhwZnDFE4enG6KV1IRPHfrkTW2mVy9TkPGr5l
C/YRiv5FX7V+BtPDeomSH/JAjgM146JyVBKUWGbbuxEoLWzrMVs9bvyV0hMQhQSc/Ctf3YFkQXpD
2oW5XT7lCEf04bne1TiULs9Vy0H2KAsPr5BpUrRjAtZNDGZd8sdMfKO/4epo5IZMN8N3qdfeYHvm
+bsSKhiGIy9cv/0sULa3VIPnX1tF2mGAOJHehl6X99/SqaUrgX/SSnT06hee/cuxQ1NaR4Vj73NT
kLgtVWRiHszXkWG/WZDCJwrgJiS2H1kKvK91LCVQNW5x5kz1GDe007gh8ee4XV9QR7cUuBxYeZLZ
Mmt+5ms5LtbCnb1EK23T9zjsoYrLCB2OQ+4ecSq4kxLLgU3etPG2zj9ls/X7k2S8Rx3sgSuYlrO7
xPuIwG4twlxZH8qzL9pBrM8uRHR8UW//PPkCrHGahTm7xI+3QW7mTS+QgyzUMxcUS24lld8GgNOD
BUrz+FwfjI3uEUNYIJvyOqtXAL2a/FIXovsWVAJULyc0CCch3HVfXZ/AuwH/PMubdO4wS1RuUCMh
MUsuKMw5SWkldYrytOeraA6G75bALFpZUXaAsIImYUagkNKBe94lPBuTek3bXA1UAjWV69ybDjDU
Ohs5u1rlt7+pUSn519G/Ynj4LL0YlWE/MFa7JZUfdjJn21aH4qHIbSqEsmRpypw4jHcjTUTETezo
njQQq/yuw6Hq0QICcQmr68ml21QiEcnucDoOblBQ3Bey76tv26BfqXPYjHvB1AHZzn91jYEXfvC9
4Jig6mOjQ3HbUTVns3gekSyWXiRKx4yh6iWNEOpNzGiYGrPZhHBHOXqywqsVcFGVTiGbKOdx0Dqt
PQ8aXqTIYirExT81W+5VuwiA+xf8CpzpUS2gdd/KaLmPEdOfkgTAXtxWlTShfKU8RpG0s/eFt9gm
+xGptQ/vojy0Cp01j3egkHN9ELAXhM8VAd1W3lK4qOJwRYG1n50oa+LAPi2uAY4FyRSOkw/cX3X0
BNx0hbhE68iYaumO8l6BHh5QpqD4gQShwn+Kn4JMW7SYQdujMp03rTmYamihuHjFBC42BABPUcKN
QJ/O7E3BrduS45pQRF1WwnMmGHEAOIr1iDaaKyzl9YzwkzKq+TQHbpZMU2xBeEYka3KbnFoA9I3i
y3twiHfFJMwTLMnSqAkV2L+Mt8XTvfZF1PlDcpYxjUTMwFFTN16od7BiiFpz7MLVGPEvjzbDG4GM
W+RrScGIobf2W9z6KSTPY57EEhRRdlqd3drLraV3IbdI9qoyzgibb/3tpNlFtZ//Bov48tL+K7AB
EbE9jCuHXU5ZIwGnFOIqTzc8RK2z0EThr7S0ShAB/N4JJ+AUFWCcxhCKgKM3RZVePMnhzX0iuCRa
wT6fLxHL1tgRayMdFgIc+FCnWbwBaYLx67WUWMWVKVnLVCzG39kYtvDyb1fP436zdvsLCoYFFoJO
4CgKWvEHwseC33R1hEnytvDupEIHeCbIRYw4telNj6iWNayASXKygG/NAV/tNO/cVxGIF6Lqy3gJ
OBO6Z3JpekFFBvXy/zuTQTYXMnXkGeVQyx9N1PdZdTHIxohh1lJTjGYv+7qIov2+uwrFnlJlAQIw
W2cO4Xsuk0qSn1vbinFUsI9nTbzz7iqPGopSu01nMTiIO+2L10J45JNsjPVvMHXK5fH6lbpDB2K/
kbQKZgxt0SY/3BG2loZxu6HD/vDV5pIAPWUGUthrMhwrtGOAfLBDGrP4nAsHAXygjHQVv6qoHoYV
Ulk+50UeEn25FjXi2DsXGknVXFp9g8c0cm1tfFT/uGDV6Lrfa30OrM97W2ZTf4QEtaQOeaCnOnuo
j1lnW2EvnUvrVXPP1/JvLbXlXbKYuZLS8MbJj34mmAbgRBfMaHwkqxdUIEmws4UCZp3KDr80qD6n
LT6Uf+ApJzbuDCG1Yj1nl3kj2BFx5d54lypl+mmPEluRthC5hCmBk+1nKuiLbZzzM7NIK7ytKp37
lmffkY0p7eOSeWQA66Tb1zD4xyl8TV4DCOTU73L5E3urSxn5QYvH0+UhjMO+4oN3DdUG4PAkCTts
EodSf3d8NX2DX4qbX6art4hNznFpfXQmY6cLEr9JloKkHj49ofILuaJoSEQXIEKWBX7SuNHc8dI3
wZyHJt90KqtCumDs8OMoo/s5YEe+FuZTI85wYv4l2AqJQUicV5nIeuo9vNqlTRcxqSR1/2mtcOLW
pHTKwSgdcBO2KMwZXUA/SMNXfzSnPrgJcIinIHM8zUW1BGTPI+R3yAjFrFOpXDDM4Oy8+MxBRyMr
1KiTN60rT0pmwmcV1yx2QLdQbTHsZkwS0m/DD9VxL5PfTWBp6SlNYVzf7hajUlr44YaJwtrhGqfA
syFFsj2hNVFwr3QxmdmTZEnuLvZpwdz4M+U/d/BpmxgRxHOkzclqYsNz/iCBUM13RMD38aePvkrO
v6TrCFWNw2euhW3A79b9nIRrjE/OWU6apI5DsF/AMN5/bMTRlXZkHgG8jS3IHhhU/F4saPvdToh3
TVc35+uAceq5xz/VOm1hYomDxeTj1V+Fzr15alNfvTi0UGIacJwpGlzvU1eGE3VLpfMHhS8WuEQS
wZrlcI/7o6gMPvcxUUvcShfxsVZO/NhLxfArNZao7pB5E6e80NR+yq4cRroGqLOWupwfEtPv1T/P
1uWu32Q06E8uUusm6Dhfn0MEyOXClIdSU7CYaXmP96IR6+Lhgr+qay1dD1FMaZxz6oisA+feNN/r
lz5xXxxuy/UXUxvHUPdW5ToII7F7nPWJf5rCQv8mHoRSd8Ku88lbNduBrsHOkGnm36TUg+i4yxiO
yLzPuYX84DbhIXs6G3VQmuSe5249Q7WrmgGA7aHeOpZw9qE3A/vAEzjz1pXhoA5kaW/h/psgraH8
kb0w4zHhY9LigmGwYarQgBTHTgHU/bxTfy6AI6akA36pIDs0GC4cLRKKVIajCE0X2ktyt2I1ntWv
wPOlGqZGAIm3r+epybqVFTHxAyKLbfaZ0o+MoiA27CBm1bQ0YWYFM58OneHav2dFFE9OkTk2BEkx
5LLF+yMRjo/huXPt27uziW4EZZJS7kRLnHUB8E4v69c/8w721oB4jnjeBngPse96B+aPmsgJNDXV
yJBxH1Knwpl+/B8fI0obhh0JNXyYZSxYcKtm5n4T0OXP2ZQfkmrK2BUCRlRmA28TvZvTInjHAyRn
75TV2MUO2QYygYTAtOSugVJmsN8pgaKKLp9yei0t+K6jA6wZLIhSbBXENAO+xpWiHh9BudZ42fVV
YiOePnR5cDgWwwtmj3nWaSl+k7erH4XbToJUQEycyFd3zb8kb2so8MvJ6ZrOv9NMsskHkmIyBH6h
t6S/F/OQ9gchQfIK2wC4Z3yFo1zl5K2bRt9ccsIt3iVMk0K/Iv0W6/sz7Oc+tuu7hQnGFxNQlsPe
lykllDfy62o/zlJXx0wX+Euj3sJeHAdihQevXsQkksfV8ZkcuYmRZY7AhuDKYOOWb8AtTV6KIdOB
cg/d3Mrpu6fDMy7qiTgAXo+rw+gfyx6fGOcejc2ovbdROJ/P2oq1gFd/fCTwI1BlqtVtZOZkNexX
KjbR3P+nT2jVcNJ2hwte6LY/lxdK//RIyG87VP8fbmX7wg4lLz+Z1zTY3THWmZmKRejKj2OJwTn5
fqTpHIb/95/X4EHZuEO8K4FyXWPdyRPN6119Mo6hgmfzh5SY0L43onWKMPX2zshopovpOCZ1ZvPE
J/HN2w5/uJFkm6BfXK7Zx6D5diHZg8IV76qyMHmQPEiM36lYeyOAvBwTV1lt91vOmJfi5cX06VVJ
Ir9nKyiOdngwhVNJeoKiYk1oBXv2i5tIks7kl6MdtyFvmhpYgIB3EFbd3fU6p+tJL/ykGfyAV5U8
4Q4HKHF/FY7bRamEIb35l+ldt2FbCRkUviaxUrrL25xrNoUEoH+Mw73GgLTqjxUVcVBipYou13SH
Cgv1i+WJWqzBayeqErNje5mb7X+xQ66iJCMkpeZsn8MtqGBXYfTGDE6antEaHR7knrOPVMEyLa+q
mKTVyO/JYRF+KuY35xM1haKQ4tCgiq0/s73RCfSPZiq7NbaWxMxfdlVQHsLzY8ASnF61ahptq6YT
wPV1QBlROcSrIkkL5LC1FrwJx74ASBnRxLCsjwTaZzVXLUOWw92UbZL5rj2Dq0xGespOHMBNTWIQ
D0lAyM35Mz/QDEAgG7/cdfllA3cGeIbpNJYK7c/+8LZjpYe1Vqt5FFpkkCAZaC5LcYTOxGFpqVPf
VsrsiXyznNtYBisadZMKDn/XtyCkLG3NlLQfGz8LGp4NFeJvXpGYaHBEWqX5W3OuQtT8+M2+1FbL
SDZ9u+IUpFD7AaKMSOPwLWZYYtHAzf0ki4TRz+mP0qVfMtkLbXI1jND5a2G9YG42e9BfXMpjL3w/
lXkizXwUCOesOdfyEOMoH+ULxB8+QPRlhOS5goRUcIpMfwK0qLYwAt9za+KMWlA15YR4/Ymc5jva
0Kq7y+D4WJLtCZBKVofxtgqDcOqGl6aadBFMMiVy+bfJ8vX9iemA5198MqMjm6JU5nXJV+uUJWO2
NFVlty84N7H3QgtjKBquDKRv5kics97RYMamL+/jKoTC3I/jnHQRBnqmZh8JvBzV7XQQbpCaywWx
yeFobE8818amaqRr0l4CPCMgOpyzWo2sOGi1lTxHdXGhVWeHmn6RY4OYgNgw8tF4YPBWfkHWNphD
9ugdEM1+anJH8IIyHrhf2J2kfGDJ0UppO7oWwTQIHvh3/WdZ+A7TiHYh4B+43ELcF6WIG8ILOb1z
JNgiuk3+jne19/RCbgCFgPCyroGM7JzgH3q3qmP6c+zPXSXtXjeyQ9FxQKVPIoSQL8RvdE86lkBC
I9LrKUPdBvzYaQywt5HaeBMu8IN4nUjBV1hLPk3MZnkqF/me+71whiwzR8Yhz5QRXhxEZ2xml/Rk
Z14byhmLvz/nlTDOf3jKUQJPIJ5B+VreERbq61HPE12EDGRgp0yIV2tUpQIVkG/lItntmexlvjrD
HXV2t8T/j+0SxKQtkIK+anFpDyKhvvHe+kyqh4+Jm4j4zZV1bacRSmGQb05J9D1GRCmRvQST0M66
th4YFRVDreOBwnnKEyLNom1El3p4F3LU5gKDjSaMDFsrqiuafv1mIbb8wBn5geeqFck+jSv04o8z
DTcsD2quv1ppu25Nx3z+qzaUOLIUXU9SE0zyiiZHF8UKvgLRmCWx0E6YKx18gZj+D+CFMzc67bhz
imFoJ/ngvW88lnjbN8NY4GBIA/K4hZEFxBsXbF4HQeiEc/y8mQMEhPH8JVKw+p2BGXlIHidabpqQ
CfQEsIYF+rHrZitp8i1IuiFk3cSWKomcLcQKlSBGbh2gPfwIe0gipJm3jk2fBkqCpB8Ig91A1D2l
0mCiRHj4VkNrYP6/EPzT6kBkkAJBeVIThPOO7AZVN3/y4Gu99l8EwCAV8i97XvLg5UFU5wRLDawl
8jiGglo/6JfAIYsylLCKTwoJ/m/CtO84DXUaeKYpJ0fJFE7t1Jh58zplaELiMeQUtMtxlC+SATTW
fhspjjJEaI9V+nm1j4wIE133IGIhlMtxbxww0wIVRHGntB4PmCoUjPx7zrSkigO0TFN1YVeuT8ye
ezyLzJXDVRH+EVDspWRgaJsqtgOcozZxISlJU5IwnuPCOkmNgWqPy+Ljv2o2GYBngXAhHPVc5zTG
0MsA/jFgeVW67nf3FDV17yQu0OgJUcK5NgKi7RVSuWi3LV16t8R7KfVIU8+p+DA3RQRf0l8BTmTe
RBl+vXP6ZW1qVlYh1EkcOR6jO2YVSNIlgRmsQkR2A3Pn0RqLjMRIg5NoegcGe/wxvm9gbK8nsojE
zHvR4OwMngiiYBxf29gGreiQd0UkrC/Wfb0omSTHdhvz7zKSSxB+iTgSapGTf4MTUWwM53Df/II/
CceV4XYIqDEG+GYLQcQ6cDoBOenSGnu4/MGigVX09Avqy1pEn3lp58ad8wuA7VE+1/SSOL1fk6eT
/EPdYvouApza2Pt4xzh8WHe6JRcAca7kj71WqEA0SDcP2cBxs/IGeEsixoB/CP4mtDGQ7HInSgmu
GnYLnDbFXoNQqG2p569mx/LzMSJqNARRTG7Wtipl2en9Pjj/3nLsA8K/lwaHA9OoVfcdknjDBXoM
scl5ucfHIwvcwIFE56jV+M5jGB46xdvbnbAlTA5I2oawmciv3i9ca5r4seVRQu7ULjAXQkLpZpVg
xqDbBqTuriCtsPIQS+6og0n5J2N9jhmyEtsMrBiIoFgmzLLlDsqUT2jT2o0ni7aqtHjIC0oo4yC1
tO8x2qs+4GWziNsCK+1N/UcJuO/Sxbk6ADf+34MI8sS3Ft4pxwo37b1pk7rpvkc2XZkf4aVH+ucr
4N1gcq4dNUydDc7K9asR/iFimnc/TJtlpjXAUXTTSDtEOU2SC4PqbahopjbokawIFVBmjscO/fCB
qDZ5R+RlaziYvU48s83pQFkKwlY7i3OLrjBnmRfz26TNvjhKNir1F3NgBKMgQO41q4MHJRSu6jRI
NfgDUShHEECtd49D+m3xxTq+v50EUUxPMUXQBuZSTJc6f3yR0OceqMA9MC63EVi/Lkz3uLi4L5s0
Y+dJJqhJKuaGveOHr2Y6yFjVDU7Bjmp7OHWiwbgCn2yO5M2RAtfpRJHASANcLgk42MpMjZdEBSFB
5KrD/bTjUieY+AIUAUYez7rrbmpQde+moDKCDJM7kD77KTCzA3dSUKJpJOG7zklSg4DlypsMwZDz
ZBJhOqcmo/Ps/w51HcvCsSw3oLGGm9BQ8u9SZUPqfVvGjgTi2I+JohR2L9aVDukkFSbnKalGyKI6
2zhqXpE4Qt42auKFcYYGeFvre5K4i+AoTabIV7G0PZDQUsXjnmWdgh1X7S79HCE2kH1FVfPfzxNP
dWsr1hLrSSApTFCkQn+RgScb05xx96y6weB1SJUPmsilRaBX6sytY4bJPcSAU6zlAcVMahNywnw1
lXLga+aujLCruyKhrSO4YPPNKo/ALUYDqLc6W06t7E+TivPiX1sNyL+zYkKs//WFapEgI1Yor+bL
ddj/uZItrbhz6ronIAVD8+2f4+AL7jvWdetwaM58W3xDjwiG6pBsSBN7rLALO7kTsxN11kPWBZpO
a6muEaHkrLfH0BOAhFBd/J10WhwU12LPcelxoAFxw4QG6yubVDqU7AxpuMFvvtqfrDNFRsrys7rr
LoK+1wI91QECph0+DcHXTmIbKCQtikFuKWHU25RayhCM0P1h0vL0MtHZmlQkSNIC7fXQsReC/4WP
sFdNrJQUMiQG40tj9yATsJGLmVrMcKvvS7y/W2yJjPTKZ/yBR+aGBI7cKA6UBXFIyLhCL34lICwy
PcWWiDsigaPYA+/D67mYs2nDom0jZrYjDooU54xluUpWOHnkrr50FacWRyzxxadOasPHtc0gSHJr
J6nXPsCnHQzbQmTQo4kypvhgPbSaPOmQgK+jhG6mx0ROLwzIsp4mJGeQ+S2/4Cmlr4i7RX+7Wb3M
JF5rZuIGXVdp3mZchAsGq1gZcwHpl/BCVfpgYP3F1NoZkCEE9N9Bwuv9iXMXxfWANh+FYeXw7EIF
owZ1szq6AH4ltIZIXpu9+uwGa/bWsJAbKKiGKcaBz2BzmJSgzLAt/j2VQjumQR9gKWomTauGnMG+
Tb/HJaNPm3fr8P77NdHtzv/YKxQDBwhKgx9yMwgJKSrdPFCAQSr2hFoDcDSUE2/zjo8P/Do7Ngmc
gY0C5oPL1DNUM+LvDIhWvDgWrO2HDYOc3ukeMWvqn1GeUAqYgrzoydcA5oVX1Oq5h2TwTN/xXGal
5naxqGl7oD4raOgAwlmqrDSfemRq2n9aNE4xe44zTrzkuW5b/JhnBiwq01/vzSjbfTbaceBtttiH
46SQ0+3RWirZucXrP3GTGZHf3GLAYu4lb1vwIwUW6I5I4fr+tPMd4JFaHj4KswZIrn3OOsN9Q/Ia
4MbAeRrzFS81KvPJPDAFLwwupzyTFaCml7vuyF/Cqpjvaz10JnMAhv+8dY901WPzBhL2m5+ZJOnA
ytbT5v7JwwOmyyxz6aweY9ggfSaREuT34XNZ1h02wUPP9WWyYlfNOxels3SeaP9xMfftvstuTwU4
3r/Bl9Bkf8yQaLYFPBv1x/yeFMoBYg6a5ZR1ViNVo5yvRz33vP1KWrSW3Xg4G5CruJMEcPsDZX5W
KWHypuMwwLDK2iTgnBaNMxGuYnjVhT/xiXjkOVo+SzzvlyE7/TlTHO5yBNThKeeeqQSnu+BSsmbn
W7fzbpBrdxv11fS1oZG+zqWmOwdDgOlY/4CsX7eKiU77bB9XzPu/ewL69f115QL6FIRlk8qU08nI
r0rtpbcIVqfEEBd5IA7uRfZ9vaZ4N75mB5ROAtKhJ4UosXIsWKzUcgClMs0AqJuoOiClhytkvqX4
jjtdbQZLfLCRFpUZ+xRDNvBC0xByvZgSQpq+Y4IS9o8r1Ll+vo9fRl618gMzcUotKAZhUikjFYN6
RPokeIcvuJVZqqOJEtrr37GIZ2ZTJky15SiHJN4beC9fAbIp7cxtCNMajB4VJAVNT1cYSj06SwKy
7SkJgGI94mXpon1YIkyuVINFJ0cqPyCsQr+o9O+UNW9eDW/FlsGOGw87PThDFDFHahhGRwFuxAXy
Vu2Qoa5cABCn42/3GP86VSXe0fUVrW7a1MOxv9Pv2WkulH8btoPulHgAk2A8nI5KW6pZ1c7WcqZN
tzdTqCBric2G21sMu2HAfWJMDw80ZpTmIrWsMy4dNp77Bco1QJRcAe6hmLIT/x2j8I+z2a5stePP
4XJkZaPOJQJlHmYt6mwzAP6zoZdKMrq3hgVQdB36iyFHUCrLH0r+RddkJo0h9iZHFrqJJmbdkmN3
R2vscro/M6jTqnZIzofR4JlmFjGXenuPIzYwQK3WZhN2Ta2Yc3eqPt+lNGhykW6TVtrTPd+t1ZVh
XPfA8gxs3sic4GTUjQHO06LZvmH9x8XH6sTw8zh8i+jnyRHi+tyB1klfl1itTu0u65aR3++C3w7F
TX37ei5KlzSmi+dEVyStfIdscE6WIkbygYiF2G759oxCLdB5Uo9jMfjXCn9PRo8HZkTxnXvvh2t3
Dfk6VoOLU/lBbHudhf2yrSKnVIoNb47kZb53abxWJy/u3qblPSRRyvTTezxC1g3plThHh7uwGutj
Nk2vv1OEKXnwdW4FVnGa3VeNKP3ABCHTqRqj68ApLruNQTw/HMdXocTkAPS9BJ/BOAER/Y1J7i9m
nLQB6M8PBzDhGN8m81t8g41FBzjrzuwAFQPic/5vGhpXEV7cVBfKmcQOowXZNS6qHmINg1HfqHkm
nMenpiLSqBQh2D7BumozeZhBEHDIVfjh5Vy4KW2op8OFy2kNGsoJWzNwcFB/4AYQvsiEL0UltCfx
RbONhFiE/531wJFX8NSIHYGJeNvtybxEbKc1DGSzMNXpUlYDoR+jXMJAHqu7cW51HufAQiRHekTI
lIZDZCLfptc2UbCsbmp5knWzVZY3mFr5ZcwJWMco2BZSHWOhsdWbSZ9NUPzhrEKiTxK/NCM2WhT+
CKPJy1N5l/14SSc6axv2c0bEdYPEors2YNzKCFfux8zxzcxBW34M65qVKqrW3c/H0y5Q9+EpU0yX
CoVaQj2xux48Z5peIIvnFpxvfQP30qdMv9fcIm0iSIn4fIjI/fmZ3tYeeMXFE6z5XAoUBuyHNosO
yyymvWASOu70ThMqCKFWfTE5qmEf2HWG0MQAS/9i82D1+A/zIEZG5Gz8fX3UPqSqlQHd6MjIuqzj
zfO2CB54RZa/vYyLxaykAIVxriXxpJxsjgV7beWfeZ4J9QdxI6R2L3oZvETmo35IC99rg4rPt+Yf
ruDAdYOij/2vNhNKeaZSeqhcoqFis+O8qQ2H7QbTEC3q4D0q3jjTNRV2RR2DaOjNd2+6jMnApMA1
QUvu7uGz5D0EXwkDrgDq43Zv0gv+W1EvjRTSbonA8sBjcc3LxjaDkNJD6TWd/G11m0s+DzU0bt0p
XdbXBVgh5RKL3GbYU7i6bSp36WFIhNEhZvEqq/iIJsEOrmjQW4q5MqEI7GgoHwq3ZN+S+DbuzmZH
ZzznKAW6EsN1ZzJpCRcT6cQr1nP4LNF6D+x1wS4NrrRX4NH/FRBthxzOGh1z0uXkc1WK4FlrYdIi
rg0wnrDucb2wjow8oO9pILO8E7uVzJK3dmyz2NLbhkoPEZR8HUdcoe0n+YDyl8cMOCdK73bhK2DP
OyYqYhXprd6boqK3RlqqFq1QkUT/qkuy/40msdp4GgH1rSvObC9QqFRMnjc/HEUBbnsg6/ZoiWHl
hbRM61hLI/mQRp1G5JnnTN82GNMUJwPfcQ6M+tmgU4AOpNRMemheS66mdL8FgjGxJyCHCIfWqZfL
R3FmD7TTTefriyIxueDa6OUlamm3skrHjsuPYxSnocYxiQs+yx27d3wyZOUkze0GId9N++cLu2iE
7PrKNYpYDHCfiFbiL1qQFdgmstXrlgB3lfbv4xxNk2U8oBCvQ0q03CifT7ngmXkEvq9gaiXNWPZB
MfUCBD6orkl9VDTIepIxSw06idu24kNn+ooN/zmg6U0xm6co3Y521NbUoTIMjE7oZHVX4hkXobg9
4af6DlqgrIccXQ9uYQyDhaMz+fbHSuJ+97f9+RH5R48UFfBcuG7EwUQMxuq7Ty00Ecuv/xgx4rMe
JhyGIw3xRM/naHx9ryI7EuHEeN0iAtc4Q/hKtK2nGa+KgRhAEKThy33QMGNPnHaJ0xmx6eYe4elZ
pOMo/jLERsmF6wnofKLIsX7eV9a3oFtaM4qPnU9vFKJOWTGTXbTITeJmXsY3FpdfGnEug6amtr6k
6snXtq5YvXj4yn7hFsQOj1hlHo2yLaEwZlsCgIjcZ+7i2zZeAJeUCXe1AS/J49cXOlyWwQGJgeO4
w1G6a2uqcqhwfHWyqGicfi6lOhh3ZQcSqZSO/01GgQfQ52oDthsgpI5awQe8YVhBJ3k+SxrvSMyK
5iCq6VofPWaZ3enIaMcDV99MKSSw5J21aXu+/gyTxGyaCI3uNmvj7NiftfRIBro4G80Lwasct4FB
sQBxfrdlYqSH4vxpjUgxjQOw5TbH2FX/OCNwgvkR7HBbCiKMtjnKlmnlvEhclYvVqDx3ceHNNKsu
dJY24mdPnawOXGrHwKTWUrofEXaDYaklw+EtPJZdf6uip+EkJUYR8qjciUBvJ4q41oyc5l66L2jS
DBSvaAQhClH3SZ1VLEfkDibiUhmdZ3QBK/ycoyJtrjLLycvHXjjwxkfYFdckKCGBcaF7DqNvSQdF
hG9R4cXx+El7tqBK2gyWhGMA7t0mqUgZj1rXgNJHHxhzN8z1LzQ1g66pQmaTvRFeB+FpZ1rPd3Wg
o3/tTYsjBMYKxomi8TMObtubkNPJiWr8Oj1PZVhk/vbOsTmTV0dljewgDIWzr1IJXqtxmB3W6Zkb
ZDBMI/z0P3fy9degkir4WWjsSY4fPL4SUqvxzueqcTuHNUWiPUJ/PtluZPcf7xp3v7S8X/M/G4Tc
hNI3ObYumZtRBm69xMSmNahruuN2Dsbz7vGFjZCTYB6vi2pcwWzVbHJdYQCWogkebxKbuP3dIbPg
MnrvyIWTr40WHd7ZwGsNfADsv4AUkpVPCVAYAu+Sqmw35G1s5QYKfQ9rTJWwmLLHXV3Bxf2xgd2/
k3wksSZVoUSf3UW7J3n/iu+PbFunigQxl2S+OD2SDM5bHCPmiAcKmnjMaLOpKYN530glzkS9DBFJ
cNFt2wAksZ+d+fnO8LSnnnWgSBDgyv8FWsyAFx/04/PXjGo1OscDnK09Zp3b08nN0Xqz/9C7tyb0
Oc60fLkXelQOOQS0llEyVREtZPn78afcqYhXfOUNBmCjEEc3tFwB/NX2vNys46216j+da2yM/W8Z
OyiFwSexhcVHnLm6yTDqMIlP8ekrL7fi/yQWGKxdDSRBi4dfI/5+DgJV3XtJkVXu2VbHlFQpfm+l
eTVUGeQNG/qJE1pf58VNZ3E77CVApfCK/9GsKltMTboAug5HQ9QNZDjucXkUbs+MQLyJpaLY8Waf
5qtIjwmMHCRz/6zD52tgmMtSIk+rRlgJqWKGEe5gOIY7Yq6ht66Dfw0UrGbNMOvMCk2GDd5K3ZLo
Yx992DgIi7mr3LkbSRLskEoYJMqVeVgOzRxgbdz8ihNOWQk1yi5faG/FUNaB1Qn9iUGjswYUVe+R
0bDlOJBN8uXLHQZSmRBhXZ7vQAykEzOqvTzBKYC3dFCkh0Se2aOtZaaP1c+jOhgd1ib6kHj7vkZN
aMoDzF5sROc1+K8ICOjr3K4jhWRXkO4MLq7oH5YO/GNl1hs1cHEr4YDTsG03YFUA2cZRWixIXdwO
NdfO6218d5jw/YY4P+PxiPgN/Z9sDljBPa3VhSfFR/nZ+UM7gtwvZYzyCIJfib54raC1mBjOawaS
mTZS2i+DJGBD6Cf88mNtiNPwDEjs5ka+FkgqMLArH+1rSLxLhKGnSSY640YDoc67MsCxOTn3vBl1
KUY7p4Bbgta3lZJZE+sOGf/Y5gatE2ikBe4SSIo7iRsk1DW+JiGjN/6dVXCuoD24cCpN9uU6TasW
Qwo7+DXTwicedXQZF1mraHh1pa5ZlhkthP5DHWX46gSlvVIJO/HKevnU8a6VBnkO6lvCG5WJhUyH
oN9TfA9T/4ih/1BhWBqy9SZ4YCZ8NvpmRjc7eOvPvtJO3l3BBjpE3K1B2RYo4SMRxoCl9wHG2hGj
ZJraei8RFcRUSHRkf0oJak7Ow0PSD5q6sfiJDiApsaFrGaJebX18jEi7qUfoIrSSWiArQVhjXgCy
zX+Zg8bi/GuxTlvk4StKQ6QSV+dxQsYq3GgXgpcKMv5lAD4jdNBAh6hCyZryWu0WdqaojS8UQjMT
ghOZNihLF6ytfWhSMZelqBKhPeBKWtMo+smkdQLURr6ruMa/FsI3mqu0ak7x7GJS+8fiZ6SsZGDZ
5P9W/mjcmCbQv2indKo0UR+08t7pvLEYEuBQyFiIpxOENEmAEvRe9ygnSLC/VMoGbXa3aa+vR7N4
94WSWbNnYKJr0IsM/izrLDlk8Hmd71Oj7mhRKc6KAwVuRgwSQtQ3T+hJurWEZAqdhSQz0NZt0xCe
/Hpp08stsdK5XKKZ4nfwf7wtksx0Zi+thjKJmiTkZZ+KR3PTNr70mh5wXLSTXnLg7eARNzrOlRZ/
ONFZWHDWGfcG2jVFSyDtk+i5FfnbseCH3h3m3SHrtWeKGpNqvL2OaPPhoHnT8L0nFF1FcB55R9/V
LGYG9/RiEKCpA5kmE/VRabD1RgoeZ0iOFZKKXyM4linjpJl2/ZCQVIYEAk8f51eRqHm6/tEekWOG
OymP6fKSDhkmJYPOlOg22fUKKA4qh+tl2SxfmbiYfhMG2B8xfhGw8Wx27rPOMin/gISG/9TgPKSB
udVRut6tEcsle/qhOx55gt0DEpR1l6YNzCjLquI3w4RUTbRMMuyTShHNnmRjf8OFI/OKrY6qF4HV
bGTa6CdgSOwNQSewJ6OJlVUu6/BqQOzsW/liyDterplS4iPckdpQ8pQOOYIjFusIHXeX3SaWnYLM
7F5NkAdBdlUL2cVU1fRLhhCrlBpdnWYFbLIVwgd/zdSxktuuAVpdscJmlcNkgdvDVbwspWpgobx6
3hkj3uTl905wKkJ2FG0HWI1QLTIl9WWuq8MdzrbSzocDie9/jiEGoH31vheZyxPtK5THb/QYFjSa
N5orBqqAfdA4JiFFoewg49LVF5mpADPVDoLLXdjrjs0nIf91cvCAMVXQv68KWJwqaFWt/+sDVTsH
1+Dj0Y5G+fGjb4VWWiCl7TX7iEfByyKRx+0xc+xPDIqPLHlld9mCw5cPP56d9btBd3hOmCcNKHyP
UzXYKReHAYfmewlRaiKxHoAYPrPJdfPISol8OueQAOyJLIZVo6jtifBw+bC+As1bX5VJ7pthOTvz
7W65uslOStz3RvCN1yYungWujd7HVkolQ9A6UoT1+1JqW/YlF3/elaxWL0Hd7tzEe+YIDj8CEnBQ
M9Hjr7IVx6cBc6cB2q1EbFWeUeiFenr4026Y55pnHj1sAgS43tygw8v2ryD6+//Owygqq8nYFsiM
FgXwzt9m67frDJak/TNWCWTjVHy0zQie6ND5s3PHtFHwTLwXJPq2ZsAW3VOOPOATqBzWEN5EXmF1
dUyZjEnqMTT+lqyJaq6lb2fGkyI8q/qIBA5gXMN1AY1VqGfPITNg09UaxBXJ6q62YMOFHCPzceWE
SyumvPhEdRbEPIBO10cm25lenLtHIm0uh3bdqgpqQOavgeSsu/UNj4ciUIk4Jtu7jcYC0lM8xq3m
xC0gQ4z+AIjSAdh+Rirre4XCJhVfW7zzteOg7LeSJlEIIanMDPRLkUHhzE5i8rtRHr1xnJLSotTE
1wWWZGeBmF6tyGTmsHK5QdDTy5bvo7z5SlBbQliRn2kXBg+B9xUkO3l5hTqnpNQ5utei+CzqCmFu
tT6HI/QnJEVPbeXqUaqtUuMky5HBkvXICz9f/2aMbpaBeZiUAU81vsFPTXqEjVetGSLN3W0q/tdO
5wPMh78g4+om0+lkoGwuDYs7UX+gzb/Z2JJJ+33XCebAu/31lkaiQLGeLcsmG0Mqz6ABdWSTITLr
WhChhHzn8XJqlXHhcxLz2OvrMSGdKNlGO+Gik/4P5fiDKfWro4AJ6Kukbym7tGDwa4SAZBqCSBxK
ttqQaUif8xPmXFGTMyx1QXnbQKeaxxpE546ASBqJpYUK0daivisa2VoPG9rMJ+wrMh4FUxJzU+ho
9xJOQ1wrvuMSoBKtvHtGjBCLkcgL9lEIVT5Uk0YlFLojsnHQh8o1LilTww2XpH5id9RwQez3usUb
hP//NuTdtQFqZydjDibzqTcHzAsnwBF2kL70FvnZHEtovknt92+TiuS15HBQjH0vGuDXUn4aTaUH
ND3pSxSCFEDFfUbIUz7ErhMO3ZpC87E0lQ9tUtDytDORsTbhIyqaQZ282AXcJkvweaLSAciIZqWB
phOdRlfSE56nAkT9tsbH413lOTi37z04R+atPeH3W565nE7hnUNTWwyxW58GOvbxwC3sr/vIuYJi
U970lgerMzcu/kUq4Z38sVG0TVtUvRUL3ABHcQp8avvXF+Lq0PaAXF0XGON/aPfpAEPgOd+a6wvq
7+X32pOPHVGrWgFQ1r13sBj7VbV3XClq1viMC8zbOLGkoWQXoaEUtRtC5eDp8mgrKV5WweYMbC4q
Z02hhDbEMlN37d1DU5mlMTi0OxTdj72vS6TnNRwb8ZI/Ak3TUYRLgyHEcEwP+G94vlzHcsouZmHx
oN9Lybmm4y6nDraP3gXHCXk+bRj7gQV3f8C67VUfspLd7J/eBKUXJHbgwpIk6DXMqNmd1+PxHX6n
zXRaVU9Q5Hk9c6nIgiK7n0XYjFrIAchLZKNVbaERo0/MGtkwMYPcMI3jJVjgnMrmw8eGbIbfPI5K
t5BmFDZxXBwRg6OAWY6KuKzA5C6+Wqe1/SEV3CZNIppbuZQFmzzNQcE3XeA1i4uFwVGVP3Uy8aaH
GSGSk2mXHG3LOGoNK5pNYP4kLvRj0FDuZSVcrn+5NGjdm/IvcskiUPZyUBWxeenYMZWK1znbn6pU
OSiQlZE/oNi2nxvxi9X3PmEji7vMrg6Jg+7awPocR2BBrloRWDCH4OMdW7YIH6C9v1rCiCyKp4h9
kcp8ryHl1wGiK06xT+3IijcLhmZsgPYwLEGtnkGh3FWGgIWUhofFu2JAjNTGFm7/H2iLP7mZj928
kx6ZH/fRrH4YvDeQvoaLEq+89UH/WdhxGWIDBXAJcwLcxc3+YDU+/MZjEWuapB8pfqzwxTKuY8RA
58RtDzM56Hg08/e5D13sCoLPDOzZXGFgGPgLIpYZa1J/Nq2yrvexszeqBXGOfEgIvnhBVtuoJWYs
BsEpHD/bO0AAof7hytM1kXLFLkBicYJa2/BU3QVAlLaLgAfo5yYDwyCwsp9JeAXIHfeHYKT+fxHd
4QNoTmAZNXRqt7rNgSr0hAkxdLC7yBzu+z+SeFz0miU8p/9WM8+42ODqQsK+vXdLwEIeZST/859K
qZxvFaV+ZpeXjP9g0K/kdIt6itveJCycNcuN8Snk/UylrqNyAZIqYEPLAPNU9ssvRKb+HsUBOJnf
e7e5TYZGQh3vjft757G43YnPKb1Yh46rU9/CZ4PJKHeWR/pjvzYDNn9580ce+tS8w+Us2/wAFYUI
ex6dNFOFfGbTqxhYFAP0RRxh4l3000Rd0t56Oo2SAK40Be0/iBmY+xR2O5sfUd35WDj/TEu7f3Kc
crJLHSfm2k4+U0zvVQvq1yCdiv4Npk93TIiDhbjzWXTXaoNkA3xh82ZhT+r8MzS5mSWFequVqA7F
eNIExi1z0QM8cCAgpWRF3hVu6qptzLSHjvMzEF/G+h003kq2/k+ZcjyrOQ8551C71LZ4UfsAgYVN
3o+ton+3NQDACobb/xa+dkGHRjrnJByi5JB99zjXovJrN6B7DXWNlNCG8Mfk+wUcK8lqabScDk69
3Nu+pQo/vePtfkK3nu/HyumKLKfA2miTba5G5xzYPY765xFB5sQxlfssmh/EDgG/oXEzeAQ581OI
/5pRmga2xK0D4iA0UufQyKuElnvBGZsRJp6h7QbwQxsIPXvD6Dy1JE4Vilrt7g1D+FVMGROUJVZn
/ug93ZITJaJNO3u6QJ1E4hWUl/jKHaKgpXm4dPXwNuU8z5K9XObKNRRM57mi6fFXaFF/Assp0z7f
aze0svJyyY59iICX7T5Z6Ka2A5TMd+cYx0wMTuc2OMVZyXPDm1OMGlg496kZ8LbSajaclc+1jNrB
CLRv7c+Sf40xVemsVuZe4Xuk9tTgxXpGFK7Sx2k2TGOzIXc7VDpoqO6PK0WCScfc1TMa6dS54SgY
vaE0NRjAbCJmNRrXBXb1+hx0PuyKpakKRnTVzHQXteooPQ1nl9qyoutbyiNSpI67w61l8ljXfxDv
9sFuK0mVs/sJmqgqWSrYz5w+VUavrcQWv53r7ysE5T9tnzHP/Tzk4c0QVXyrOacwSaq8zPgdUP5i
QeeePgrroVdaKG5NwyTjQCh0XIKCCak6kQMfX5I9hKo6CkoCWIQxRYIhftHmrgK2zJR/7l3a/fOA
H9qEZAklrKFfehOpq+D12Hvu5Ik9h1jeJbAwEe+sHVR95oVJZ8gziAeJ7/ejYS7mAP8KJ7ZFdRHG
RfykLKCr9blm+ufUsvubB5hhvmovSK45mrvxEWIcl1/X+TmrZ+Mq5l3wRHtpXTZ8eLkRcLxKiz2i
DmHPWNm5Y6o8uZBjbEANxk90c/SASYev3fDNsatIWQTin0OdhwEgYPOtqYOEs9ou+JnZ5GzaXV44
wUqXpit44CKHUtL5Zy0Z5MbpSXIf6/3ieC3X9WreNESKOWygYamvX5o6S4m9P4p+eSnoxeFhaALn
DN4DxqLipMj4sZOO4IYCWSgeoDqfU+0F2cUH91vgOINMGfCad7peiLebdBDvS0GA4fwsUYK8LzIZ
mMZhMCRMj4AMW+ybabuR20klQYqwUOpw9reOpbFOsKYZyHSPv14hxCOi4OykPeoYBnCZaDVDC0zo
7Ylx5BnrM0Fk42vXAvWRhO3BVthhTsJ9d1kKGsqiurfzDJAtoQrt7XHIkbj+63A+o/F2aBWJxMmj
8tzvfQtf97IV28jiCt3NgSEqudqI076grApNqwPI0nQ+ciRV7AX4UCDdvZFlNTE7KtW5/tXnGXzi
LF3HT2/f5BM4EawsAvIzMaSAcLfPRpbHmBIYiVJpj/KbKxtUqQ4mfEBPdvregHvNP1F/nwMo1h5u
dOlDUxLdtCgUTq6wGd8yUNJUtCx08SoGsBcTfhsXQ0RDWE2jt3yO/27/jSvgAYtQKSS8R+BtEp22
UmfrBaWXlNrVVJv6RSZ6QIiiYQxWC8iIARTAoazZyf8syatzRZEXla9XYgqYMX9FmqILAkklHT+r
ZFjxxcImlijMm9f4FhuYLxem/pBEonurOtp+iXFkNNWCtwD4vlg2gV/dfard/iw6GkSQWbsJXK1A
7fXfN6aFFdX6/NGFQ78KUdYz3/kmCzowPm53tmT1okcXBrJz+TL5rkS/OTUWGC7LS5ZUIT3nh3zE
WWUgTb5qub+COKVt2CtxZzqZ7sT0yXTGPD3nGMFPlczuXzTPjkhPEusxm2IydYcUP25VZfsuF5TE
HKQConbn/qS7I1onrBrD5ZKMQztB1kLbNG3OkHEDkrX8HKEuqcH31f/TeOM37dLlgU+t/X/LxWFT
KHzPwTCdNABOWdTZD3Eo+MGvNZU23F91GAaFyJTICFVWDR8TFhcWNzyYEuisrsLY1N0FWdTxow3T
aF/zyR4P3vXps5Y0qUwTfuHvypzXYddmixh5HUumMSXWFuHkKHi4bBcQj7xpoxYsPlK3kjMEDfPP
6AsMtSbrZ6zBdpnvvNGgbNe5Y/erWoZXdm+8oIY1FglgtGAzvTDIXeJAyFH30LbPC48106qXBHWB
SXPZtgEIw5SedzFxViy+Nu8sgMc6tOAMxinJCHWbZW+l6JM51QxRUbWdaKDr/23ritMoQo91nEHF
LeuQo/XXdiOKs9HtxTKQD9SPbkzF78h913Yo8KTglksb83FGBjFBs/PePeEvw+jKv48uYEBpGLWP
uQJvzQd7bPx/mAacVBN0gZH7nh7st5yMU+hKH+qil5MkNIfYCrxsjDTu5MUPOmlHalexPHU/UHVI
9YJE6PiVxX5WtCPkPU9AUcxiRE/QRr8nmH317xWvzKfFQmUBk0MQmGthHEHGM2zC6zu74Z5zQLaM
an+8ra+aeVdHdZyDssaSUY4k3608O+LC93Xhm1ZKdmFhqjGMQQIDW5V1ocmHMIP5uZQPBnOY4kaV
2DeBHizcku+ajQ4kFlHluuOn45aF9k4TmEFcJKLNmtTpA7xrx6ToV+Zz/15cLu8euhLDqrfz5mNn
w/VUjhbPJMY+Nw/5FfKMhZ0LR/uhEtuqGOMSY3lLpcpc22mWsCNeiszjH4+Wn8AOlB8qyQ3OKvUX
9435fqkTSRKR9hsPplY66mfF/FTYtRhuY0Nlk3Vh++lxrFoDpGky78o9mmvN8OIFVbkZlt9Ittie
3/igLTHFfKMx32lnofVgpNU7/H+jgqvSDohQgP0a6aV/vpt3pMxfnKQDakN90CMK014keC+VS+xd
cS1WU4dlwSIoJUSg8q2gb3R3JQ8Fb/aomd1VRKJBDKaLrWKff31v0S2ye9waE4qjj+ueO145P3y3
JlezjsGNENzePJ4L6LHNEfJu1hclcpZ8aX3d2ielnxxRVYjy3EbRuyLhMglH4VNexvk5Fbwlnf0b
+ETiGaMX7+Z0yl9R3MT8NM04UokD56gnPFrSKPWJb4/9Sj6NdHAO+GXyoZCkH69dpSqg0dZeu2x9
wktGLr3SHm1Na05EqSB8S4ZUD5a76d3Yx2AsfWvldLpP/3DdtXm2TUqlBIvJ/dTFhRxp6ewS4Ipz
mm5R6coCwxGrt/KgSG3iV+pl3PwHWjz0KowEgezIdBNwYXkX4564qEsafrgDJcM7lx3Vmg8dLXVd
AEc8OoeB1Qd4/jxjCDHGJZvy4GRkYS7Pto99QUeE3n9gnN6U4VpQ4cz2xkQJXsutFvwYOaiTOvm2
wIKpmyOVHOPznVWBYyQs3KUtAetpX9q6/pDICDpCESay6teSKseJuQPyUoLhstkkm5we2nVFJ5et
V+sk+p7kvFrHWF/h69zdKpTzk2eGoKleP/HSQi51JSNJ+/7TzIh893HfV/3rUMPgknZeMCnEpOuz
EZ1JUeYwx7Kr2gpciMkeIy6/76igJP428y5HepE8l1h8gq4p5ZOS48EtM+rdqZa0YA27lBkvKnoj
BVtXg3+hqFcQCLpp4e+xJ8Z82vxcGzSBNTJixjCz+HE+xxG2qQgyUxjduwFujqio+ap0fSNoTJ+O
7E5sv6FKmHdOGKENt9JVsk2fRDd4lhTVSU5PD+LVgE7X5SlIX62XgtRunjl4twvE0pMgz+0UFT7X
q2Xd7qa3QKSH1wBC3IVKW+sy+OyDTW9HJKENmNGi1PYg37cwdio4FSYf62Ofa3bJ4/3M4dAcP8pY
hszTBDvhBIKJ7rGfqzS71BIEvNnCd//zs2w2gYj5h/4hwtJKFZpWoEnthkF4gZO6gYaqS0xhVjOV
PH7DLQ0VJuuI7eyxzhhZ8rMhGErr640cYZSoXyqzIOCDyQC0svz2by7EvNJh9P6b4Zfw9Z7qix0V
DiINrj+ZecMafTDAhm8LPZquzdLF/iEY7t8MkQP69Ud2uk+MASNo2IlHM3jK19Kbn6Scfy6Eku1N
bO7BZcxh1xE0VGpQ9no9tl9OF/wX6sK5r+0/p9bYmXnpexA1Jd5q9AYqiSB3Uc8roZdOVMo1++Kr
3KmZ3nwrI7OnSyWK4fhdnw9b7HC7Qexpv4AdhUhb0aRo+pfNA5gToNc97+YmCrKpIg68wO2w/0sr
dXqv/nypj4tEnnYCRBy9AEn6e2t5mUQpldudaiDYyZms83Ileq5DLsBBoV8rCi0N0RNL+JP3jmfi
ESOjOhJTTgsu1maEvppKmxwOQ7AdFp8UqLpnw/smgqVvpc81W2MBSgtDFBgMpm6w2Lsnz/VzZRyP
OGT2WjVZCOSJ7GKWZIYvZmrwi7ywx6PUJkvgjlmohp5ydQju0EMaEfQ4o3hm1jky3u+sqWHWCKGn
5agopSsTT9O1mNUpTPVSdicyejsbCjdAMkoNWtuuA7Oy1eftydO8oZSdcZbo+XpHG46OXJPIe05c
9xzYzwLoMDvCUIlY/dqlKXYNTDF+wHx5PT3LEIDP/gmbzd5ojYmMdmD/WAJLIDebtfswfLNWMP7R
8GVP5WpxYdMyLzippNgoe/ET78vHZz22YRjRtsorLNttoYhV81QfNvAAsGieTwc8tYHwtcOXK1af
aW21MV9IPQPcGvG9RxiMDuO3cP2ns/HVcJ6Pnb1BpnIZrbHhmNDsP2Y89vIOmR2Ou8VPmqeIOQZ7
KN9mC4ATmhjL4gysIgTQYEVgaZXtd2jzn3woT3KfdptK4fr0DM4rFPKUrHo1cfba0KAIFX0ImUdN
Ls3AHEbcGfgiE7PswsPjiyieehfWdMPQavQPlG+kcCtvU+3CrZw1XxDtw95tUrWpzOQFUEOyM4le
3W3WqvpbW8YKsFuyyaGZ8ldhDb+xFkQrqF65rvh9oWiJOX9AI+Vk3zs3xOokhE/OsDOKDKDEZcKU
hACMN/jrjpi9tH1cc/RVJigawFJ0FBWfRAxbcGep6J+KPDgGk9w2GcVd8Z31b/iTkYYWm0yS7DTc
GFEwX1GoScJVo1Gl56/9PLGLqFmE0X1QIwmC0+RCBivLIMNdAge7s5/nFTFKI2wEXNmWv7Qtr4qH
aF1isk0+m7n2dog9/NoJE11DZ8g8P7jfFSCFnjRHatR7Jh7moGpGXrTP+M0x/zbrlbotRYJkr1H+
KepOSVROG2Skzt69FcWnNiBmlVdP6ljKpzrlzmjWEKS0q4P4bk8TE+3358qXPFJL9A14O0EFQOgD
4VgiyuUZjlqxZnAO1Pe1VWJaSfIHHIjpTWZR9r1kFO++ug7siUTu6zqiah1oPYp6Ujzw6VdjZeRW
XTzdj74NLT1HDgJpKMWVItbM4W4H0A//9n2jA1cj7GraQg4dYE5BDYhIRN1uabUPfysytiZBnedB
wDhVGTQK2dvwooCKMaQ8GbF6VZZNm5uBcQua55mVuFELNsbJZJqz3NYe08z91XMEgyZ5LTniHTSG
I1mXtEFWJRylolW7jFVcotL1GImkjxX+ADEv0sMkIVfHMlqsU8nMwh97TXb+6Z8F4UWSjyNinGKm
6CGslp03QgxL6WatW0N4Dkb3iZsBh68qqKqvH5gP86h8dyyX6Q5XD9mASDGjfSN7hiTYUM4A6y4i
hpHZUrerY6gFPrZ/61/9165cXQOgSpL41h6rtXDkIfK19le5MM6etPri15TuwmkiOl7iUb0Mu77o
z1Ehaupqg64uERF25oycIkuTbQN5X8WGjSd1DDzseNq4TzD5DJRhJOjRACD4gvsGIDFkPSSpK0p8
fSeuN94DbDzc9vBzWkSTadXHzNbRG/Z7Qy+tB+UiEOl78pE/IRx+y9oCOABKKzNSx4Kl3s3qky+R
zt+KB1SJwlJ+mGfVRKsY3tjYBNGX7N5KfV7sc2u2DHR23OGTJaF4BicJJrbFbIUqSQdh2VKtkLN+
AQiNziYCjQ8X5YbgvqFVG1jhy008atczrPCOzlnBneAu7aVQzvMtXCqIVZOfn/GqpFlu3F1yKL6H
U6Okr6k5oU8sfele5IHyU2JoxYF+l+YU+kn2TcMPe3xIoosJpdnz7Mr1h1cK+z3L6lbQqxetZnBn
LYNW1pPsrTZIJyLVuxDCeP58uU9KqKnsQf3bka2lb2/s0Z9Woinx8ILP6fnL5Yz1YWNchSKkyP+f
0h2jBMyuqCYtSWcs9rPtVCErgQ1zLGDX1U9zAM+CeIjIw587qJrUT0jzJk8TmD4Lv8TtgaeNCZP5
PksrEVkYKjz0MRl8Npa8pAkGp2/cVp/xCinF2s0H8hCIr06mNqBoWbsplQG2spuPnHlXY9a6FbX+
jCZIsFRsYu3jFgZcaonEa7RDVZqibL54Rtku7bCLDt+N+0Tsmhe377PNiMsQoKoAFqREFSt/Lzid
olQG3NK9naOsvl55jMdXO5/bpxRyTr4kw12c3icQxZcrog5jbZ2Fiuvw6G/ARDYnTJFnkYGmRbCQ
V7flonGfa6kDRsrDWQkSiMoAO/YQUE/Z8R8ylg+LKX94VfHNqPdrJwd8n4n1TKPeftJ2jJWvztyr
IpE2munSH2weqLWDhmRGMVFkSEemsxDwLtU2DS0hu2txTR8XlokHEmuYslXRKMyCEeK8XwxiRaJu
oVnCUEOqJdT+rSSWDkW0D0tKTyyW3+qlNSW0rAuP32B7XS1rHGdqUdMCLAYElLqMpbuFbtetmHg7
AeJZG+Mp7vFOhGQLDnqkL2XJfqb/Ei9/YzVY/DDdO/ToUwu2ANclA1R38rDw3T7X6qvZZNMYIsTy
o7kG54Rr+G6P/IT202BjYwqx23G89tNIk8oxl8ZxwcWb26lKIASvlse5vXJSprnKlrKCs7JGzBuZ
jxhoW4R6YLU7JL6sAwgXWkXt8OP/iHzIrIV/gn8HrjxJHDdgrcpjE4p/J8B2eFFM357dLfAWHFKz
eanLDVXEIA0U1TubtA2JZgmCVAOiCee2ynl8HwuwMf8wWBe8uzJpAUhGedXFYhbXV+Z9uSLWqsMT
aa4zeD9CBg4rlLAgEhQRRJtso66pOEFw/72vliwTwVATMJ6hFb9uvRO3Cr60we+jizVjH6gEHrsJ
CbHHHim23Y5pSZcEoO4Kqeii3TXMc6J/kv87soP/Ogtv/XVmXbsLwsKC8EcRGECtOPnRdfuygZBP
1W4fsj1Q9CgPRaN364gd/hC2xPBl4h0fO4Oucesf6YddVsdaOo4E1qpUZTDlooo5NPMKpxk1WpTt
gzcafdNGqAB5HiJpQf+QzYRdTF6DhxYj0PvTBUAupz1srYM7gS8PutJvU7tGCDLwFYfNN/7cIYro
evrAXpkPnP5HKROwAK7Y5dsr+pfoSnZs52vhgPYYRHsX/l/U7N840s5E3yc1vOhVdKLcrwqXi2tA
AZrnGqCrQQmwjYuA38Cnf8NyVuuIRxIGpKiFvRzabwjNQB9yraq+EZFleC1oQNU71VKfEcHn7Hun
ie+os72txeWpFOegz+LHayfbqBQkPOudx2D1uNtyjFhKbj9fZEvhckrg48r9gnNugZtbe2cXdUrn
WRFMyAgm/OMPTNfi2y8oESEi6qdRPdwX6Xu21Sw9CV30KvDIkCbSz96ZDTzFAHDrdP/9nxFu0ojo
m0QMKjLo36L6n4HZbxmeiZeIqThbpc5OUjtbj+pJCiyYP8rXzKhMP2QSFPPSuaU2OK5pHgBxalmi
2hQu1EowgWdW3bIlZJtwTCi5fvDi0FJNJfM+uveX8wfL9KtpkR09hxg3yKGTucoOheEuZ+i3DvMs
3tDMOw3aBkWBSgAFFVc6fhpGSBTq49pocGj2wY8+8vx+Q9hrZo+vJGo+oRoEJXhBdC1wT5spV8rz
m3B0CKif+xHFrcJaZimdY7lCugZaWC0HK8CI/kPAUHUiaiCx8F86UnhbbWYmGOUcMucDwemwBBVi
KF7S7srAbSq4a8zvxG6yrPGhYeIzxfxLiP2krZtSnuJsaeTHwt1xxDSvrYVHLIPEAewne8RwkhNV
WFVVxMzsbHacGJX0TMTOTrzeVfxUG7qQIp9cl8afgH7mVB0kmNgzXc0YcyF8LqABtXKM1JHaZCN4
hkPKFfTn3lpP8dIoDTiXASceKtN9WCIwRpLY0r6s5jGETKS2Kgt30cB1azIePh4hCtLzo9TGUYrh
wK3ApMm3/vpW0joy+oY0OC3OJDVKR0XE0emRbdA9O4czcAPVvG7KdWoiS9ZDr38iUc8gMyvuJvFe
3TSlSw9XiAfyqRBaRpKLv0YSlCn7+LXJKxKZHSUjMHV7w8+ldeuknytAtJVNB7acfvB7b83sD3VO
IlUvJZGizoTo2GCH5OuHI4ApLiGpYcDluE2yE2qtVyq6GiDWuUO04qH3PP2zpYt+HutgUl3zh1S+
eZhVLGzg6umJ+R2oNwWw/gvvVdc7Zediafov4vzmuIRIK34CsY0vf3NhejtHsyD/d4DoUyqQXqO+
uJZJ2YDph9FeeHk8uaxNBGND1H67hpzdhuQAqK1idWqDpbP7EJmX/WLRpPidIOYdRPWWRotcCp1A
RMiFzA35JDfM9B1XqC/y2ZcD8OYr+oOzmta5pM9f9nC7xfxvUq+q1RiT609d/qpAkayJU80SuXmq
Et6h6fPfKdjsdYFuVsHiE9iii6HmAF/hiaBoRWdcvINyQWG0/bGF/G2LjfnPvx/oCTPXJA9U1rEk
Xk5AOx3WJyIO8K9bsIMEUQmarYTvUd71Kyt9tWRgjwRmFdmUjdHqtJXbrD+GwiUxI2+qVMYSm0ZJ
Z6qukYhnNul6a1oytMAWu1NlVAgLCOg55vS9eHzbtG7M1sDJCjKh9wqiPOCSsuSwFRuB6bO2YrFB
Armn/Nwhq6NkoT061bDqgIZJYk5+3wVCV1RHhJ6ruv/oluF7Y7h7YJgBmIF9T/fn38WqzEin/c7W
Ey2P8NT3aIHJJ2N6VGNzZgjyn+5FAJjsHlEPiL8wwTaxEipqjt9woM6utTH7sgtC1AvOGyrKExRi
i+Zq67T6lps7wplhQshxd+C8RT83lvTm0Ag8QN96ND/BUgxPLN8hM7ewx2oB39KCtOzSNr99aj2C
pVWPRlz3utCukoStq0z6kRO0BuupT1nJkWFpqO/YdH9Cjfs2VoaJ5sDSndxq20GjA1HW+lp/+Uri
Zh94WzsqpvJ5AagIfFnvyK86R0mUAWKBOeuZxNV0Rs2/Jd80NYKxLOdu6Ic2eLsIJyRa4jWgl+B4
b1bx+oGgapaVxCl/dBOqdayQypMnqf1o6AwNmSAkgQXrDzmMzoyL+Ncvm2pBOLto79JLbUm5/vjT
wybwV64UozFYF7zbuoHVik66X6YfCxgbKFTazTLEVGqTvp6YeC7IMT3T+6nSW2C4X9/V7FQCXdqP
F/IbShYwTZotEaq9r8eNjaklcALHDz/NKQcjXaCvSF63MmrWum5MYt/nCD1t9B08X02U6kUdyfU2
m2yHSeati7rJvkEE0JSCc7MuBvYb+GP4/8qk1YGmpN7Q8Ep5BjfDqBPB9tFBhKWYIppCuBYxJS46
RXnVCh4CIxOU/wQdWnLJBpzONGsmml2tCa8vDMexqyZC3b7RWofIiW9M2vSgzTXFClAEHYVmoJub
LX8AT5KPMO77ThlQmap7ayfhLykNW3HOLOkMSfx1gc0S2gxWEM0Cp/HrCAFxwkfINNMuHWTNxMFL
1hhy2TWZEQFdIsLkMRL9QdsZ5psVC1S7Ske6XtsH8Vle4jjh4ohaObXHsa6f4eGQqusZUeXdxPZZ
bb2YQLxMmYnlKN2RYKBs8qg1Z4eI69AGs4ZMPzoQ9ST2QnH+9xgov8vsE94RzwUw36v8Qia+Ska2
LeyqN4wqWxPLFwHGYoP8t8eTeirfEHAcBMUmcO+jeAIrYWfCgKuyXXfg5s51WpkR8eWVS4bDuX/w
lwlv/oGblG8ynVKUZpPUcLyWWXt7CnJH0zySCvcXFesu2aexMTt4JAkBBfjXqAvKqsyXOrZkmXKP
GfUU4P0UFnK5GKF8jB+mAec9Pd1l7Z2TuyuJoC9nCGrNT+WfTlEs6LmTn5AfYW6efPZPFGzX+kCp
UHwMkk9lrDLqJIKoLR8Du3tQKRnL8lKSQfz0KJTWW4OgxdbX3sncsg25KEM3UFUPoP2BnMsfuSuy
YhzVZtrE6A++n5L49URksajUdUwkqm7Y4uwICZqkPFt8jOHYb/hW/YFPhNSq3G82+JAWPFi1cv6O
qBJhzJJV81dZerQtRzpYA1YGJz3L66rUNm9ukOY4WzjG0EP0HyhZcxlHQNsrFH1nncgNFg+xtye4
edW2Pzo/yVk+AuXjiokVb2kqAMmeaQdXBlj8vAOr4P00LCK/gqpuo5xzLUDE8MQrq26yiMkF5VA+
5q9dTihVAy4IrCiNxmuoXWUwqjxKl8RDchryhrk9YNSQywEAEaq5gVIegJOWV4XRLlmANmp1q5o+
u+2donJn2FY5yNrFwmWl5pWY+lMMEFyCPHsN/OZe5Af03wesLVkNKy5acaBq9n3e4bivoPXHrhw+
fDPZHifNsF5GpoIA7EnomIs9f7So0MepBF5Ilfcko5J8WjyxaArqY2dTDooZxmr5KvH3iyE0/PVH
0B2WF2z05SjJtUVTG2YVLjOc6TWsE6ZUnbBcqxqoOWqIzGXrb9Hq69yAsWuv+ue/OouKkAwnQeRK
gJixCGXOvmKM2R6OoXpECgI86stS6iX//XySnyQMiG7i8+9mUfRqyXro5thErMVMXQrO4STz4Ali
gRX2XQVW87UN7VKEyd0gKPib1kSDnUr2UHlNL8tiMvzlfh6ZStRpjMafvyqzW1YH1VOmg3Aknqr/
CHSoQtL/xa7xY5bvNIATbsadJIcvbCbSfzrUJdbrHLnp6L0QJLKQqu/YfTxe/gMvjAlQahQu06vG
VJrFUcjDm9ikUUIuj/ErcujaIaYCMicaRowNz7AiOZeRf6y9t9ZKUJAfwA7lanO48pPXJi6ddDuq
ueKZGih23uwz/2iciiudIgV9/YKZAk194CPSdzZjSEDPcH8Kp7C8GcwLlmtsxN0fcUf13/izphiM
ucZwC8UdP62YSU02zYyHKSKXADkFnrAtqCkVK6fR2fQdXPeMcliNhnea2fkHritMf7gCAaKHW9TV
Ep/9hGRk2iRz/PLUKTzygZ9RUnxf2C+z5FG05NYno7VFVOXV2V6JM7opTiHkNkvBw5CINCnHncDw
X/zKqjvHVyr038rfWjIpjx1Aytg+vQXMjRjbUCwDnmYoSbSa0GxqoX15lI/cZh3WbwYEOyCJdCax
i1zH01W9mxEFHGN2hS5No12SdA4LPlw2kwPRIyR3b7EQQUg4+XasomNwcSvivmjYxQFGq6CE0zn0
QPS8kgM/vW1WIGI1GnoZbY5kq7i30b2C2jdqqYbzH7D4MlGmDebHsbKb96OjxJHFxGOI/HiBbXKr
wbrm1NKVbDQ0//wlRw+SDHwWRYRXPRAJYzKw1L9nXwGGpHoClFJ8dBWyjYxy6ITP8poNkHc6/dtw
1cgHrPWNN9NDbzfWjING+PaCxOAjK0rYMg28j3Q4GIWVDJuEfhxm2OIbxkokZlujcTLa8nHXQrzL
BUP+va3XHLXLRzIA0xmI+0SHhjLcpg6VRvL9ugMZGIztAKk2vt32Xm1FuFrVy6TOPWPfvTTexEgu
+ThvVyz/30FkHeoFZp0bc/DoCWEnCoeOlN/O3hdywhpVXI36vkEt7U2bWcVWcGvdKIoVqfFf7tMY
TYIctCus8uOeAbQOO1lgsc4H8RnayAi7l8iLpP4IfbbV+uyb2WZneiiGHr/ACfRh9Zch/ndtGjgK
YzTzYLKi4QtgGY1c3FfRBKvwAr23KcHD0ws1IC3NDcRIe9M4xzWhz1/CLxfBhc3pu9Kes5KH0Abv
2SpHrtlJh1zJv4vQaH2hy6wXv2Kl5+XfJngopd1ZpKC3zZJqMZwCFuAJv5FU49T/LALOXASWshI9
Wbb3agKSSO2YmHEBVR1uK8BFrJqzwpzfzeh0q+wW7wy5plh7iU1H0DwFlH+ee76vM0BnOKxkM0KG
LEGXRM+syq6SsjpBQDQRl6GQL5CK8jqc7pE0hSU/YgT21219atPyVbOYP1EMHwVPEJQDg57OFToB
qQKz65oKvanjPrCXX/LejM69+LSrhzY4hfLhvB/vfFfw2RpwS+SYfFH0pA/zHa0J4xx3JzTgwq1t
/XMqX3sAAj8Sgq+mGnYJVf8bJh/5AIrW0KNaKft72ts5FH2N1jh/aiqiyZVJWQ95n1NfnoDamnld
yn5EzjbBV225vmBVcyFujKe3lv8KPO7DNpoNnIUjnQIo4CuxoJ1KkZVxAFH8qFO5IxdhUH3rx1wn
EJiYdEzlwxQTwPdyaWFfBp758PII//soCOKdlBMmFOgF230hfgMtaPlUwaOZBh6RrWYn6IbrX0js
XOI52/yzojJlOvqz5FGSWGxuaJ+nWaI1FAuRwAom8531MoTvezNvq3YUMb0Xq7byjskyuYJX5+WF
ZILE7DEocUIyThBtqUS55bb0rJ6Q977kbtTtUfr1jPYJ5lbk+Eyx/GjeEetitsXYQuXcBYHMbiAK
cn+dsK0xKGeUfrx0PKoMm6aPgsSSKckJ6l2CdyTuNCB6qy8m2jpiDoxDU3YvqWb2We8SUd7WDiZb
1cb8T+iZ8quVmSjKR9dn5AX8rRZ/SiPx+qD6UXoEndhkY1YMpjWwuLl1F9gEZht6u5CjpuJz9pvG
G19nzJr8tsRMjdZMm+Uaa3PEAzCsZp2NBRUotpcGip9WVuSThTkqmBUDmf7hMex45CGhmlIAMEWo
hmtCQ1SlgjRufaPcWVrGxDQ8SqFi6zt1l/1yTIp7XG4WWPrlmOOW+bVB+uQlyvmRd8fUeuD6b8ne
kYaIex/d2No4RfZ1BN9GGoSQQNLiABSWVEOCJ1TH1mEZ6rBLaZbF0SrlxvjoA9/3mqmEN2pnyDRS
7SKeBDI1Z0WrYWBcKgmA/0ysRawqksDJz3ChQTVoRHOk3g059gAxUA0TVLsLdnyMynhEJNsPcpAq
rbMaQ0aY0JW1uPfgpig+LbAV3qPvOhxqg/AFMAtie84ZTdsaooi3W8IV2pb2+2lKIjy7OvFYzwEJ
3bpppCfQJMT0JR4wFO2/knslhPWDflHHqe7G3fEUTDjwR+FkcABB3AJ2Q3p0N6sKIIdTt4+5jyI2
rDbDmKwSLaOq+P9kESXYs5Nww6FP75871eHqN0Sq6QiikN4dX/O5JDtwFZ7W9REkC9RqZ5Aq0Vgp
TsC2CE3SKvSjnQ13qyxHDEG1tNquL0iQgpZaid9Po447X143RNUKw/mC9OlUvc2ut4Eze4hIMwz7
SIZ1m8w2QykvkgJRlibuUcHmN85iv1N/xaWUqUNRTjMweCn7mRLMSJSbI9oztFhyY/A5f2KDagME
f2FWJ6kykdpS4qeuG7Z1uoZLHLK1etnNStkZoUbtamO54oNigU6jHSKBnv+Uk8OPrU6eOoEvyNw2
QtbdHAmpXQYAGcRmYJCnET2/xS2Sxq0Krhv9mnWXgRZ3WFtaeZMDCnwum473EaBf2X9aSJqGeM9n
29aVs63KJS6JqJzeXVueLPMcAHWeRcF7+t8C/EJpQ0E8K22e9TU0Wh5Zvzk1FWd3hfQxnNfAR9vV
COM9s+UOymVVLknC0g+Va0dsZ4l9k6gH90r5m6jFcv5eWYVlORozpfCzp86S8gqOR7s3STlehx2p
73bai3T456ZHbUpaRwcArTun04rRCiU+RQYLQp7lvdTZAqWA/KaX4mXpU8dVJQTAXLiY+h7uX1bc
8hwWez3SwqB06/gO/gEDIqfSAT3xTmYIDMPOLK5fj9LiBazTxCvVDtr7rhD38kY9/0TFNcchoneB
mGST+GZIjYzuRAUJD1ObNP7fdyMsDYnbvz1FGhcs06TxkccLygi0VVWqR/380zlaIFztpQmCu3k6
OeBmzubY8wSazXGaw2RPtujxHNDhgBRBo9l3wr9beq4fvJMh5eeOeKwBIAruPgLtdxKOoeCz4iqI
ZgdfKmc6iLVgziwe9kaUIxO0NINwQSXzg1XBbEG8BgWru7GSsWLHtyB7MzO4TbXMde4GJGvGV7FC
YfdWg0j1ALSNphzZqirfgBEFjOHJYONI3K1khqM2+TQPORw7IbRhwsVHPLNA1YMfxKhEsT9YgxZ3
1y5U8cK9diPNaaC+gCvvGMj8PZDLSJrQB3sKkeMmjPTRB1wYWJNwhMNZhRECjkS/ckDCkNQmtG/q
1jLOGl9X+QTRBmwDN/CBtHi77gWsmzxrdH7vNxmpJeoh/DJGxWUAa/oGMCFPJhkfeMul/ItIH99E
UElrcwEAKxr6/8fuFZ2bpCwYuB8akNDtZcVh0c9aal1d46xggRHR11FOCqIOKFcihBqK4TPCCgtk
JNxa4e86VZT0+WmHKplEBj4zFQOZYc6J39tQkSB+JgrVt9pt4xYhJ4xvc8sFko2UPWEQe5AJ2kO4
5GmRv8ixmStG/xA6R1sOEe0X4rZ6t98FZ8JmQqUnRm2prBfrmBN0OuObh+g0909Spmjo/8BaFN+V
l8qR3Z17UK35k2st2G8p0DHyPza/adaPmfJqfnpYkK3UtyoELW/NgilRc7OReT5ikf1PKUiCXi+w
mNMpDcMU0+PjEe3xh6QySHmZCZZklA+zXOcqa851JIhOWF68hGFZGDF0qE6jdHv2E6NxwA1DN0/S
fpAfiOnOf8kWhQnCp/29AUDnlod4FDZNReYQ3fcOfYJqVTVV26Rea9N4I+DVhFVYImLc1jeKacs7
Ey7Vyjdj3g4NlzeM6DRULOpzPGs/nGTQ/CDzCqnGPo655j6z9GcGHEv5uwxPOTeiwOEEdyMsCDzm
upNDKqPz/RKg+u2nIrOKN/rqhZ+V75hTAEtVyOxZhaIkTz2GkeZUOm98XOzOfOvhiedG5JDffT6n
QB2d7mmuGhWFy4p+7WyqJQRSHwK06UPA4aGG1hn5Jua2pIpu9TqmFGe4Rof5qq2jb0yzVihN3RxP
w0A9X430QH/nugA2yDtYkqzLh97Y/zDVIqLfUsQYXT8Zs4Vmbp0zuK8YsLIugjj74r/47uXYbPDb
s2iAnipqi6OYzMffcb1gaQBa1AUhbX6FjmI08rXXLTmjLl7A4D9HkUZKXv+mAKTuJWLuIXXD1i7U
8FCzOzlXm7jaaNfO5ugTIskutEC4uyjZmgpmFbGwVbTQj7Jgkm2b2c4g5YSzkHYh6zRcttrzf8ID
68UcRY4McWeJ/onkje5BySA8EOAmNqkv0xhjF5GG0XGY0oJTjYAa4ufsD3rOUoMytAJ0PHFtcDUw
d8ilg6JN5iSSN6ERm29fATPd4mCFjWAmA+K2chlmW85LRaHwJUyQ/m6Ah+YxI51whpXxM4YUVtia
J6UI5dtHdMDzZbt+8geVZ4VCKRWTUhsB4C/5O9s1IwJCgxzvkE5pfzDfPSe8Eo1Vo3dHLqNN/fKc
6PPc/CDYJUOElpPNMW+y1Pygv9u+aC9IhJZuYhN/rduaOPnce2MipWW8mtTQq2rLrRaVG5ikc5kM
yFTWM6JdsydS9uy7u9TFT2T9nBKzo/GaGMY/J4scAprXipxIVL+6l5kxDPMslktRJqFZ9h6BdXrQ
J4cAHuuLUGwNfQ+RmPzLtYGS3BXQiONeWop7IyHQfJ0dskcwIVJQr/zXP3+kirrVxUeaYMoY6p/w
bFE6JuBmfjW0Y7qDSQ52w/OPP+Hc8jTjNF/CmAlSW1Er11jkG9KSs1hbBv1jwY3xp0xIWwcefOto
SSszUR7zQaFpgS+W3OwXmtZUPz+7tn5/EDKYLsyYgqcDkb0EG1jBonwywpgXinIZL6dZZj9g5spt
mMAsSrctgfJ5Vb9nz3sdYRlE4OVQVOUdGe52k2/9w/XGcs156hraTGjZ5x693xelc35lqMX8ayFi
NAIoZ6lJXl2fwkOhgIi4b0yOYeZFDCsqVZGfiUmqH4BBTmylzDnSzizZGWKTPgEcOROpgbLgKHY4
gkpT08mWXfHCBS5PNQ642TOXzexFmNfqzahENrO44ldrkGnfGRCdl5IK1wpWX8BASKEahMLNr87Z
QYKsG+dOLkStxJN6Zw0CrO8pTsz1WL1jEUmf1/QFcusYGurqJpX2/VaMYrnpNUpSBj4eTuoRPZnh
cBFuJZVaexkdFSmlDxn10Nx/X3jO8UXcFXwejz3eEXzGicm8YeNg1OvEcJCYSI6zZlEYf2Cup7lK
u4Nn/ehYJXo/7/oubUfikLklV2kLSKPdD6Nl55GNbjqWrBS21x1MwNi/hWQe6x2V+8YyW98TQkH7
dEc/4WChnu10ZWmCsXDp+NfJ3yU6/vm0uw6qhrQUGAjHsYRugRQTxj/tEr/eJB5GX+TyvGo5yf6Y
HSTsYUNdDsw1yB5FMI18pJ8CKjIF09iPF9iAGxzo05gfH67yAe6wFgVMAH8fQqevIsmIrtYjbwN+
gM4SNz718YQVXllxe/Wv/I/IAA2rYHbUkfWAnTAuhQN7tEG7v+cbO/BD7X3X3DSpftqn1Le8DNY2
fKBFY8KXEz3v+GkcQnQDTZh5pEgZX673OIemut5hCwXFupGbB/wR2eXMuKoa6Ovcgmzd0MF8m/FC
KZnXHJBT8vwebeL+Zew60gJZpEyH67/L7DPp6dcjFuePf4+8S0n8yZThWNHBpd4KCrGCdE+B3dc0
IKc1n+DzHG3gwAVerLI1yvaG+KkNU/G6CqpNpvjX5pvCi8ahqhgXdemCPCr2WN9ZvPnr5PLMZnbD
dOgmmAsrsDlCqIQi5w2eS3G70cGzcR7GFnjpR9fGdLunsSHCJ9jFliGzDBS8bjJIm9+4imyyPXo7
VUsLJQhEG88VhUO9vFoRRHsqyQL4quv4p7enXhbdWVvDV6P8B0KiPhX5Wm4rTUr6XyczN9fDGu3I
Z/SXPbVHlGCn0Y0as4xei5lFeNEEeeMo888LuQEBzuShW5hek9WDGkQR3i/khHtkI1fweMcoJO9V
6lK30W3C/8OPMxU5z1umyMx+CcwJL9A6AnM9MxV2cQ3xl85ZiOdFsuS/MZvZk5C9K4CbDF17BTVq
SC2bMKNJcIy0Cgluj/lC1KwvAU8RmAk2DRlcr+PpGuN4E/E3cCsXwuEkBs53EJ6lRVrabwwtabk9
tL4hjgN0bzfo7pMaqvTbe24d6rJMeQtHDfwTYFDqu6n2AMUxuGgB1a86UL8P684Lh8CiObOhoZth
6XIAYXJwyBwWD30nr3ik47WSORBl69KHZvCg+foK+eiNXLLfccXCXQnZ+8PS3zIWtNYPh83IUz96
wfoCK3f3wU0GHFkKg3+R4XssulrEo51vxxmKwMIdMf//bu+PNVVdkGFj9pE1BKfRB0pkj2m0nBjB
FfbIceqnWDssvCVAPjolxW2GbdlEJBf7E2gkOWlx+qVcmeNhLL4Y40h0+FR46USCWjyrcnXYxoqs
T1vrdfZDsC8qavuk99oEzLrS1tv73XLq67prRZSWw72KouNa+FIyxLLMrmPPrGuWKDAHIL2DAAXs
7j6GMQDmwlcc3ysB4oIskFilkqeOTF2qHKWLCHcAgmPN0xoDhXcovvzlmO0Nuadl6HJxE+fTXwPA
gABd7LMuKNIJL2mfb80ZscOkGBtp4+hWU79ZdZZSoU3NP3NS8vQngZTNXfBr+MQwYtRrMGdUuJc7
YvUhFvsObtIbilw4viqcHrmclvL0MjnbS/w4CA4cbXCdR18NOg9Ven136+0Nfdxx49Kvn6yfHGpN
icgfHfCGGvJvIasWtBac+V/KH4XA2coZJupJ4AbQnHx7AFY+tIuoY8qsz4xGwJFFzxIc4ZsoVIlr
ICD43FmB5s10v47HsQaU4msAxy/9VHDR207DzCl4LaHBU4flVvWG4cC5IIC1YVR6x0Dwhsdmx+07
N/lyHnTl+SerrP/yWseK2w9OPn+NaPw10zoWrYyVZyS/bkCdj/2O9ptGUf3nxEQE+mFTXnb0Mzdz
t6UD8Mb6raPm3w5JrPNaGx1XyIBTru6hJD6LY7lBwI5tNI4YeGuNVI7NHwi2WoQ7Q1Rx2+H/B7HV
vuCcZh5Yj01s/dDfeP/vLpflViLlXRu8CrAH2+bctP53IZ+aFqUL4NqozRusHHz230S9J8daY9iO
eeYKoU+H5z8aW4Ypj85xkYE23X3RJQ5XwmZKK8BhkYz3DZt+GnS2EAcEL3UTt6RzXFtoHvi2tKWr
iQoQ9F2BIfK0ScWJIEfEIlQQNMcyotg2VPv+FnyoE46KvXOQtT6NSuODnPPcpRYJ4jjDBX0FVvZ3
UAhM4FS6W0Gk+VRnX6C27k0pnRH9Cn0AqY0rlnafayKcoB5PaKMudP+F3THeOoUcnKT7BZgXXmrG
J4XLYfSGKoPS4XMQDkm9TJWRWS0zDx1IE3bckW1visrPm4mgB6wDlBSUREBnh0xVp9W7xwSoGwsj
SScl+giT/s8mxKhIBynItXmIo4Als11C4EUKRHmnvDSzEATcwNtyBPqeeLLlC8yXtIbMmMbMs6Kj
dEp/wUG3Fiy2lePOg47upY50+Nxk6+N73HR8BDD69Kbu3EOUGVjdy8MVsABIHjj/GApbmFuZddOR
NleSDguHfSZa7CDjAH1HPBOaq1yi5yl3wdfr/Tt1/fBFRESX6xGU622Cyc0z7gsXFodLwPXBjHDE
CIHMxgGBNr49S2E32d8F6QdhYoBDy/7hIL4HhcHAxS3N3psdP9ldi3ZnvzRhO45bdKbiYzXubzV2
bvag1uBRZL7/Q6iguw40qYTQDh4E0xC5YhJwQWvEEVMXOH4tAqQgctEyAl9adft4lwRg7jlpfg+S
fsgv8kP8H50jtOKJa2o0TAyhOEgQejJITZfS5e4feaJAPbRraaDi3teXfoOBoAhGpBXFEEmM94dy
NvY7erFIhWYWo6QXIk00PEtU97x6yJ+tDX6jaLnh5A+q/hRMZ16U9gATY92rP35UxgssS84g3Obc
geuAY9AFFgEczmjvHrK7YCgiJL9cvWAYVctc9fa7la+J8o2cJXT8ehqtH+avqIX1tNWlhwQxM1mK
Olyx6ZlItu7hOtN1ASQQivYqfn/wbOpxuPwBPtJn7TpDlA9wx6AHma2D0c2YSwWnjnapqWA7xP6k
S30yVu3vANmfXNMZbW54mosoaq5wqqutbYRdipE6GpX7lcpvV6He6nk8RhFU4pLM737XddJhI6Al
WY7nbZPSlSV1FIAr2m008KhNxflL1w1nLZQ4Hk/pxYSI1QEoj2H15osqbVxPOtCq/khgWugxq8KI
7ogyAuV3ZmhFzChyQ07fRUR3cIJE6hKFRu0OPs2tB5hqNJyq69dh39icF6tXiYP4BYoPG1UvwGUN
M7KzNcKEVaZ0SKBYEiDkg7xC4/ajXDDnl0kD9yae5j3U37OCRTSVafw8P45JFnM4s5S50Ar4gBjP
jpRtD5fxf7G6KwKofP9SQzhS2fdcMMET1otpRagex8HOxsg/oUFgSEyMg9c3K7v/MhlMdH7sdriu
SEGu79ucWnuneeGCVM7slpzBk5Lt80+zIzzr5whUbjLNpihtP7HnCtkKSWk0lHDfuGpROGdU1UEF
8g6JnV2MQAtmhvvvzjj6WzsPOWv1us3focXMr1fiSlPBKfRyTofzbGFSGvg2Ssbuh027POgz0s7f
R1foT89tx2Unz7iJhZ4Jh75L+l4ersYuZKCLThBqF7vro6O0UlvcLrN/HLvrwAgwxmq7GWj3f8l0
v6A+Wy6LEbZpSUyTEB0u6Kvmugrztqnq5gtMlGy+n92pt2gXFWK2K3lT1fHpUnEVJvstcd3wEw3h
NKizzmbQcSizmTGjMySSrcTd3t3my57H6udn1ZtZfadP38Rb0nOl9sPJIQcqT4DNm2Mh3XA+ul12
r0EyYSMaqJBnkFXWTRVYvJifavpj89B+Uh1jExAHNK7kH1cNLEGI8YSSncJ1pf8I67PvsmeEtRQ6
IkYpX/5ljDwUS9sd7V594rN8BI1wKyJNycUw/aq78NVitZle/V94fB/7Eq1M0fQ2Ry6KanE9PAew
noOikkDfhi/Hr1Yz8u9FuAQcyp9CqEMvwVZide2h9RRlQqKFUBW4MnEUWlq4T3rkFoAGLTwIZAkk
UGuYbaNH2CTKqNENkgBCG0Jsc9G/hD05VW/bZ6LyJu2wiBjyNg9Oimd+W/O931gYyVxIdNivG3WB
jqHTqa5CV+Qeob94XbPgNVzb/xhy86bwJ639irPnE7kANpdu8qQ2NclyWzg7JioLChMkxgSnTglU
7aY+8ugi68OZgglbYvMJjPYFtR+XUVft1uei95EJZ47TgxaAhVHbN1E+wspHlr6vCFuejRPbKQhj
eNPPCJHDLVOucRNYLt58XxMsXSR+npqeBGhGP9Ckgk8D9HwneKuScyRl3ALAxEhWo5nFatx/geub
IXNLbTN9XhWDxoLb4kUXvCHqlwbAiBNC4xD9/VsuxK81E3Pgsd+aS4S6ePZpTJM05lrCg3ghgG9U
ovVdR2LaqSG4HBR+yWDwQiS6Znjv5tF+UeUbq52vXknT/V62rs4ejtuIn6pgDGopACRxQvvSeo6v
nBFL6LfoA6MkLSBi2dbngjWixu1qv7owPNleme3NnR8QpGE6IuLvAsgBqmQrL4HR+vk4xb5tGPvO
lMKVOhvR8zMzuTPjrT5cCQ4c7kUig7f7ST+IBR3YkPYcJh4pzri7HtOAqGHyEHRzFF0sUx6mdxn3
GDcGua74yY4djmF+Y+rwG9oXGAQ1cWPzNBk1OfJsa9urH91Rc0k6DKO4uj7DMySO2GkILEm3bOPp
Yy6c1C1HvmOv3iNXQjxlXRIxAwDIslhVfhjwvy5C88/uhvljqbp9quxahpJDphHff/zaf/6keeGu
8whAe0FMasciKs6yLYfccWo4CUJRYRdEm82QBSPWmnPjdFk3W72AL3Wm8qnP8kpIZKvA3AQFIFq+
kn9WO7ZaVCAoCbYqQZCXeRNjTM/0fCnE55RfJwP0TbRtTryScba4tN/ehIpf8AYaeDLDUYHPIvjV
09oXCJaDfcYLZLchbNMbCa6Wb/etW16Mw0FYqCgZoWninpt9e1lAiZgFMSUiCv8lTA54U9t94KAg
3Mti4mt6SLS42AV97XDpTZ1xiO8KMt+46WurfVzIO4E6KLXco+bA7h6ApAfIMdjrqAgk3Ho6T+sm
iF2b7ANNrgZV4uEMQayFCug3ojSx/luAPh9fAaJvKX8G7j6mpcHKsjD2Fo3Bnt0K1eX+OMVd0yte
G3qm9GKdAmJr0vIvhfsQF3DoclydTWEOesBXA5rNFKSLnkPf+z8rA6isBovv51pDAqv15IjMlPm6
b0kmxrHTgIYHe87HM50exEgcejtVCU7jzfGa7Z4KkwWy08oqiPL+ASnAw1vJhpoVdjQkzocyE93F
tJKn0KQacujyLfq9KFI7biSrcLq0C0r9iGBR1j3gfqN9+Ysr485fExwHgIqi/LfLRflBXpjmN8wm
Dmu8ewbdugcB7oEJT0bdwSSPuMVhrVuLaO4Mw/D4bBDW0QEzv6XeVjOY8mJTlGijyKMLCeAaTe/O
ucgQUSgc8HfZAK0Zy+QUk+TEZulI41e45zAFG1Gn7qR9OazuN5tAhDkDFyk4m0Sbw9wyNxgtH2Gh
BcBdadBnWBQ8IT/iNRBtT+KIEng6GF+1P2pVGYGaxUM7/gf5DroqbLGAElnIqAVerUt/D/5awwJ8
pq1phdOmlT9Jx2ufd8XNhgUo4Vh1d853rBBFnqk/0Fg7uovrMKiYLVIZ79Erj2a+Q1sYFz+oRcg8
DQAh3zr69wDPswDqUP1KtVK0yXbFTSdKgrdSgMg0zre27GoWlFbQionGs+9TOV0OcdPQiWNz9R7+
r+1ejlppElRKWD23kx1TtXpqfJ/9OncwvQOmTHdGYNUy83gP1wd+wG8mZsKP2ycLY4JQWRo2aBup
5WV0sFsAG1aV25QxYnEy0tNKRZBiC7orQHRjb7dF3Srwc9cH7bemj11QmtOAqlSwLffW/fEPLIt+
hiqDY9OotJ1S2+oDVkc4qjeJTxegPduqPWiFVqoFKZFXVE2xF0IVniUXOqSk+lbxiCDkMzCNyMYL
9t0lpDQiWz+hh7XszoHT6RgaqjaLcIASnR9dlOBFmKsxeiam5nzGZfd0EsEgxdVSE+OfFkhAcQ4H
Pv8gDlgqzRssXYsIyxj/+LY3qb3LVF/kkzuo9khdRhD/n3+laZ7xUGtsVORz9r3ngQa20qLQxQAh
1RdctoSK/De2risfVgdsqiDHDhTyF0YAzXbY18vSm6uoNO7K1s7z7oVFvAcsJyzwKStpCjXXQqHN
QEusZHtSaTt/z6aJOoQw0Z+KHkjcyEH6nmKhSr1VCn9+tmZh028JrpisqDnA/Lf7wQIIA8Q8KiFP
2OA/15bzZEgoxZdu7ufmpveW25yJmw5sviE/KkpQCJwEyk7LRU3ON0LspA1NWDirV9X0L8GWjCYk
OP7tjNJ9oOhQYoDJTIgilsQaKR4z2beah2tpf+dqzJXBxeGhsaOTysfV1nDHPsdzXv4UmO2j3H/S
ZxpQkjjSodbXuCIZ3qrknUCrCxyZC6jTmSO/gd6Ws5A9vFZ8/bh4/8fl5WX2Nl2QJgxTxfUfqVN5
qklEoy5mQmvmGZsUp47ZdmvAFiXRIdFfqk1jAH/inLvhf4j3HwPMk/DnyaGpOmJ0jGgZZngwZ9yQ
lqkyHZf5Fl4ZYp5t0VBUNnMXjNt4v+c3WTTRYJV34jjdgxIdRgAxa6TKKqN4PTNl4A7QOhCAyWwo
cjDxOGjy0u6zRxPweDs94Pjkvd4cLMSLVf9BIL51NuuJAz5WeyAO8i1nTaPT36v3//w7KMy/Kbg4
RXKFkA46p+yIi/gUhwQQhz8LV9/w+Bg3c8mjOyLkrSyRENEu2Mcykz/wvBXe7lZ+rwiVBhcgnbhx
kB7X4+daW8R885MmtQ4M6JQU9cNmgxA2Zif2L3CiRN9R1Jal5wOC6MuRPCD/8u28+nz3dYGvTBW6
haWGlVUCoptLuv2/+DIiukbKW7Nm+mypwPlR16fZ2C95/bMr/uV/AGPLU5aJWVspGkeIg+ZLnBPv
wjhvVpHdsTZPVPWXaqmZL10C9k1Js8lD4k5x66zNfGCD5AYMQiVJzWjEYHWUMG16wHCRPelNZngn
1TpI9zgXoaSyOMR7SPwGhhTaKgUmRHB6SupRZEHUQirEGUWUzPmMQZ/TBiQy9+P/5nIOJHz7+S+d
sGSxefCbgDUbhy3R1QXau4vvhAkzA8PQ01YqxVmfi+NLLQeR/lEwKFUOjjPyar8wg70e6THGrBKS
yGo0m3YKMM5sZQvaEeiDJye1yLskPyRhwf6y3Lk8/+RjLQaxOdp7BECGL1YkcsIRT+ag3DVcGLHJ
Qwtkttn8s1uFQnNlkfVbhEqcT1TsVfdJKlSyvDxIrplftwG+ZEtWfIFaW4Fx+/PvYIfzALVWzZ/l
ymivtjBIEGGEG2Oxv8WE3sSnYryj8UCaLj/kFlgLORKiDgWtWMT0NpaYkFoihVaR/y8Kk62KWLFR
QA0muHNkgaGA9Go6rFiaF8STJVFr6Iz9QyzOAoXDMW2K/NPVccyMq/w/2Q7RY3+GYx5cVNrPT+83
NhXUOHET8LptMjIGq2i3dtxKxLaTl5n+hUQZj9/lI1r3jEH6mpT8xgK+5dMMC+agwno8H96wgt8f
0jmmkbddSzZAcXWzBP1kwzjoOZPa23LDxly3d4aoitC3FsWIyQG8hkdd02hdqqpp7cXxOQ00NqCa
YA8gCdZGm09mR0a+hsayuaYGYuuNJ/BsV2N6qv6PITi6lkX2PtwGbySq1jNHxr7+jAsBd8F5CWIZ
rPrsbz76d7ODqWnTLQ8ngxyd1bR110crA4Uld9DhIxEQ+vmXtGFPbZdsGyyyJLoK6I0ss9gZLVWw
53/8BOb/sM7MkO759MHDEyemnRefatCNvsTGUAJ+g6J7LNYbsqzJc3zyjTKzLEjonUuGVaOLmlH+
/ftgKJlHOQ8/OdHyvc3x9+QI6mT0OWK9TSSvhPKSNi/9hxRhfuq0kijXo2kHIclDuOCLn1/TcUHj
/DKGKO6MiAJAVSuzfWkKhhBgaBnAaqrRr1Kg93q8m5WPBhWC0/NJahFb0dsAiRII6LhEsfbMOFQ4
oY6wxY8ew5I11BFl0xcZfm4MOHrl6T+NOhVwwSwwqqv8wX8B2sOoPoWC2lW7zZ52W9puiwcsOWCW
D9KCPpBDFpJAOwk88jqujQNJiht0EJXZALBi0Dwyju4DMpAS+ei9l2OFjXCINxou3kNKQStZMZz2
5q3jAIb6PVVxRwgLnBs+QN3KWpi6pPGPtY3YUwhX97kg38jWQpkMqnyiIGDYa+R4h6njd6bxPQBQ
9NcFn6vtIbbvnk5k+G4Zm+RdtBLRkKYeVeEWuXF3xzvI4htE1wsA6hnR35vMpJRnt+Su4afuAwv1
y+MHUwSgX6/poAoizn254Ig8zMCe76qJsqUCJsCe7i8cCV+OpPjACle2BTSmbL81ItbmKktYjb83
Po0a+vVXvgkFKlMWrrAjAgG1iZx6B7+f5JvTRa5HD+LKSuotHdnYwGPKkZkdecXA48WnnKiQbtWJ
39KWq9qeMGk56wYK2tFZV10uejGGx9zg/Irh/EXqrF1F0azj/E3eYSadQxC5/Q5Uc28m5olGVFpx
AbgXKelM3utuKcFtJRAN0TUOvwBih3dVPeUT5mQucF543WtQhmOb7FczwFcmWGxrRNau0jRpMJTo
Pw5I3nXL9dguKmSPb6mqO3539L6Q+E3ZxGGEuSDO1VilmOYG8wWzXOZ6D25bTC9mFoB9fJxmQPna
9ck0/4A1kXgJ60KbAAgWey+6V2d06lcPOF0ttuWiT9OHHRjp67YlOpyHsktVbRPh3lh+OTJk+NM6
2R66eKLbQNQ2DsGf9P+4lNmvvnp02gV0zXHCfyjuhUlhmfCbdN22Q/FbBjTuFMQybmHx6TJtOOfQ
2ZJS24YCzq9wUHFMwVAWwnXPCTuUYORL6sIWayEEZhHRG6uvGFmFprPHqR7J1/DHjYFgwoRrrH9n
JvEr1NW7L1J2DUslvtTKEujHxcDNtpk5Btiz6kNWbLIvCpErvhw7Uo39CEyAXzGhEx3KYrqEX+/a
ijGc01MH+lOMY+9gxm0LgYt9rtoCKg08PkiRJmbWgbqN6M6WA0McCjcdWiqH9L3UrXvAaSfWCJWP
6mBftkKUeehKt04ZWeFZDPToCk1LLtTLXoxT5qKB/DeZYTK2G6L4cDSKhkdaSSDp0cDcXuj3Liuw
Fu0cPS5pSxyNPxfovHLx7V5R27+2xyyfzBb1YjOuvDosMWChwEAEDAYCTT8E7OxsWmv3647lpYKW
rJRoS9L8LrgXNEFV9H4YxukfCJ6VwYc635ybj0exS6ITWg/OMB395Z3P24fV830K+ReX2jl95KKI
oDFNiHCvqDBliYwFzmWOu6+HQMFL3q0KuwIrE4fseEzGEDAqmPP/EAsaf6aP1EuaqrcRVOAHqZWb
a4jNLBFTVp4rXySC2kYAXhxRNrhsDJps2SVPz7ACAUo96qGTr1BOQWyYjIDFp0KNTAAFBSfagU/o
Q5WbM5SaWXsL52ZkK8bCeA/TgmQ+X9jQRYwAOkl0Gx7+08tYgFynvCpo9EmeFkLu97V1I9FVvzpi
eAQ2ZI28wRofWLMDwyCdFl6pr8cMWmoLZi/WHuY5oHk1/EDrrKJmXqJrvPbTNBSAjWR7CAF8BnCZ
uyBWOqUzZfTlOU2KGhG+rYhEP3f/Ti+5kO97PMKZtG7Rb8Zrtp0knOI7Wi31ttFx3z2ZdkmzbWqB
pCMFAbpqScaysoy6TW4WikZRkhI1FT9L2zE2sYWK1JlVHH/wa8AyvxYzM2NIztB5W0CHF3FRe0N5
E+50p/lXvHRv73cMMrtkEW0IBOTTxmOyjZw/tGESshY6XxseO0CEFhRqENVe6qDOS4TFtxvms1r0
KcQs/VxqjwDVo9yh7+eDMq62Sts6Lm1bmpcjUcLe9qUt1QjfjMgsOJ+U3ZeONRRg/5C9KtMA68SX
C8bIlOyV89agKcvtKsdVBKLXL8B9Zl2uy+wUYDoF+QVX0Fcs+/IzJk5195x1lfOk1paWahUg/HJx
h/VTRzokDzzxhEj7oCd06cdfS6K9/sz3Ft67YQpndw4Sqijw7X/N79vRXfIYrsUKZ5cg4WH70063
NSGrUDORzmY6RLS49XGOihtbDDIpPVy1F7p0Dc4wQVCu6ArybxXGWFzutVaRUc9h/j4//szYwyGQ
w7+KSwc02JGE6mLRJYihJGBZbUnrII8POWu1otFk/eUxrZvxInG9Tl/ygj4I+2b2XmgLsOZyzgFj
ncQnIgjAoUjL3m7fRZO5vSyap7bf6Tcjo8R7Cfh7EMOgrmuyovakWl0fOWTAId9yHMzrpQ2Dg7qB
V641S3LhoTojtXDcR1Yqy4MpkQFtNar9lMVyb/bwjOvu5bMTIhX9ceAt1sja+9DRkViJoA0LFRWf
C1huQ6A0N4gpza+9kuMVtMxCP04ESb02+1N99yWIWYFjYPwc+3ZcEfBzHB5ywcP/tKIfWvq3J613
KAYE7Vp5VoG3JQUyzZnueoR+deRqScmtoC1esGjOmyJnPg4oOlCKo4MTDQRwWt01Ct8iXCGNBUOA
IS+AkUEQXVv66g2H4VUzGzLXucZVSoqtJy04CEOdXnAqvkplmmclX2VTXUiwhtLu2uJ/WSe5ATeP
c3TnOkqhgbfxZpqvP4Qbnahy9c4sS96FgvTahSYgnTci5CRbzr3SHVuLeLxOV5B/2LMd50TNW5KC
LrPg1Dw7jZHWEwxNj9HShmkVUU1NprmMm++Jsx72gXsfWk7nl17TkqzspnEbRZ0u07VRuYbR+oMQ
QHTCZlAl60GM3Q7uvXcU/9IDxV1mtyCw0fxqiRN+pbnlEtvyvFExCViD8osWatlDdMdfZdbdJtli
cm5tu1ioEyxC270iIGKR6zm6DlPIhCJYJvSYCvLOUQhiOq26RVnyzYbQHdY9DhFiwEnY9jnaFvb2
qA3gREH8LO/cMvBnfNmrM2oj6e02B1b8CpEGdS/KWqWdT8xUh4waNTD8MLVDpQtHBAwuOys0Flp/
t1XbbbNp1n1DRIwxHbkmP6o/dkCt/HOJHTZxAVr/VgF2mc78vi73Idh0BJ1YxIIRXL8gdKhvJBVB
yHei+7SEYAofIZ8nO5HH4C2jeu6N5K376X705pTS4GKx+VbYRrRGxzW+l+LmBbGRsaqxd3XJF1zh
zi9DFxogOe/vCD7FktBL0eY+cyabnK6i7GhMzhZv2TOadxsEGMdhA0QOAsygF60SjSQ2YQ61ukCx
t/7evxQUBzbOa9l/fpl2A58UYcdUQN4X5JXtuaYqpA7AwmW5NotnGJ076uAHcBJV/Hd0E0vVkAA+
u6EwDgnajWyBkGH4OauTc0400OLijFo55EgBIB6Bft7RKSt4xMxRW656qc1wijKPmKO992O7/zZI
KvxTL7mmiv+E58Qq77JXy9Hn+fMWLfp82J/0pTlwNu3uKQPFafQWNxAQRX3fnmbaR9joOVebVJLr
rI/ZYeuIeWr6OnEvFanrashYt86OXzvNLI8CEW4L/M8JjUOb/7zssF/kp4JHlBRTPeRBmTd+w86N
DdxjGYmiuhedKiDPjNwg9+jA64mUN3D/+v0HBeYYiLODhWqH5pKVpL/NHzHsAwGyqbGzR0BFHJXI
fxMckcgMUzBPCKbM16Wj0OYbgvWMM4WhtOnkrb1/T6jcDMBmUlgpqfpDJmlaqyAX/p2JqOB+BZZ3
KIVao/bACePkK58L2lA+NCMLAlv/H5nub6/NqRpGdU1Kc96j/57ini8yPFZtDd711K3g3TXdGw7U
U2uOnfZ7Hr9am8WI1PKkMXDv9iqiOKjwX8p003GHUiTQ/GiKv2ViI17KI+0DTkhrBST2LDbXPkxM
ZR8VB420g4EpeA0/7vsACtsbkeJzKW8uCvIesGhtTtl6AnOxWXF9pKYumYv/ZN9LYa1lQskVfNOy
737jc2cpKUzWfw/osu/KC6Dr0/8cj/1pmWUg8Vmew4WJ7ov78w4XL39YgZ4i1/cFlxOxD4dABqnd
/9rJV1sJyqPHQ41QMVDV3PMIm/6QU+Qsm4S9A02fPwreP6ZyZJ9/MzdzThydxVm+CVW8tTPDH5FM
eLBjCysWRurrRECBix3/fP+/KDZGrxRdPnR8aqIgPsBiL1dCx2Kh1aXPuQGCMtGhwlx3j29qKdv/
8PViqGJFYTKuTiol+XpLdErBHal1BKEQRcHo4tNGmuu1ACwlolWcHT2pxYdwvSu88pHGzAq80Z1S
bT+4ko4skjRJFIpV0xEcjrtO/n0IDD6iUhWztm5mTdmWA+miC6rNSEgJf+lVCR5TfTxLpmmiqxlP
N0EFDm8RPxFZEojNqjjKC0blhZAqiTjWpkropV/6XmwlyXNoVVmrK1izKS592FJW/htLamGA9qpN
80ieDlO7iYWd9fNeuTM7UEGwpivBl0bcmIr2TmG5JHfsvytr0tUEgSkeXh8TOWuFNgmLZHEiSYNi
g1woG2rcnWTXNQqY9C7KDTpgi3qRKrTtCENlsI0eE1YvdKVJ9azfQav1lrPYBtrasBh/5krXgcZq
4g4SaWwbWHWAvoKCL3NXbWdADV6CPHTxgIgZfAA+tXHMrNdpUUwJ3bczOkKMlOC7C2L0jz286ngT
o8v276m6Yg4Nv768r58d/a/9R73s9VJOMY7lYKd3jvBmYshk24FqxJvxe5I9BACRXcSU2RXoVfZt
RC84+1F0zimCFxXpCpyIrS8WcBfiaNaX28DigO+lrYI7djQB4XlDA4NANQSLlUUcX24lwOm/Pq9I
jdG0iL2Ud7QKAadoC5AnZv2T/ozlMVfD8XS9ScLHHB/Tg0hTfS9h9Q/iXJMsApYBshDAfKK8xuox
YuCX/SDAcFSyx7QDqzn71XAngqUcbvoxty1HOxN5qF7n/R/1cAQfhmpNTOMZVFZCz+00zinTycCO
VtpvCWXFYgry/lmTisVyfjPNTPQqymeuDN30HA2ZycK6r9ozSZW3TaAGNhSh8WSpnFojjNm0IpEc
mwiwZCz+FSEMsHA3diWj6U0Zw2lVlyJIyETTRaurnGkdCWDMc3phpnv39SxengZb1DlOelJpi81T
pbeDmx+MgfKXy66de8M6GH09rxuq65n528PB3TYITneLIaxQRTJ++NfJQNgxQPTIZn7nn6hhllij
VQoxc1XpLLaY5t4CMbwDvW+Yy2wzjKZbzlMAdtrpjG4eeCbndGuArd2LjhizMNOnoZJHdqdwfIpP
EurzcylmV+A/DIjqMwdJ6ZGZ90ZGYZqxII7YM17c4WwutmTh/trIzoJcw8nlH38V4wk0a1uJfb5S
aDDtjgDI9d1bfoOeW2gG2Lc8HSLrBYcfCAkdqZwY6Xs2RSWLH7agZbyavCOoWcodC4R0ymbFPsnt
2Whwpb2kWtXfI4rouk99KNTwBN6DakesmzjksJFMivMWh4kMM85qUkVljXwlif2mFndzjs8zV+Yh
EwHjh1wuPcs9tZp/Xyoqcd/WGLNTCAZz784PzJCe2kF8KpLvLAuUTEHEkyrXG2AW8UJEaYxx5aIV
SR8zbQdh5J9ePjJPlKtuBg79mkbfNYKhbIK4YoaTD8VpXfViKXEwz5UViGyq/Q8xjmJjg+pzC8nL
6+u1fl6ohOJhcCfGaiLFOvH1hMGx8Q6jxtEwhuc4l9mcjnZWHmoHCtjD51zDyMQOdAzb7sSj5aiC
Iab9twKtrsy0ot3f+EFmsX0pfs6KP+Rbb0TdBHcxMzKvSroUlGj3ozal1RqThlEy1jXmn2r+DFH0
MC3cCC5+QYW4hgwNxW4wJhozLDWyzJH2mV/uo6PB/fSF4c+cvbDxaZ+WqaAKOLcGXjzGEnx38W+H
fCbA7DZqBRScOF5O2x2mGwLYaa5/YQHeYsmDL1FDuV11V2ZRdZmsNlOnQDgzT2pNDwouy2DKfRZ7
RtuUcTCzgJOrxMZFGI3GM/XjM27JkUgsO9SVyS4vHEPCqqvNPQ2DiHL0Tr3rzKvVYapdtIN5L1Mu
/PrRgKqbhxhMUKgKTLCSaOXQAJjIAhZ+OiubSqxPOB9mAq05Bcq5GB/q1HPy3oUHtWewkF2MH3fx
kp+3YsUXRbyZyzM2bxfWtwQrTKlmdXe6jk/+iHMuCucN2geE4ZaeZsjVAjHWCgxS5fNV9YvJ1BBB
zFig2wGunxjiEdzTcgvvlFSmtq1N3vOJtpHlr/RAIjMQXHDXTHe83IkpC/OASxE3OAdRpIhXUehm
hSrEuzQQPxBNNXqyl6WdraHWnLRioCHUtHSOXx73HGmNz+Z4E1fscV+B0mfsXm4n4UL9za5b87F1
9HEWVEOTLFMvhnPAiVkPvbb1oMXJsehknqlcIL4JaeR+ZuZKdfyFk0zzepVkiqZDhAU4MOL9Y10+
7ChRU0n+JMFomB//OUTrH/87/crnCGDla8A2oeGDsIMZuaDdLY3eyFcKgYf9Na3Ovl1mNxRT8b+D
bQ/8zHw1GF5p8VyqiBPrIsAh0imCpo2eLr6u94NvLwZ3UZQJI2mdtTgGXZlBhlvPHPzZ+XNc6AH4
zp67Wahxy3xMHdFtBkiYIuQpbGsjx9cRP9KayzxE904slfm41dHRxz0U/FQadIGsY6MkEGNxWTqc
RRT0xiE8ZKKmb9+JAqeeJeR3ai7YG3/DeIoixNAIrvbWCcJ8/FuX7xt9dQQY+GJeRljDmxjURQyY
OLeMEMGZsHBhGJOHnaFe9sxPHmcLZ1aB8SQyObZj6Lo2Dk4+jicMa31w65U2qCv+U2Iqc4A4XB/h
lgmUK4NkSajovx1kcr93u5tNyLLL6MxlZ7w4g3mftIxcatMSo3yF0+/XRsdvNXlDO+G34HsiLtkM
mQsdEFOR7yrZ2IREaFSRCC9k6g73urOzieYy7po37bFzeNT+EB5PX3InWJ2pQEvI+Cboc+qEnUlk
TRAikm0cjluO2PE+i0q2jqc7DyYD4cKgjRUYQETf6oVtphWfRAmky900CNVcqXPYDyP7oXDFgBhT
JZnyndHkt9pSHtTfkIJjS9eyc8biceozLy2Bc5aF/zc8ohqHcdNmJOX6xpfuppe/lhz7SHoTDyT+
5lEVyaybahZt67hZaBiN5PapLI+m7MGymNtaTkrTyV7WU1H5t4slVTjbWDSiJHF+S2YdJNoOUysq
Em4TDJIXFuB7DAZDdPsTzdvKp7JD3CcbarJ7MaKrwYqEtwWFkp/NQmDYNXAJtWFjrn686HurZxUB
9WZOmgQPRjVY/dhM8hLfiB/WmuK78I1eNndZztBxmVgR80cNhGKJlpeW8frWwPs+cpyaTfeRGq5b
4O35u17G0HDeRvKN0A9v7Cu0od6vrR1L9l0WgXNm+a+m/hR7jarr4YdlJ01ZhjvMdL8N9wvtTQ5V
MAwjCL3IKiepmxlWTbi0C33UbdMMVHbYCL/W9u59HN/5/Tl8b0nz10I0XnOzxkodt35R9+SxpCGH
rBZFLirZYgv7EJ5nywpgwpF56Ieh2BabbhRTJc4t2xnaRyaxbPaagOL/Ecf+B2fAp/OjvJ7Xj+/C
fkA055pak2F9br3isGZCUuq8ohQu4wPV++GPBU++Nuof+URWdjZ3h0USpvQkaqbltZO6SyK9NwgL
+yujEx57DHuFUWx4B8TveZzqFUB8QpyB28CAMIxRvsmEePdi/gNsYmsHSQK4GTLTqzySaOFdGGA/
HhMsIrA3LVT4QwjajN9VAa6c/ApLQ64dhxOWmndUU/CShxiU2+PpczXM3qBP/V8kGcV+xAe72u8+
z6O50UhN9pkyEeFPZ8AjtBOjMW1KPrL2lDvgTmcRQu/yue/y8Wj43LLRheNcMtZhdWaA5pU2v7aS
lxTlergCzbI6FmIjlSONNKwxeyA45KA37hka19u1pcFfCapaHlPF3Fk7Av2LLOQYZnQ5zYYHa2Xd
KBDZgfeM2kj8ZVR2agwwHXZmVcIhMaBbBL4dNZOwXgdbduVT2R5cT9fP/+rFwSaQehxs2iirAx1N
3oVrgQJC4ouGLDCXFpEAcZUawJvvO9rYO0PMUrBk61w6dYUdKlPWuhfKIQPMKFgokWpX4hMrpKlU
MEJf4tUl022xQiYYgchKBkZvVfFMn2YAa53PdVtInK/v7zDAWwWT+qHsccE7+NGER67a+HdyUb0S
D6aNi7eg/w2y6xuefAK25tMohpPZyP8ISwTKqU3rgZddlCOg0PMfg5aiM61axEgn41iSqpM9bRRH
yXdy0jL2TyM4cp0uQat6puNF5uNuCNn9AMwiuy6YBzDw52yaTwvA8IcwlOYqQIYcDZBDp5vNFbAs
QdVePyodIv7Cyc2TC67JymMAd9GHo2ntJrjuOOrLamOrX8BdvWS9GmzXeCw2waly6jAWuYVbhD8c
QRqSUc07AJDKuqoAIaXnMsqpAiTTybSU5Ta2d91Q5xVPsyOwDlI4+7nPlPWFcKnnaPBLc8+KclRL
0Dmh8ptL3gbhGAco+kRIMEyp8IkXIiaENGwOmgb8T2W+a92uSgnlnpIcHs6d5ynTjl8nyHQpMaue
j4qJ/ywP7mULM9g7PPfZKwIkMJpLWpO+c8lo0wUXfcsvkODnyt4KjJp2noFqhn56+5z1CnDy4w18
X6j4ryZSShZ5CCCdpVJ19d/lrq/Yn1N7NXdJw+/C4aiOPilK9QkouL3/n5diFTFTtpVlCPJwJseg
2IgF9cfgVZJRxYFYaXClMcNSOG3mjaLCt4AcdEa434G8JzgCufP5OQmBz/hCah8uuBGB2k9gpdsw
31rF8vYUvf4/qNNORKXVOcoJFv8s4nPFEmyu+7sNeRYp2oYb06DQu3gGh+DOjXJUPwWb3Xvn1MPz
OfIIiqR4waFh9cUuB8jYZVVAzxaigz2IWCxGv5U3D490j4niVW1JQlkB84ii4Cj7PyDl0h1FnDU6
ZBZo36EBggPGfL/H8u+dax5MxBcybd7wG86CZ4w5cousMzq1Fv3hFVOU1q+GoQlQAIK2GCGUxx1/
hu4IKBjN1lRHPY+Q7BphCnI+kPKPDXTGAZxQOJNoSjspMSXQK20btulfS2IjW5mFqAhqzuYKyUGT
Sp79qpXGMMS9PrHDEq/0fQnbgufm4L3XbdYco+QACj+WGjbxbxdoP/LRA/a42JOSq162Unsq+i5E
0RmfUoI7DGQRW6P/aQCEGMzquhHOVK2yTkLeLqIFyq3w0UazNNV3LmG56I2vC17eOLQPfRAnvTpg
HkurWxL1skHHHKhuCrq2JwH2exBz5fGawhb60Cc29sWVOj4NPmEmkg+2IyzovLtYRppHDHgfes7c
8zXHI6EwHHMv+kcc0Rebw7nnRKPlupJuTLDHvUnZBpWiB+WoucFX085jNGn46NC6E1tYuj7epP0G
ojZGrFflOyyoqByr/VWaAzrvLnqPe6EqGvuJr/T+WXKYmelhVqV4wuY7QKbUmxN8D/m/vbnqy6gK
ZnnKfzIWSexUIlefGCt4WUd+YIOCl2AKvYhyMIBjgjt86g+77A8F5NW9bDPS9KGuGwNciiloQStU
BMEAXJzrxoYRph2ygeZM7ivNHjLeI1ZfbunOkPWZHLKBEH9KKAjmSgD0j+1/oOmZh8bEq7SXdhMQ
qkYfow8UB5FcJ5nXODmedkSVNU3pDTJ8R2lg5aONTZP67opsIFCWUzuqUpaCNqz8R8hyTqkuomti
5w+iySCmEK1fGjDYsi1vXJrMTIe58YiBE5azfB8spGL/sbTHe2hSG6/pnfIIPuxsRj5sgq355tip
wmK5Cbl/BKSUejQHNRb1BL97mVFOmVoFJkO4LVrlDTNXttRlpCcg2mTfMTskNuI6lzGyJFBnWyag
DvRASHWYkpUCL5RCdXcR4Z9+FRREs1wjgGpa6pj1r9QvzaqZwFAWiiMRdiwxt2+jbpQBgq1vsoS0
MVmNQseNopgeSXnFgXvOjUIKn39TU3O9mlauR1/DkMgrZZg9dQWhtDETnY9Jr7GgO0UHkuGttVzr
R1Rjd61GFUwC+63iLr1MpXJk49jVz1ugT7Xh+8vGhLY6+bbcLz+WKr/GOXFfPGKxNk0dmgyrQ88x
BqSXe4sZJ/TNuzhBVCUPO7uWw358moXe1ocV0vaJj+uwgZXfiRQDQ8fvoKnQcVwsKTxLCVXqIv70
iXZWkfdpSyZhL/ueys/WB5GNyTxr7o8xHiIxtfM+JaBLP60XgQUdC4RJHlzN+42rysK4DBrVuxfW
3UZ8N0Quh+5ffn1A0WLfE4WbnxmvjDPJM1h0lx0/KrMSnCZk1H4fdPPBBkJtw/5CVhwv0zor0H+O
8ex5x3F6UrfonhLTa664soJtblIVhN4/7UnxEnZPTGckTtw/TRJEdbWFUNrIgnBswkqY371vE8Pn
lvnlN+OWayvQppjzjFkO0q7i4WpWEjRZg0ABlmR9HBqmIkANd8WLhBfrTbzRcOFsNzRo+/Kx0+H0
QxhZvI5LvzJBcff3MCGChQjxoLDN+PmjFQzHTxRQ9Cid6ckIw3PLkmxabSQcyjjPcaq69CdxMfqu
wyh9B92QBWLGEcYjo+GerrY00Jm0LpVjCR4mTJ+o4l4lmuPyproDL2OyDlRdCVHsgF433UTjjrbU
UG3HrHos2XsmdLqi6NRLym9A78br1k7Vxl7wAuhmqpWK455GN48muQT9dWs0VG7NEhVAmqn1JWS2
e/a6dzcTV9NVfjD6sOB5d2XHJ98u4lGkwPINzoFFAjw7NFSCdPU7XWwcIzTMnMLItS59b087zu1Z
30NKnS+YIFWg5vnxxFndsEgq39xv5As+cEurUFJJDVMh6ygty0z7mDOkjos+jwxCaKJaSfTZQmen
4m+tJ4Pg8kB5oZ1Ab2HvNGIB/tJCqRMqsULk3T6pQruGROvFeQH8q1Os+sZ2+7zYD3H6im8SXd93
JKPzaPIEm5nJboL3mSCTzIwNj5fhlP9AZE9OeG2Ca0fqjFWn25tSn9a6dU5iODa45E+93aRqFbRz
DXoeeoilocKXIGrJYCp2ZIiwiqbr5KjSqHfxASIJ3+nQeWLZWcvUQlP3KYun3Qlk4f2DLNzDxN7Z
oc0pDZyWF1fI3wkZv2crRM4W++2g2Na/OzTZZn8oGOSs8JeZX1EshptLfph90fKkRaaGTfnI5uQx
p/66X9AP9zWKzRwXsvF8vqQBUAyBMar6TQc9h/CZhFWwIjjcRjzz7+MZUmJrX5gw4UOcaA8uvnC7
D0BGiW2AZIa4oVI8v4STMjIeC9GU1YU4By4LYljZb0AoZXtpkuL1F0bDXfi8vP4yGuuz3NU+JYeq
h0Xgw6N3Nf1dNpDtlbiOdJx+MKkSHYaWwTRRMkhxP9vPkZKfNDX/0kzup+bQeZQh444MeOf1s48K
nw/cbBveA8zM/W3J046HvlGCf5C3GSCQeyLfVm97ax31CtSp088inpzWkWGiUOgfU/uQzvJLchsW
zOOMHOOUKA3x0xDkz2DfxfQfi+3bo/806Dp9stZSQIezx7Bx/oU/a8uJADbPgzBk7wHZKc7qTv9g
KY2Gf4/7kro46FbLIvmbVt5UycGA6arw5SlWrLZcnC/SXR5VbrkOKTnVG6nqEa1Xxl/OblwTbJeJ
ox1oJWZa07CqrNE/WjAbDZTLfITlvE1o5PNpbmt1P4wRyAy9p20kRi/lEYNkyz//OjQjsFIEHLGB
sRhulWWq+SU/X2sL5W4/poxDmJ2O4KylUdUrt83xmKxqn5KJRBJsOOuA1At1rTQzdayeEAzZz2do
TOx8VNqHESguvbmaTst0kw9olWI/c4Lmz13yQhw1sS5A1hN7XpBp2aj8+bhHW38gUP2YcdtVFDhX
tWKA7oNrr77Z2OUX4vUPwkMcntDYu4szb8UKmRAY9UfKoJ2xPtZQqKzHrlCCC42Jx/xIAMMwxxEZ
0zMqyq6nyo1krWzpK7yNZ+4b244R4cE0lUt8X/D6Vag/+ghsnvaiUZzMGQTG0ZVCTFlyxPYxTpKx
83IsVBjlkxwrIUpmaJr7H0EFOjFSieaG6Jkk9HYnl5PhOd8o8lxCNEbMzmN6fP4PxrGiGt/yGOHB
VoUJJjkp5SWL1AC+5FFSJIwMVvH+8oYjHh40S4lzZai0Z0jBjud/57Yywnbus6v09zpdWNv2LKEP
0t2YhZfOOg2bgjGgK6JsgS/kpxWyZTLZ/BwcaKqOvGGrrfy6ATCAVo6HlkcE00vUfYaJmTO4OfWm
3hznFXUIZ+nn457UKlAMwkm5TR8BkaXG5JyY7IwXCcZF11GJoPCD/6ktZh3ttyCz9fbAln/KzKI+
ZFbsoG4AtTnfiUXl+Ce+GpQmqTgJIRhWFOhlOaBKKFiiuGnxATvzzs7x3BIGZdKDAjJX+R3hySqP
a0Cv3qzrHquX4LqlsBoL97GXuQTEdp8r9mpolo1SqcxA4YkcX9u9L7vKzEDJ2s6t+ajSYlIfpC6G
AmJvEkP2MzPY01iRAVDTcYE7IVNSyw42lEyjalZNIRkY8bK5mYT/R4ZU6gX/iG/OF82yl7WmGiB4
JMRgjuFzJEi8V6PGL0K4MvBn2QFmF7jp/d+tJrykwtPhny7NXRo5yAVIf5Mtn0y2Ek0csjXvlYfh
ZxaPBUBfCUdHX0yzJFFqVMcH9TdzEilDd4mXktQhD3MZdH3nDrv1GXm6fNYZNhD9OAL7nrznYRK/
E2af1s8VhNo2M4ygaj8RcXXMvCs6CqyXzOa5bUIq1g0plnB789CVo4OabdejrDN/2Ic8wAWJN9R7
XS8tVZlOHrLeX3xbej8y6OdNeHq6uqAGp066p/J/YQcjK4EdaqFy8Wr3z5CecC6E1bhssutjzHMq
myuvsLQAFY7ujvzSCc41SDflDtYom+66Fj8Vlczfv9TjCG68uI8/zCbdpZrhuXttLDWmnXeMzvut
6n4Kqm5UvY3Cgw1hicbxDr7I1IMwaB16wt+KtW0+QrSy/jkygIeQkH1eIf791LVQgQHf10Kj3fSU
iBzxVWz1UH3D5lBZ5wFCWFE4BjnJ18uvh90+1IBrFTTp51k51sW7KNI9eTgd14MVYW0TLOugXjHM
OHFIDbGRyxBYGoCBVCK5b5vW7gyEGyPyN7TqwMLDFss8ngXO1DgL+XOIqu5elIphJsLaPYd5hlAK
BBJOaxuWtnHLujlfQEXIdm0MhwTJ4ys3w00oUiEkcg45/etNO+HtXptEXa/tgTnDBaEfQb3lmH1t
pBGVWyr3f84Bfd3wPsGjMW73EF9fxcbT7GzlzgLDvTVaZydQGw9JiL3cduWb72FmsqqzS7r0Z3z+
1GODsVhIuJKRujqVPgONiymW5WTmDNg8CextDHGQlihOd1pnD59cDf6EOgB6t+XJFy9asm91Ujrb
MCkyWnLdB6Fx7rRnniA9m/Mv0pU0EI1AIitc4BuB3J+XLtn1FZd/qiHzfodM4ioYSBjXhvJHGO7e
lZiB3DzHFKz1S9rbeZ+fKk8tk4qheSL4mW2uHjCKilGws7Eu6sd+Qci8nczc0GcWcaMedxfQwd4x
JfwPPAPOhSLb4dsU/dSGeEzPXstD+QM4OjvEfxAWYhfQEVucXxsJBWx4FBAQwV+GdXY5vsEtcD8E
5Ud4n2zJQ/g7GKjd+FEpo8MKro3pEWz6C56g5VRSZxD0aqhQBVXZyESxRwPOfwbbsvjL2mIUz3xW
gWMWJ01ttWthy+tMimgLyVqiR9DnIVsTLdvjC0MWvvnDSVnO2CM0GeJtRL7kSe3149GuM0IAEmXV
f0ow+rcI5gwyizoDYnmI0TZOcSYI9q9ZIX6XwH5Zyu3Uv8AatMs1HX2We6aFvG9uM9mOTLDBP5zO
8CzIh+ivrv5pcRm8k+o7Q7c2smPx7LmsVUPjOMGg/vJtfsnKImbMtNvuCAOoMy+YfpLUjVm3vGRQ
irOzvDtuRUSjSVA6WRgtjOYMejrqbSSpMNrQvLo0kD4pWanXup1sxxhAbnWrVoA34hMaR7PxDhTp
faCz+5jtItMOeGJjImcMa7ALzVkGEjqI8LdtQiSdk0z8z7/bCEraJaqmnPgYRiCbw6e6ttvRV1k1
/gyVMbspIY4TGq5SPVUhx4SWJiJ09AKXwj1YwMmnOgOW37b9qkJMYG/MZrLer1WJgJoznFYoM/5n
5TxvW/lpvWgOLQogINpYbm+dAgR7kd1mhHnzGpdcDUkUM7dpI8GUTV3qUJ+tZ4CJbFATV+wBYeKZ
xCB02TvyxE6tKSPdclpN+ykLmx7npTzTy7as7o0LGfrgF+RgtFy/RIgpkpyFEYlM3LDiRMQjWV8D
8t1kOJakOssvB9f2ErbNsZ0y0oCEW65N3gcqTimpspbRTEKvNqGAaH7LvKIHhqHRrB2m4EnSsS4y
5hqETUVGHWgBqrRuezj+tQss0yNjalMPtpBj3lipALfVGD5O1R3Mp+hk9CCECGTjmyEbk4HDc6Oa
vkQroqWDhcR4xxjN/0ItQRccfcNZBTJbkSXizhGXMgxjof7zfjRwQGOX+upLEmfFNqI86GMgyQLJ
MsSENmMOJWDF/EMIju/FhLmnd8oXl5kELl52xQwF7HrP7QRWtNBqK9zkL/jqzQ3HUnoMYQdmoYzI
PWblcTzZZ3KwzicsrAs9gkDiWISeo/bwE4/8IAL8UZwavyZurEzADHTU7cQ0J4hvYY0CpXbMK2na
y1tTQ2lvlEEaDtolrF76SO7a2/8Jk1YjlQpqWlWBQS5gPZw0jW8z+4WvQtUqRp9VZ07IFWMLwvQX
RSsuLfZcPJOs00FxYJ3XUENomxnD9xJC1Ria2Hw8C5/ip5SZPkHNSTrgL8TtEcsIaPot3CaQlEbS
XVkd5eEypaeyK0JvupgsVxC5cTts0WeOqFMVv2d9t4pd63Iyuui8+Q+59TEww2lg65Zx8NoCybOh
A7lOC6wd5TjntGBXCyaOfuLChJfOjIfi+ZbVRXpJMS5eS+TxbDNdn9ArfGu8S/GRPADRyJ04JPMb
+y8lpIy1k1TJA8f6xI09SEdqPzktV3ZyOascLgtXwrejbfBdnEJww3l7ssMKh0tIRYGqdToUNSvL
zUUzJpnfNebTcID6XNJnIsudkgZn+c0ogEGWn+KuxclYl2Z2ifE+HFGCEDw/OSCC2uzMXcQ5Jqbq
rVfOTVg0mWp2C3amatYq/RMH9L5piDggpn67M8Asmc+Bw/lly9Syj/Qbk4dKgmm7TZYL/Fp1hvfX
yGADSE0VnPazwvTqrJGXnrF0vHCTJ3FHIMxKgpEg/Rpxxw6uHIV2zX7SisuFFse+xr9d3tXXsVn3
qql/M24GUPcN+HKkXiOPWFBEXJO0sqZX1qWHwRAA0BQnnIM2hbvlL58Fh8SNglPYB/wvp46t6TK3
cHxJRQi+sOS0nUboUcs6YeHrr9Gm1yzUUWALBdDsc4zpCDVaHw5eayiQa6T4ona+o8SO/CM5/ljV
jFtESAzI2+OXzL8LQmk954h6RMDDEbk2sUvsu0jlczZgtVkDhdvdFh3rmWEzgbj3TAoVbknDxJEO
chgF8Eote49s3/Z2o5Flo+riUNckSovEk0aRthCB5PRivGv34BlxTSl7ck/qkGD6SNG6w81X3C6e
ikCyeb71dXTTMUhMN4UMzfcbU/qP7y9oaW3U6DfHFj4C3hBFVuRCawY6ilQ30XYLP6nmQipwgk/r
McDEGRnvxyLhtd3vZwVCLNCJUxJ3MsVwAzqxQ/D2NDbewD1reDTApWSxtUx+U5dPU8eE4A3l4G8r
7xyUzGKqaHwbcYYl0qDjCRwtObOKCnC0n4vGNG8v57BkGyL/kR20Utk6bD0gxHFDB30UisSUUfEw
ZVOFpGT1mzlEq6RSD5D63wYNdw9CsO8dkqJg7+EUtCzC6qm+yT8HyjxbcwxP+tqv9brZKwHMJfOs
v13blKg4FsJDFNFodXb7qLzr6FjPvHp/8DE2RHWwjcVAfoeMT5kD9NG66uToU6ec5FBK9DoZdbRI
EilOlBbIfNS51ta8WMBEaQMNmfd9nJGCZWk65dwZV1KnScURY8bYSLjdDopfuHtQaR1g7I+lMALi
vACuaJuVmkdKx4C5wtMr817Wbayjs75guHSSt0zlPxXaWxbKEt8dh+N9/kbnXq7Vv1LWWfBg1ajJ
EpBGAGCIV1lZARYEChSgwJvdA1ZCoPcVFavnR3hhTbIExTQgEOImKRWfHCSHdaau9Vtcu5EbJKs/
HuKeRUyviSPH+Dhb1GFxwGlgl6ye8M+JsI/shaX0nZMyR7jNk5fSluT9vcTsDYnUaA4L5zjQqEw+
I1DrDG0EiEXwT63kMeJ/B/krLTWXbmIXShE/MwxA+grz07E4sSPgW2aQqN57aEkofb/DojV7q9/R
7eqGQZO4blsl2Vm16mSVKNARglx4+69jkXY1FkhuYSI9LahaOAnmYOOyvVQ/Hy64CiNHpIa033lz
DjJeDOzQCnWF+wC7p1o2ZAja4H/U1/VL8p2QtC5Msp2jBFezpFIHscigMYTRvtv20of1QGJHt35W
5rSbwZEzvwv/rAtnr2t3e3DRD7vp6eBKeP2YayofnTwnRA9AZJXIWY0LK+lIa6AxNMbBYFtrhgJq
YrnP2I1N/YOViyKBSwNbt7+wIbOKAUpU+xqRttoXiP6ZFOhtZtzkP/B+vudDb+wvejxfiSiZvdBA
ZzjpRDcRP7lUp6HMLYWkF8/Rh8ji14HRK35Mr91qvJyQcfDk+TXmJ3iY9vKINicSR3cpm40kQ8Fj
gNbAYZlGYIzhONsfPyNYRs+Ab5wnZZcQRHW0E6buDcY5mqAPlSD5SilWR+3CFDtE+D8Hw8QKyr+6
MOFnITvwrpfcRnSq/z+xRBnZgc0Lhuy/FSjycGoUxvoGOI2I9EK/AAMkse7yJQrKo3c9FiUcuuZ1
j0sjp+mD3nWOKGdBqSSGzv1Qa92OdW9z6Nu89R3LRHkeINrb1+kEH8eKWyZbdXmDoonZFnGmAmMZ
E+6PQow4O/SHIIbh1gWasV/qySGwHJ/k0ji2tQs0T6Edu3n66/iGfPGgiA4mp5wawAiK987zP1ts
E2eLKlnZGbFlc0cgtqOvm2/UZqnWrDUrliAR4wBfLBomGB1ThLUkfuWnY6p6qUu85JiYuhj1pYB9
K9hB85JeqZICxesOajcrNtfX/us9O2eTPuiqiGI8uqw3JCdYff7hK9HAmOWLKp3Z3/4Zj81jTKLg
c+pAicL/kgJp4bt0hB33buZvX2YrtC4DVt9FkYW5erGHDDnGigfdD2WxPQ+TJnqM+MMwYcnnJSXv
gv8h4aykwbNXBlrnL8BBMIrz9VTFLv4Hw47yV7XN6uR+wa2ZScnlZRTT/VLFxJarm0aojKVhZ7K6
sGCIlJanTWMI9Mp4JPfeOBAr16KkEpLyBttcb8+1/76FiiklG9mneXbPFMTipxwhSjYGtPrQHXsO
CpSSSFAb/pcgbUEO7zBc+Xt7rqzYuT9uuoifod3xxMVR6lPybv/+la9EVssZlOwauaROoVUtmzEy
qUY2iWyJVMMziGV2UkTNGWPKSKFKByz5eHqnz9txPlj9gtZVU4jDemKGMsaZlTGti5/X7ku/l3Ew
r6A5ZYCP7/VAZucdqAYgChRL4mO6VpXssg+OUvCXhzeiW6zXnVcCqjG9tfpvuTvxDAFRu8H47H6P
PgekiRdW/9G0I3gPR3wswcDB+NUMxpVND+D8sTzzgD4UJmkbdl07ntPMlCab5e+oUcx0kcu3E0Fb
WXWa45HGTZjAP7iuiTxw2hPKxzvx7U8cZpLghcf4bqueAK3Gi9FJQX4V8BpNs/LXwuEvXbvuxBkw
ihQvAh1YKdw7NNk0glEGGAZbAa9Vl8e9v+0gCet0gfXuBXUucMarahfAw3aSL1/Mi2b2zS5zkTJn
BFzYztSe+VBryhJDPhb2hXNW/bGR/PrnKlJsTAtMpV9FpWF6TfS75lgd04wfSM1XH+Z8zqRv1JNu
ArOT4B8XB9gFfwv0yV00523Sc6gNygOudBqufDBEC889kVqu0j/3EfDIVHaPinXX1zaB91YqUWyV
dhK3dA/EzGyb5hjBhL/a/8fyOlBoe4kIKx7cgiNf8PtVAXpL5yqevLPIoj6yiiOTHXVu6DQ3LcRV
2lsl3UgjZ1i4n7vHLkeSoo1kaH9ly9esOpoIq55nmiwGJ3AjZXpJR+tJbqacKmInT5WbLgBbBEib
PNXEFRR6R1lBZ76Qycxgyq9zE7c+SmUv1GNvc2YIeEVHrTM7JibQs8Gb42NOpujxWJA18kI1xnas
IoVdfby2g/AuM2af8oi8RQok7f832d7pWr5sLKKihvjX4bD7lkR2Tchm0LgdHJVSrvF61uMG+RyP
TEyTZCAMK6DY+i3LrZckqKCZG2qEWDc/Enbjoe6bKPrIE/+Vs9/uppMiMORtOXdzfSTgYorzViIi
MXtX2ij7jTHzR0OLKgYCUIk/nqRYF39LojNBeU5fd9XACpP6jNmxVejjLA3ynw+OgHv6+yq2eNkM
O3eqkE+sbO6tf2LzwhYqIX8MyBeTkIVKI/KpgzHn6ETL/N2CdHQcCdDHscYgwPXzOUOXgRAzMRKo
O8KhB1QL/YGiUfprtXWDgjT+TsQhqKiAAaIGd0TunEmFcGFBOZGhHcIDzgBElHab/yWyTiNOQqEG
TmvOA6SESzqi26tc5433NnpoGSv6pAtRz31wt03L3huVBB2PWALOG4ppYc6TfqB+OjDyvki9ZIcp
0CqQaRBtbgTu6BHx3PQWe2xCF3ZDR2CIzWD9ttvu6uOci1DpAFk9ua70qsFuf/RLoN/rMFzGaxlV
wg1TeR2TiHO5v25RL4M+2MCL7SlXWuY1RYQkBghZAW3bCDEDAicHxlxmyq5QP0GOe65aNXL1M8az
8SP9X90trVsJ20ktkgnJms3rEHytwwOZaPdL2UqWThiCqOKPCZ22rgUPmODV0trARRbWGf4t7lcC
hD9iVLglMfehWS/uCykcg/i/Z851wDtRdUnzdXhmoNwvU8U9xq4nWgzx5GYJB2OviDd9jqrHS1ML
jIiBOlipXPidOTBOfK+lTLM4Iqxc4gDPKdwg5LrRJj8EaTc3KUvQPGt9x76TX3syn0n0jvn9KrDg
XkCSJw4Hm5we32ILKkirXCV3LORfxn/IkisfdxP+ZVsPcIY7FEbZIjv6/VcJ+spTck34+CuLI5sW
kpY9Q92KnhKiN66BABkoMdaYOXGyiekTCb+qfrNkbukgn5wVyH9yV7B6B7Hx/7FpDoUceZKErhhD
yowkYlSXXmfcxCT30+RPgJqF3FUz5tP2yHEF9WSaW9a86TB3nkaDjPmGehxWKFLAIPjgop/sJFi/
xN/0K0ZiTHyw426MwsNBqLLOrueoLOnmH70Ba25wfpP+a/1SLOXOXvjIjrK66ONZKlSDtoqMzVSy
bHiE1E7dgIDUqQ5iwitSfE32IXIcNykYTzShzxkIg9b5/Q6ri21XhW5P/mrnjZ83wLWb9mYUVw5Z
dvB5pnREBPhhs2mJweu6nq4FIEI9Q98CUslo6HJeAqatk2T6bR8+hcWHVuevpB0hiAjlNIF2917v
RL6wJceVMw2aKfNlvmDs4p5sM4UevCANZeowRAE6JCW9X2m6KLd60Ja5WaGK3ljdZ94U4wYdWs3B
TqpAAaH9YKMcED2ecwC1n+O7qV/34dWnW/KkgJ8e6tbkRjhc6Fs81PB+QFYkAvgsKhluBrG6fTek
R5jMkQTFNuSEoOtxlpKqpy3CFvSQm8SSNwq4xOs2ryVj8q4FVwcqNx6N+BNpR8bbC3ikuQToqwwN
DvrbFnVtRUwnLnjuJoyquwL/uFTxosQ/F+oOt2qlKfvrJZZ6hs+Bydt0y6+hnxUB/14Nk9Bwu6p3
/8zHkg9Iuo76pqgtRiSKrQJL/1gklBwlaCuUkfyucE1pAj2tfOhKMSgeuFsXWots1ccHy2Q6Xjz7
cJdPHKdx5zJ5XJwTzwSMxhaBuVX/hH2+xER/S4zl+5bg6PdKUvzPsrFCqOpW7fi+T1UusUF/upj0
piVsBkUUt5WRiK04VROXyCIJVyT94Lc4/654sn3+KesrfLa9Hcj/XWzeke6Nlm5RlSqlK5YUq860
tzTtJPvp0tDCbvBeftf6xTWTBlJCIHhIIwTQfJVVizDGawkRcY716DIP2BKOQQUQHTqX3LchVxBB
KWhImMl07Hs2YdzQkqzgFy6Lwub61ONvNKGjsLbi+xF5C6zwdszukyxnQok4g4srGsgd/MEzXW2f
+0hEdqDgvO/un5K4xTBG7GKwFhl+T54Ji3f6WFEKnkAhGGW1xH44WDReqQoud3axfMEw3xpLpXr9
qmBbRGPvk91OCyQZsQdxIp7nlL4WQb/CqsNKRcF6Ol2wdKy93xq8DS5wH0qL1lF9LJvXY+/ZBVTs
C4pPjzt0/tATntdR2FRsKDp7kQXjUW6yncCAnWnhVHCwOIrn5bFJ8UhjyTqw/qjN6v6MiDzmFijU
cv/an+qWVqhHryfFD6DWnFE4CwZJQJpZxKxcbrfoQ3nHRT817eguYnZWULqpxJM9xTaXhetrBt0p
9U0J48UUGN1ymrKKOwhQJ6ionza85fbTPCCPjqREhl0SCdtgMV9Dyy+aAIyL3iGa/qKNKoyhByB3
Q8mbzbJ/aCytEzSoDLtOjqPXTf6MIsPnluVbkj3rk8FbcG+PjTMnGPRB/9D86JVJcKcJhxMHKnol
F0+NaQWWZYOhPCU5ws34HQDq92jRuqspxNtoM5eVN0fHGu69egGHUOOgKGlaKstPnyW7v+/dZeBZ
A6B/trt68ILVWz7LQdL90HewChGSzn/+ozI5lPWD0qokf1B4/CO845OiqKsY3S1hL96SAgyJ7H2q
lXPnUa/YBtUi/Y3ES4pJDbv6FkNQ6PQHLHavgLMYgnmZtZZ1G15lDrCBiVshKrsyJlvbU3oqEfq4
yTWvy9NeWkYcOB4YOLNE3AmrelaGViCsZihKDj3ZLXdPWeeT/wRy0xj79xZfLggSLj6v0CPuNMgj
s664XJpdsNpqInDIbDKe+wUy2L/PVxfA8w5YFl8Yl7iwbswCCl/VoUGXdvL9nujGbtzxIxHK+LO3
RgBPbxQhmmyU7Lrr1J/P35XnNdiDkoacrqFBqrp1uw4lq/2g6f9vUPzA8+NMW59AJ2Lpz0u3sDwd
9wgcxcoZgtNWJSzI1TJKGO/E4JGl670b0g3MWnIUpQyD3VWwQbov686crXCzZZEqk/xM5fHwDOC/
xAIdoiD/zR4GjQi3KrZ7YIiCeI4cL7vKEsysznIQ3WqhE8IHreym2jVvl5qeSa/4c/Ya0tOyRmU3
XmGJHbGDHuAEU43g4Of4oAvFgNqBEDU2cMNxlShfriNlTmsR0Of9eVUYiQcg7zp4iDrD2joVWLAZ
4zwTix/reLhuGzXXvoK7X2BS8e86EoqRJwQMTvWWzQkrxFcwWa+P2luy/xFOtSARiewxPeZhnimX
Ftfa6z0YPrrjsiAKB8mBvAG9XHN/jCRNhe/TJ3v2FSNh3g4IURFqwb3u0fppHU6tVAwpSoiCM6CZ
Nw9FJhTGh4HgpZQhY5V5EsB0q3fBly725GDAmDdlDGAwZnn4UJZpgJqz6a21CdE9/Akva/onLDBm
oLLZuStS6DCYrYBBwDmXC441T61x8T3ZvjS3VGPB8F07a+IcfNybDJIuMyxHoyGI1ff0qps09b2M
28kIUFoul0ej9s9EXDrNcDdSerEEAZOGWRhfEVbwid5duvsIlTaUu8hoFkv4PgN2mqjd1gl8avaf
3dOPgvUmQmmj0UoavAEPJXYeLd0WJcJjDiTfEzIpQUVxoHDibIJxRv5OpHV/By8D/ALliwcVPtph
VIXepPoKOIzOBfqWSO9GGwylAGogRYBVYk7gBmFhs8F9URi/lM/3ug/fPz35uj0VIYpHfuB5p2c9
9kQpEv+4axUXwKyR3IgGLe+P9GycRIGBbNdbQJiHb2FFq3VRmApjFZtZJ8KRWhM0Nl0WsZAcH5kn
IMr7cunF7S9S+ZmSD4PT2o4DfHAEPSSIyy7glAOGrWWLuo9nhiky+n11B+ymBtLxH51COiS/VMTN
FZi/JGMNnvfq8C0VL1epELnFNJx57pwMf6Wz8GRC7p8j7azs/qtEWYVug+2mSLtY2+YPzpF3orHN
Pz6iT31jgbHnvMWX9Y89fizdiLz11OhzgkQ4XashIGEn+/rtq/BovwodpUZrP0kJZ+3WwrMlDnFI
zhwGwPrvB97wf+1EGDawC6PXs/T3dkfhqQ/qJrz+rj0kCgT2rqW9Y5reSXOK0s0c7uyPv4uEJCDV
44QCn0FHJ35e9MGP/Ec48+W84TZ110YYlBZRvUxYo+Rfq/g2+YMiujbb8ucCA4qeHS3IFqlWBmX+
QdStzd1XZH6g5zkWxG+ykPAwaQDZ08gnB2uirAqjBjEcjZcyhnFcBckkQD/Zgs9si6zvDfhymqi8
I3/vT/x8d8jNx5pPv/cLa6DfKUhYOqyRBweZHZYnXf2E9MbiLaB7zHTfhMJ2e8/Q+BkNx3ni01qB
XDDKI2D73fdLhg3Do6QwMF7+0/y8H0PBMBtMgHEXI8mib39Og6EnUgcrvmjmSjpg/utZ6hP22aPa
l46pUVc7NLTaTwlo3ukmtJsnTJJM2gCBZ+Vum9h6E0nl7HgtKJC2vdLbAsjlQfeAPpcueDT7n6Jm
q1D0V763YZK1wbcFbi+poLfnuMX3GcmLWFwrGP4YFBEVmzatH659FI5I3myiU3U5fIzN9SQn4l1b
wAmQvbwEnSJSPOAxd9ksUVTcC3XaOX96Q7B8el8Jy9HqmNsvpkBeSYO8Cv3ff9VyEB0XC3duyNJE
c+cC+yeXZ+xxP1xsynH32nW6OEcN/qprXvNvi9LJadhLKhC5rC+a+VlJjVpM+ESmjNDj+pKQ2awQ
qO/iexOiscDcM3IoQaDMeOn2rhwFU8ceeKyI9KP6MDjr4+d4lrICSih8OLOSmt6msVx3a+aDTJ6W
rA2bV4uIEDLJx6sI+PmQjqzwh3vJvuy96fKp32u1HCxY9s7j/I9A132m8ehZ6PjaOGD7pmzC1Xip
WjgCNs6Ma7P0735YhhO9iX9/ekAG6XgD7C9frVdmdqOod8DFRFtURmr0HtvHsycQ0UcUoodiVjzF
BWlDmaiiiWHYnXueVc4+n/wPcCfEaKnnMRl/Berh6djMfE6PzhIHjBVETvrYKwrcwev91US8N6m4
RAA94Kb6e/ITmr8IS05QvVDtH+BmbMS84FLUsbC0NQNFGE7N66flI6UxENxrAx7p/bOYnys1qkn/
TLWeuZOUez06RXnwyQcPHafeIpdoSCP1UVrmPcwDgrSd4u2jfhd2BxAYn8ZVbAAL4ehIs5IdpXU8
g7wvyf0U+FGOTD7ZcnnX1w0aRDksTgec7x9RO8Qc7mo0Kuh7KLYPY65b310yRiZWhRrb0J/KGtRU
eNCkaw6eh+PSXMQ6ZMW43otMBLQVAtp3LCIUXCVYYsAmqCm1s520BLHpH4z1aTxfhbbgoufCfseH
jim0+OBixQM9Ofo0GY/Vc8wJycpZAB5px8heYzlL9IatQanz9CamJDRetKRDz8Mi/kYuevaUMuDJ
ouJW12sndQC7zftEmjDJQH4falemKycHfiltQLh5TFTs4V6yvM9HuzScJcF0ALr5cyiKmGLW2YJG
nSZ2JH1E2FQJF4Fo+MGMjG/jeJnXtpMrNJSxyB4j7ByuKp5b9WEH8YwdOU8MrEKwyI/kNw6aBLQ8
cw2Hth22KT46/ZpHXTEbR81QYmiYh/10sdcnM+shSj3XSW+iYIiHKG2tB1lh4ZykIO/dxWfGrYmJ
h8wdFvIalsjovUgMQt16j8y77Dm/Ojh+gP1+nsUZpY6fg0hkqALINnYa+Qej50yZMTnMnGBTu2gB
9CidAjuS0EkhCnxoWip+LryLTh7Qh8Grlz3a1l/u7kfHrPQWD5HLRo7Dk0rYDaN3yVzZ+P623VgB
j7tFPGQAipDfDGd/hFRdkVCfJFoCL/1jRgyhK6xcE7ba0RzvBxSXKh1Qoo2JCN3BVItBefEBf/6+
fo9lF14NRKjlVRCwZU2xHeNa+YrJkTr/YQST2GecchopuxZU1FQRDR6ZGk1FAoi7OsyMKWl+zS25
jg0whpAkogRN3cEMOsQPYLmJ+M7SQSHpjmJ0LCEiUkPLx8FcmIW42pFeO/Ns8R7TEYM9ISih4t1A
SOVoHlFtjoaeP8A02Jb0sLjP/6xBIp3A962hT1IQ/VB2XtNGA4sYj18H6y3TLLKYTR4q7GKq+APK
uSNB9ZM225m8bvmbKjnTL7jNt3SLXGkr57rVw59dWZSL4iTzKjvvftnNY9NuQgb4VGWtOcNnGebN
hOPvKM95QsgsjI1Zlb6QOnRbuLk0YkS396c/jlbmHAx6o64OjzYLwKYfdq7z1EGzDlQF5C0hLOJk
jT/lteQOwkfbnjSV0qeFmttqkcZaWdo91DlFNA1kYNzw0GMAsPv2pdS+vfhY5mGFFKjIVvv/8vy8
YhYNtfpn8yPDZczRfJFjDIjMEkd5DRgt0lXmrkB3cfBb2PN+fMeYLYrRuXiBpCR4sfogO56LoD//
2tlwEH8y3i5gZgiJZ57l3zoUntcf1GtPnlnjeyfZOyky3yefiVkJuU9YqtHcRHSbigssepKPaDNS
okKgGoHGmJm2gPcYxu9H+mePSZHsocdExTKBmEldt8vDyYHU62jzJirpDtnxsd6w/Ys8O0T0CIEi
FeqkaYFuFzJuRJr6YN8al9d1qOizRw+PlBXEbOeL2pW+tXwz80Ke/He71YPsZeyF6ZIPXjUo8MhT
lwHuN0/5INyxxEQ6/iTb89TBJYS8EEb3PZauUxgo+H2PLayHCuEs0EFFDeE+V+QnPVznwc/EzpaN
rjPxO2RdEwtMrPCy7cc8E2hxs771DRv4EiRa0sSKtCnl2eFaaK5v/AG9Q6Lgt5YVYPxL6Qcobmkq
1FVC/L04auyxdwt92h5qJQGQflhTEZhZgyxch2JD10djDNz43rJjl9VUcwFHgTDeGGgjjAsjFaoA
kQ6EFixV6M57hg+36a39GE7xmNlvXVuI2kp5pFPu7PYTfQhIyM3DNLRyvY8SvvpgCXXpq7+vsbFr
aKxFgMUsQcOFScGgdqIRUN/FDpzUpC50DbDbG12tZm0fYXdbPFxx9zLqAeh6HuzX3HywozKFqfWV
1TKHzdVTkeIsA6nQ7EcDIjNme8Jdg8Jd8FhXeGse8v+ly7xbUe/wH7RHl7NiGJXoVCvYZ2k7XEfy
ZgKMUgj9mvWLwg50CBctqdq5oirMkFzoIpwwwoeJFe0afB1JRQjJWvERe3IQZCXIrAsc07rEwgOs
oax/XnJN1/c+ksELqPw3rBVhKXmYpgjM24BK8qHwKLMHR+5b9arQ9BSKkswXOUta1AP6y8ZEaoAQ
g7D6p9yaupN3LErQR2+BHmyqOXx5OjhpRix2KRG9hZa4eNN/UHfuCvaOhZvq9l9bigxjatUFBPUO
h+ssQNMi1ozEq1F5ArUYhUGX/WmL1Vj/UTgRoWQARzr+IHFu8cHObOON9LK0hyX4vLkAQdh/6UX0
MGe77mtXIieN4FU2wRxwBrxb8fmFIhBM+k7SvTZAJFhLdigDD5MQr3sEZcYewVOjbX+3c8cBD/4m
A+VA7walKX9LMFEENOLo2eAV88GvKVvxM8ClM3pu+QXJTZEOUC4iXYepOkwQyvLZTUqDppxpkRdE
VJv14dCQ+xGtuh0Mtg2Tr8xImf62ElTIu6/q5iPtxQYzObhROf2RHlI4diGjaXi3tdHT0s+Ow3ge
AFweRkWe6FS97pRE3T+GPKUyt7GpmiL4VC69HTEgcVof5JCXF9qbK3K5Ihan3x+a2dYCVLWc0zdS
QJ3gfAkJHWPWdjZUfupSGfD02xULa7cZSUyZlQCGarNmkw2HX6CJCgSNNH7jzcZBGLgQWqxZPX8m
dMlKeulYHmnK012CUAGxfOasPWrnU4yQ+CodHSDkg+TrG+ruWJU0ie14ataWLG6JB9wqPc8oCEFq
nXoS0dkYbLb4mJ/KTX6coWA3KA/p5eNu2wWo01KvbiElAJCONo96+WtLwqz5pIsi2O1rMcs8125w
56NhxEtYBGkNYyqS8wAcXvTFMrnwYUm0zp/LcN7uEBSVmvJfedC30UV81U/e0JFEzTF/zNFvmSTf
d1SYkZ5JrZ240jB0EMwBpVUvV5VOOOOExuxq/OIGZ8W5PBlsaLxLYylIbk/SV5KvnUiYlGvu3Iq4
ZlZiln7QAgX8OlYCHqODGXqgzh3f4hJ0yS5m073PRFOdilg7Gh4sa74WLX2b2U5/tOaVciphwGlb
Cp15EuboLvy4muBjyBg/PmXq/DEi05j/1p4fy5/wmanA1CbPPua0KeIPprnrsWi5/x9dDyy7Oh0B
YzVduQEwInWLsD5tvfLxAb+jUiX1I1lySQ4BjFQd3y3Dm3C+lKsAOYtKfNBfLfdJrPaNasrmBlnZ
z0U3xgNiw1RTaMLWi3UnsZy7rdckiVIwVMYBPDPvNo8eMx1RVajlcj2tmHdf1LloP016e6z1fp11
ooojqbYDd5sNmVPRux+sIn8USSg9bEFmYzLpqupqRyyMCPAEav7tCa7aj3TH2vRJy+ONRJSVSOG4
gW4l/D/AINGcwdOywIvW2J4Z4dQ4CIQQwsHibcqTE+34jdagBfVXMYb1aWWzBUd6qlb4wDABx2w2
qAYCswMPCoU9YLWmNUb6/oYSWtWTxrJP67CVMz3Gz8w2MUIDj5wEpIpjPvwCUAIA+qa9BI1pL4Dh
4PPiESpme0ZzjSKFKJsenqYhHXbP+46AB/DqS68sE6reprUghLf1aW8xgxfJnuoEGYPjdqnJS9S6
TJ9rvYaif8fDDrAs1qVdc5YvSL4MGSig+SmZ0XpCoyK5ZFMe2pEHgk62Fihmq+ZPyE2hBE1LG2wd
Y6C1UjiUoCv0RMbSGzs6/vHwwjXVh/CGwNPIXuHBxhps2gSOyWk3em2n/9BE7XHLN0Wu1OANzpKF
2WPtN2UFS96o1z8PbLF2sOKzKJ0wGE8JjUf4nkJ+ELsR7mJbs4DGgI+9aQ769nkleczMuJMJZiJu
HjfNSSIo7qWTDPpVEPi5JZthWUMMl3iQFT1xrxgak11odxcjoIG7uEKc7PhOR/gVWyN6flJUT4C4
5dTD4D0Q3mT7CmCjvR2Hz5MjEXGLQLON4hE/imPS0oTHQ9jmHHYprS1fa6jLWe/3qEwvO2rEj3Ma
HvrULZ6VCnrXtGxx0ILHMYFeyYecbXU1hvoJVvBTO12hefwrYmhItTz1oMpAGhjUb4x0ajghzrHe
YIWFhMVO/mnzjrLQ8SD9P6qq9EAYKZaA6b9KBr5+o0bPWi0cfcIrmGe5DAEAzBq0S0qC46AY6MLJ
uuOcvlecmflQtD6Fg1Rxw3ZAZSDj2eWTqHcn9OFPiu8B1AgLvqVMRdFZ+T1piC2rMYz9Vmr4P1Bv
MtpJqQHxmTV/dm/UiF5BIaPHNyQ8KHAHijScWZDf21/t0uGqEvgnp7YMJJFlFxO+eix8+q61v8F3
F81SljGZkbiarp9Po2Y533wNeJexpfRux+8fWoZSUxnmTAR3yxq0HzVQL4MHcG9Y0E+Qiw8Jog//
OeVtzSIvD1bCzrhFZD8R479UUYAvsUFLaU1Ws9Ii/VcjpZxqEGAvr8YVkdss9bHwuQPhfbJHb3FY
KqWG4088jmrfYGlZMlRKo2mbvd4rI0L6qkfjgrsgje5gkv7sNnc5AoeAkeThgIIhCuYBHoVXU+Vi
hXF/1dL7ki/BEsie1crYcbqOb0wP6FHDpKJhIJqIG5POXz96RzWtKyj2nVoeMUzn60wyMIt9/ayT
MfuYuZ44chDhcxBSfLfDB9/m6J2qF853cW5iQLt5p8MvfXyg8FxfivUa4Dq+bjjQMOk2z2z455zg
UaOacS6WLdf0grXiURweT+BUhnnrkPK8zZ7wt3waK+TyI0JGVkbOgcsBC1XJ2AVLwyj+4tr2M3iO
9fFM9M3FD4PncR6Fd1DsEa+SoH2fQCyuSFF+Ts6oK2yziMCqIQP403DjxA+3oEctXl+ABdig6c5a
DYcIlDJ3mnlB2VI72/Tob1eGIjikkfNcOEsr/VfB2R0CkOkQv45WH9BoqznnEsWZ3DS1quVTSP7P
SfuRD4/dInKlysJMFX2XaqsM+SQNjmm2idtL6ZH5L23ho2GC88j60Hkh8gzG+lUW6+4REDqhzyOo
oMGk5qdJq4c4cXRL8QLLpV+mE0g45mIwWnNvPWKJm50vx+75ZkVPk/8YJev1GcLt4ykPs7fG8Pxh
t8YJx3ICxq0X0RbHyHTNa21DtUayDz22i45Iak1+w+pIcPsZPZsT2fH8Ek6WWKZiZ5sW7vJTA/lI
eD1KnVv8i67Uf+ypI2/Zo1WESMIelmwoHJ8qfEmkzUNNYRpGZwXob10xayMnoXGOfjCg/JQswkEc
CryG+DJKdEOnU+jAgqZVX7nGPCVW2Yud91EQMlfjSxW+g8TKRpwBMjG9vuTJkwWzoXRWN/ZcP1T4
J9scSO/iAlWDA88VaDfOQYF6lpr2JK92ZSXZJeDjmlfBMS0HvhWZKF5KETGfk2w2LZ92PXbR1dZw
EznQvMhd0Gho7s7bJ3IrokGCuNvl8qdr1zmEmFWOWh/U2z8SFcr75l35eVZEiirjQ3fC67rHfVp3
3hXAcZpYQXA+rlVpH2QtlFZZJTFeUukd8HKSOKyFqHcNK8yCLwsqOnODELfLWCbEmYSWk5a6Mcs5
D1w1omYAjCDkbs4fc7Psk8pJDrHdY35X0WHBfqRMRQP2wvSJRdODk6nTFqsWImj+rDIIPiw5wnGI
YKlsmE4J2W5m0XKeXe/0BkKUbYEQ7hYdX+VLHx/C+GgEYeooihDvhmqFUHaR1D+WRkD5/tFhol1G
4KI+EBwZQRpAsow5Y/jLwebjcvjIe+Ya008aq+FSEKG/g+9saThhyHYsR6IQmDtUu+hYefjfcqQF
AVkKpRpxvIuK0kON87OW+8ViuoKWsRTtgNO3H20p2R2UWHCCZDZSdd6qFExEpRqs1rpsRPTe2HnM
Qrzd4Ro30P8aO2SgnMWFMxcMnuxAem+Qg64MiKHXe3xfKarA87BIGoOqaNQlB4+iPonZORND58LI
Q6Bt8zTaTxaypOLkfajn5AhEWHAkdnpyJ5lRFagPOaJ5UUIdTxY9CJ4H80V+7T0E4n2fEjHNGoRW
gJnZ2skqPErBeGhQU9S6tSuwWtsKyUb79s0ScDfsdME+dqY9EExQsiwxVSjPvgupA8uYTLuciH7n
oA8P4Hw4Ygzo5ZJj6GlvvxsMTUFup70zTSvbRUUIGyxctPRhRefoB0tfpuhSjLRdftoxT3Sdq+ci
dvIXhXWXXfTMTbLWh84PO/LUdjZbLLizNlsobJLpA7Zq2/pBZDa8Us/3ggJFjCBpqHc2ynDgIzT+
LzXqDaNDYyP2TCW3QVrNJRqdzzXTZ1BNfTWXR3eslrl4ZjHgQWc4egwZVXGPkyDJuDnS6Ncts28e
Y9QDJRKnWBRl6AWgt8ySqb1Bk4cLv9Z512NAmKDEEsJHJ3kMGyh2wkzYeQliBzgy5+N6trrVvmCN
6eeLdYAXb30BcBQ7HZJrhkipxZ13RzrBkDUoSiX5ct+gty16CvmB5aX40Ksd9Al7bSU8vi7OEKh2
CGEhUm0TMpdnQwZ+E+O1ePGF4zPS11xuWXHG/UNbqZeEfQRu0ZCZk9ngmR/5U7WRXBhkx/L6vyON
erjzXfqowE2Adm2EhAGCz0Uvd+aeIPt3h1V7EHzxwzATiyfIExBSBbRvF0iHW4fZjWj2gld6WMSg
npuYI7jQmXMeT7QC4KitzpGBtDNJtMDiDW87JW3Wj9VobG+Quiw7dDrg/NHC6juQ0/Rpc7iR9RBn
OvuwpDyXZ6tIIYgyI0ewFxdfwJT4IaTH8PzaBcnrNIZJon0npu7E0UNiZte7NyfYRU/XTiKWCSeK
XwvLktIdHgBtnv2LB7IswBxrPImo0j+/bd9T4BeXr7aaUTB+/C/qNH+NLynFUquyVAI+L9vfIzdJ
MUdIjJUCddcuuSftM4U+BDDpkpt7JSeeQjkdVg8km8UwfkIWHsH9gd72m+A+lY3YbdSki/3KaQ+y
grU4pWw0b2w8+tO78Mj6eJFQLEz9kCV5xznoMebNvQzlHyv8r0/eH+jhx6JHrlm6ta8R+ui8TQfO
xINKQ1dv/LazQ6QaG9lB8qvW3dlBiqc5e01wlxjWGn5UauzKvmkUbUPyvo5rYQoAxfCK6GVnbZSl
IuZFH5YdDsmLTcE8kOEZEGo9/fq7WyBMciwUaREC4IXTQTx2kTTi/PahuklkeANZ7BBWF+GYb2yb
mHWXSr1Eg1A7bp3TzMWJPHpacXao+vNbyqNl65tc71xFnkZDX38siRvwZZsC7/X/hLqnYg56IWC4
9Qv4kUlEvWjpZwKhQWzKn6lGCciSgilF+SoTRD9/5GgyoueU0meQYroD+7Ai1RJNS398ZIZt7CaF
FxMahT2DTfOgfeHvFb0yd6JOcSW6CN24DYLdouIHFnGwrFZJNbRMkWISMPj/zig6KN3mlFrWuwA/
ixgmAVmgSeakyLIqPP6UL1GVfcuSqAG4Vl8MBLu/SpqutzExk67+N5ZYzHqyT7wkrkiQy5a0jYQv
tCrpn19zncEXztUNi5b38KhJfKVx/o27bk6kj50ZqrEkHQ8WZ2KOx5AfuSm2/dnbbFjustNlgPwG
kT21vbpKbr/J2MYcnqHpulFUN4/0yAfJgZ99wtqZKkQYEiTNBHox66XQ6GtWObOIfodn4cuZjGhC
QQ4nbA3qyirnxUxCWVdA1E5wRBaier92bLtgkhjGfvRtgTewkgDOeOlBvQwCT+h5csJkIl85567W
UKNMzrvguA8Z74MUtZ99eOnzswF9vXDgtkUi1RzjVmrI1o22vmKTYttN/XWRq2/SVa/UCrzuJagH
ubK2BzBWHyvykAp52aquaYPNBpy8iC3qIiIAxDDMrqu9rCzh7mMcpI8mVqhSkIwLkewuIgbQJu9y
VYpgFL/Bv1a8MrsDTvuZayz/VJGz901npmfZ9E0Tmmk51yvEe0Zj0iwKw3lUFjPgQTBXHFuV38qt
qU9wuUSfX4Jk1Y0Yfsh26yXF+Kp6Hem9fAvbzU4vphoYqpd2QegGFTcrk1SEagG5YNfiGc9lVV9n
BV6mPzk6jb3gb3JqCFjFyPjroTUCRb6NC7CUxsodM/r5Ta7bmGhWCy9/I7ZF671dR80NiNOOkBtJ
x9r3ScMObHZaxcRaDJmdTu0PVoRZl/aPIFwvv/SLqBM/4XiZaInpqale0wkhG99M59UULLmxP+BF
dFGO45PSg8bRDLTGZAVNXzpwVUvu0jKsk2ftzRg3FBc1l9dnaaFUPGkQbepCj+ifviMAtDF/gORy
DQFw4KbWbtKNtbZwflII1X2USdtOM9ouqIFV3Xed/qUpDUPOOaAzK19s7Ok8rveqGmKn2vbpJ0+H
mwgjJVebj0RfOgjDKCpm6anByPcuUacPbEVBtZp9rqn2yXdy5dxmrAb4w39E6nhU89wqc9vd21Fi
pd0g7DZXVRyDI+hvycLDyS6tTpi0w7j+Whhh8A6fHsxQB6YTJYexVdLWN3AHT+ugj5YKYa9S9254
Ys4SkIKltvlegNoqJCEL7y6HQux4PF4oc+FVfuz93l5lXcwgl8rSnl5e2Hvgo1RFiVCnstQ9M70r
vD1CbylxTwrNLdBrqbfVP4jnKPkxkUkv7c0YPkyU+r0epdldf8L/hw4Rv+g+MO5C3x6rWon4Zu3W
JLyFiAPsFX/7o/O1aKRKmhIPY+imybUG4wUhyPiEBq7kTDgYfh9WErZ4N8xSi2K99MjEowLrTmYm
FGoxKSZexb87v49VLX67Zzz0GqUWimiZ5xjo5hs5PeQ6nOJOEtJSevVowPPo735xZr/ETW7Myi62
8fbR5v/g4D8w2DBEzoGeZyx7EvaGFyYxCfSmy1WTXEcXN5DpUWW7SK52/iXylL4YcJ4iENMNpgzb
G0XV9QfZ2OevFmSpEmwlGLHjuXq8ZHfTFBhSYOeHCet7KNcqmQKl1nZC4m/GUTLEpRFet7fzMOBx
UIpnTHNEI+CgIMpBgTp1lkMh49pUaVhp7tW7527nkIXlyDtdtohSxrFNcI8AcDt865uHEzer9+mo
FCts5RcChRMkqGh1LitM1VES8rqLft31bVNMuPaSYJVbBG82+RBT3t3Vl1omcUhczqqovFjBHNQp
A1zuKz4hfI3F2iUlA9mz7cwz7h+xZOCwcaQQWPGN+vdm/0v1BxyKhkO4gUwYEwj2i/f8oWDRLFOR
tSSDe3xHZ2bsaoPCCPMz1jwVDjiRRxZ8mO7LdYU7zi4RcyTW8kfEpk+ItpbHoVLD8ky/Ut7UW497
EQZw96lWZu/8PyUz95HaJHwjwdQKstaZQOew/p4HCOgBvuSCJ5KKp6HsP7SvuJBt6RZ4gkHvE/Kl
jFfyiK2Xn+PelbEXZqkfYyOcI/fmQqiRR5AUtoaozWWcYYL05CJspniBg1Z2lyIotBQMC2WCKhC+
3MYHJEhxOyvtKDpHD4WzDeoYdpJD3mtfgDlFgbjcpjcpMUbEKJMBsyWrKXj4M5a/d5hwMfqMxI8U
tejn5WgPumorVzLwprsojvWx/iK9nQHe7kehkIQtJip4NWW5yHs2lNi/ORlR1dIjTBeb3coFYRnb
YaBoGTp3zxICNaAdtmbUPLeXul0KaG4RTDnHMpxcV0szJIAE6jtV6VLuVvhkjC7SfAZfDc2JFq00
ZfrXJI7gnUlHg6xK7R6V870U7nENJTQfgwJr01Q92TOmGy4rgCCt2gWoPYA90AzzdCcQWVf3+gec
Dd7aNTjpz0CEh78LyQhUUHzoklZndGvdgQLXJVsik5VReO7K5Qiyr+Em72d/uNGKoJbdBSvjcRUD
9JFFlXMPZrYUVR00iwudcibegGUomWBQtIBKDvEWDC4ztEbXcMVBALNzbG991leck1fJKjWg7Hc8
JXzjwfFGdGwzjU6K7ItJdG+cebQ2Gr/+IfTWQXcrDhYycOFWj+FeyQVzxaXJ5An393FZN+sJV+g9
Elb9r1LhOQhcj6cc4giD4Jb71nd3OAGzzHEpYM+gUeGz3MZjfKKmES9G4blIZGkbB+O29qrn+/yO
onD4VSoX1zpJ740o9/F68YqCgVQiivBtLOy2I4pJOOUOSWLdZ+7gT1rPiIcXGt9XbP/NbYLvsmfw
w9K4ucX/QwoYoo3xgZtRN6pdUe2mf+Bzi0zAzTdfvcxcdstYuBLU0olVM6VfgdV1BppTDFpqr3Z7
onLlaKpKtjyJ496BKxPHwB6Mkk5lfXhFtJJ3WIu36be1TQZywOfJUm/hBbEWEQBhIwc+CXpPboja
zy8TTKiWmEwxABIP+v8rKAaVN/Yxj8Ja+xb8rVFjEAebp2NdFh4fr2LHEsL0X1pSH3qoXRa059iM
AIfO4RSg1Pa4ejijzCO+4Zq6E4MsIwzNhUaP1L9TmVglNJ6jyGXiwbbO9pTJmOQ1Q0jVqQ4GY/S9
QfqB7O2rdk1aEw35CglK+FRGpqY/6ClSlcZcExjDwVh98Klreg9LYZdG56AoPgDEm+1KLflCfky1
C/SH2OIrkcLGiZdPvg27in8Yq+Dl7DCG6/+NxREwOIcNl9TTx7wZZbFJ3VxhS2ZAgw6wvhb8R1XB
a+ePdAwukzpjFgZexHDQsO9+Zt2HS4TJ7Laa2T5GyxdMVDBSbhjPR/Ith7ufN3ksY/BEC4qiMqq1
ElBsrAsQfVaOY3XvrJneRvNSVMUrm0s9ZymOtspqgxjOdbNeekTyRBqattUFJp2Cr0b5OrcG94aT
8en1s2GOuL/IAJsoeB9wr0QwAzX21yyweuysghLljNlbg8Yq9wCXFjvOQRFYuJadpAPj+P1/oxwp
ANE7iuwJULYYGshsCR/Rqg4/w4vpcVQE7tCdYA6+Y+1h2y9RDcWiZhZQMgy8AOEy9vfwVfSo2dH8
WjKdAVSyEzSt1aUO6Hd2VJJYtws0z+guEZ8xwYjzVjL76Nz342XVlgtI4i3N3hrVrHlh2wOsZGZJ
yxeqbRRNL+pgYvswq+Q6RciBRqNs2EKrmNJdA7CgcpeTr4qfMWncQr5JvThrV3aiGCLyaH4brRk9
bauN4PQfmCC8pWW5hCrYAiHbv6bP7NXm6jRRyViLpEk2l9vHVKJtZSHIYXg3BNVnLv0FUPmXWl0Z
YkBD66uNe6n9ql8MN+dtA9OdeuNKun75bAdDf+lMfSfyd1pQWuPMvESceuADOuiDl9mR2Z6E1RTw
QcqoKqDZU+ytjnSKVRBXa4TChx4kaZERQAHwtvrWeN73jIoHeSQ6eTi2XAhutkE3ZbADefACpkva
C7z57m73nfmX/flu031P7HN+wz8+E/8zZTJMyk1ouPnZRAkw+BGCBIgx3XJvoaTZvm2skYFvhA54
t/CniRqxPzTc11XU/VMi+hVrrJG+1aiIvyRWuHeou4u6dnGz+/TyiTWk+KnIssS3ktw2z6qE51Eg
u4G2ZqdBVIsvimcIdqzWPCzM1H8W1paRcCdoxcPWU1GS/45sLIyBEemp+ATPiYd6cOyyA2uevoBF
5vY9MjnVI7m37N3ZJyogm2UrN8nOrzM1v9uihvkGk1yFIizKY/qDiDylXLD7slCSgEQ9UkWHrXqh
Mto/Nee6oOOMo912ffq0zf5oLmzK+uAxWzarfenROtRmFpHe6RxpH4ZPM8PSY7dFWMVVcEQHRsID
dqpmQp5a1qBwHGtKkGXeaCLnc2dD+db8h5z7y4ogFSp0deIWj5xUzH6VGtll2u7Zpl2h00+NL7VP
+2ZN4F78lcyj5zJcdAt+O+4txi+7Gxmp5ippC5OeLao50RZdWadGRkF1hX86Hhr7MI8mczwsBnmx
0QLElfWeQaAJhIDhNv6cRCMkNmrzp92eB1biDx0g9/tMew4IldESgKr6jSeEfh38krk6N6E9zVeL
tVS5PTx1tjTQVad/aJVO1aj0StROYCB+76Ag+LUMAoc6CYVjT/gNqAjk3UqkzXD914rrfbFKmvJ+
KeY/Mr5kcvAN36GMuN2zVDC2jUzNCZrgWHJDnMDxyQNlvhM8TEBRheCbI0aBXSQ7pefHv2xvbCRd
7zs0DDwMVn4EqvZp8z53FLFyFLi61nC57Fs9g1zsrAGGHzsVyGTzxY1FtxWN7OPzOfyphGfktfTn
R7gChpGhDH5i587LVzXwkZOSwxtULUonCDCf48Zsxon/arcmpUEADkXyG0uwnkUKfO669YEUCQcq
Gdhz79wMpBzQIzE4SVAULfESVcIzfPRkhQbvHuzq5R8hxBYDe0Dvt0ofC+YHQZcbDsZcoMp/lkbj
I98hbDPNJVRROUTxUExwwcYdBMAG6TKzKPZIdthZBBFcc01QxmhOjzTFDXmQM5m3qMq8JlhgjJSR
lAO1EzWbfzHzqMxFJ2CNhNo2JLDREoRkowRhxC80qnOnsT3h32WDDWfFMepKPHrH3tE3bSOHR44R
a+0P867G5taZs5ocbzDZKLT18/gtbk51LB3V6WRcS6/wr72BRv+2drYGenpFkpcNckbMK2KsESCF
g+xhwldQPB7d1AbRbX3m7DzsCcQAzWPgD0fN4qK0MRP7fGOGnRvmnVQArH0UIUKw5wYU5uONSrRw
RvStLS2j8etRBs2g4MMJlwIKHGTTAkWXfQIjXrXs8ZgW5QwKTq2173rYg84F33QaNgvxQL6yjp68
WmS31cTXaoJ1Uov0tPxlDDviWDDm1QJXMb14CDJDeoYlGY2hd1bO9eh1zgPIhwiVe30bsBCExPNr
Y41i84zQdKRXlPwpTxOAXOSjssSPU96hwj6Jk8e9lXOtsfCyV/aqRXhYQDSVr8GmyrF3xHyPpc1W
smR0ZTHChRT1PgyxTM0TvVnyTfXIkesgEbT5Y7ItXAq5CBpYZ85Jo/wvExUiMSG+vgYyw4qY8hCI
o19WkKt6hHor55vu7ExwRnmtwyohf833x0At/X0ok1EkCXXTxBIdGak6TGoJ3PLRF/Qq0bMFRTjK
Woqk5APoxVgQBA8cP0FFUT7rSCmh05mLxEzGtZXhxuoN+0YWi1dB+EyZtBVzUe3O0Nt1gRIpgdz5
IneWx25KnmevzE7VgWCK0LZ01HC19ZjOXpHeY+pI5AMEwTNOq0GMb4mHc8FHqhFXqshPn+DwML03
xX5L8OoXaF5OSWw4FUMrsCnNjBwbCCNqhS6Y0t/REc14LXrH78dl8vc5CVdJhnkYdVv46LYMR3PR
9b/fDXpjeRULMXteCDRMzntaAw6dJICacuvYQBXUfn0EMBxVW9SPgo7NXHAUOLE7VrIyN5lnm6f1
rzN5D+Q/i56gc6dnrhdIhZq08D+RsW5aJGcX6Rb8br6CcKrLk/Of1vC1XtA1FzZDFzPy1Wwm1UjK
O2bFYlkbc2SvS1qZVW20E6+58gDnGvl5lgoAyFkANP0SaUt8ztum5vPLAa+qvhPFSoGQHvov1ili
VM/W24ZqHs1YnlN8Ps296lr1CivKhhOwogvWzZ4ciqcPwgnrlKQKjNeb7WMeJbV3frkvzIDWSiuu
Fx3pYDHZt/BzMyPjkyskV9TBVhPDjLfWAQbPrEpLOb3vJlVFn9WD4FeyyRpwtQUD1p+Ftl7G78l5
TXYddhKLjUoNRjpNtHIQS/dtWusFn9MQtnMZLBeZaDHYESjEnENaqkxpBKrPSXx8XdyJhJCHoCfv
TxhfdBZaYR9YQx99iWyIBqJLC3K0LqBgSGVX584GVd5DHHwh27ZkbFguYJASdp7C41LOKFapWBnD
qjXorN7p2co11niJoTrIc6JGwXuAb3PJps2v4atm+xZp56J6NOlLfVSOncoy48bzQMNE5Eo4+bsI
PoS1IR+qlTuHJdO9FMh8NC3F1Ka0deZInxsWyOmf3CL4IiraU/uEJK7yTASjjEVPsZfNZiX60XiK
nec7rj9KcIs5xQQJ0CL6SMYMp91T1OzKGRePVADLQmW60BRo/Zkf7zdeB/9qKqKyEqrNtspXO2PZ
xJUJFBasn1mio5f0r6droBCo6JHURTlUXVppK5tkRyT1GZbhKFUqQE1XDshrVIXEOrP/Pd+K452m
0DMmdF6oLJ4J7GI0LiquOgJNMyPWucGj3CjJQkyUX4aGRIx77t31VxMRzOYD0llLpuERzFjjqWPB
kulXzytRpgtoD6INgCgfq9U4xB1mVQ8HqDmsbnJNqch3792cJwmNNk2pVs4cDR7n5JHO8GqmsYeH
pJvpaZD56fZ/jCyCnUllBAfKzJSNVscTJnTIA2WOfMSiJlDX0BojLYVvSZelOokMJBXPgBP4ct4f
GjvoPITZbUQFlsg9/n+DqDKkMUo06KoTSvblzxxAQB5JIdh7sW9EKiuMVaHrA2t4EULquT+zjwTu
JHC+uF4WY+ciLVNMDH3cbs7t3lEfO9TE6cl1TnTZfNeus/qjqRC3EPRBVoMiEsRH4pJh+S/q2bn3
L/wgQ/OOBkL5LjutuG2lFFlX3yoeYvoin2gaYugYSWuh0BKpIzvzR8A2F/WwyCAaXj/mBQTUpV3L
nXiidt86B4hkIJymqs10OywKCZlqRKAQM+Gf+GWAqF92GudEnKyFvudohdPe2KbYZr2TFPHvy+9A
r1lAfG6H8M9M2ZYneW5pJXSz5asJbaRX3kMi/bTxzU9H6ZcLOQkg/obXsYaH4cQi8AHkCwi51v+X
iWk157EeE3rwEJwuejrzBfBRpQoZgrkspeTXbRcpb8pVaGX3p/pXs76yHk1spvpgfXdNaeYGjEsM
8ZYTTp21E/6SsMHX3bfg+ARfgWpk1EL/u4UizDTTvmgbJUN/3bB9/7R+eRViSK95vBP3LzWSx8np
A+A4rKC6EqXxjCr7EVgGtpis7rXrCjIFSlv2FoKhjSeUQIH4+aFlpsVBajItj363pHnEKwjyihs3
59zmvXDq1ucUVP6ka4w/XgXU8/zTNc0MfrWEboC7KeZq42QK+PSxrQmlbmdzxspKSKSUGkURnWJa
y4djKEWC/kQxRtUPPlY10/gLElx4O2qLEzKXyccs3XzlGrdWmf1VWjPwsSxYbaDf0sl4Y6tCpUJ5
2/A880CO2lQR3ldc27Q9Jj6cIQATVdSi835mHIvWwKlVLhHejHzSESECi3Tv9ED7/qRlxajLqIT8
ll5jsm6NvVYjKxemFV0oGQzqovIPpXgCaVxjgQVrlRdMwrEurQA3E5KR3H35di9dk6j6dTla8e9Z
FDcir2EuDBAKznYxXeayMTWdTVhWFIRuzjpY59elnXlH/7xvp1QOUMZKN3LJYtNYpj6z4K2EnHVu
g+rzuMnL8eLIpVllNkUwH6E0t+311WueJSCavz2mLe9SNE6bRIixxRTwrec929suye5YqekGe1YM
9HyVjPkingjW3xgOARaD+UGsVal43nieKczHtMJO9uE0NNPlPT8Z3O09Cmiaew7F21CmUEUmBnRl
NRpeXlzldBazEV+NSaVxMWHSd0VEHa0LQx69EqTnM4LVBkbW12O01uxVttYTWkI7gSiQK8IPvVQd
osNLmAMS0yTxb33IVaMg74aPZd7eRTlyQ9LP2lIjpxclDhC6UJaNjcA4NVgH9BQDcm4wrG5MSe9G
vkjNoS/mDn+VHOHp1n57VH6SU0Zg1MbD/m4ne4c0nLkAwlQ92MNx1NIAIBGGDxquggSQo8LdlnA9
W6VGNGkqrnKnQJKJwobcsSpNgNB9tTPHQ8yLaWwN5fu4vf/ais3yVoogGKq01fobZYHzGG9Yf2NP
prK4dL2qXa1goNnlbroCXBp0WYdcONQOOK6bmiVE0xFo0dvJgfCQIgKuLuaOAdUnzOTxhkfjaix+
qdycH4sCRkDXUj60YEWvJBrS20RiXcFTWhR6YuV1vpTkF8lEF679UR7GaE/iyHzHm3knGEeMpTD5
R+Lluy0/iYB0EAZKcbbAPBs4oRftAsd112LRn+mKQr3jKg8+MkrPjEhO6+cytsf847LElpOgcdVj
0+C9MWxNrlD4et3ZkKkRG1X8z5rp+Ii6FqQXHTYfyi9HUwU6CIhblJiSf7WjBQFwBFb+YvkQZ/Zw
InNeFTC3Jm5X1IiUGdsC2Q3fzRJ2Tud2F63HQJyrTs1gvXln/CYM3P7tFUFjB9jFqI++gsw3P2lX
PqighhEXgaZro8D739U9YaZtmo6hLAMWfrpiUBft30H7UZ/GWWDeOYVYNljec4EvHlshTqRNZF5p
35+lpYjpY/qXZXMhm+OzLG97nLxYGfm2WngBFxk3Vt5tSbLKilGPXgPMwdVwfCjfGCXj1vHganAB
pk1XzrB64+Hehpnhy2zUXze9GDvwtRiyVmsPjSSC5tt93FqemT+DV+xPTeLzgmxts/83GiwG4m+c
FdAMVsrCnEBFKkSSBrSBV4fDPzp4QLduNVeSiy0LdJoPzN8Jk+jJLZMLJuXkG993oeaEV8FYnmYH
uE69Bq3KhrdhfGM9ujgO3ji3udg1Fmtbqfu1qVP6hEr1L8/ON99RCsawOTuuzV48DLN9aYPT3Fvk
Lbhn4e4DKD/iDiPNJ6X5AdaEgi/TJMPYJTg2+rRVK1YO3xmIARe9Jef/QkSd1qTnsV8loqnT11kC
9XTVYvwXqMwkJmhw5ZsgskgmSo7fYYql1m13Vl7OZ72TKQ0ilRICpiu4y/JkQ2L+bBQ9cWAHL+xB
9UaURybMQ7yAyQ6MB8jdCHom0CCypzhWGl+DBRc+6ZOjGqw3ly5mxdQWsXdeaYdXFAl3DkewBqRx
vglSrcHpcns3J3x+3ReUYc5HjGP2ECevNOiZydnzW4f8IdtvGClYTbBSHZNUG3a14oUwF61BVh1u
gDSkgvfklVTtt0uxIFfJlCTsE7FGiyEURnUbCW3C1LyL8ITM903NUQLz0sm6/rfGp+Vw6xVx75iW
zWskce7eCNrnAnuwYVS81VevraYio2nrsyoNoKyIFBVaRAWZSV+RdyXJ87eDy//OBZsrWieZSDue
NkMGn2j5ulV0lFrnAmpQU4aquah4QrHDs7UD6if+M3cesrrHJsKlyZShsdmz/6DHCBz5eKoPfeuQ
ROo2ni4f1x4HmuaVGQfcoWRpXG9EFlW1Fax/g9Q5vxbDWgBYD7qQgMpxWBNT/TTB06k9KUctOUpO
r8QyYybytehs+J2IEALbZbjuo40BJq7utvVFutKmftLkINJsAQYkeSpyt9THs304UwH+Yyi/057Z
2LyiSMVx6sdDIF8SVCSbH87T5Yp+r8p58ndU4sW+hz8S0iRwDASb+I3rTW2I55l7tfD3io3SBhaS
WlakwMEuKFntnlRVzBpKDHfcSdD9BydT1adjoPOzw+XJUevZ7Pe67e544stYl4b3A6Xj2aXoJdWP
wChtfiSQvptl2hhLMaLlTFKosFOfvAOPBSQ64rBCrIASVePK1HoQAwwXTM74IHQNFs+GuP38+JS1
4si4nS81GmdbyJ5vtiKeOyN4ONThHihzERAVYNkNkMol0ClMcUmCOFUpc/8dmdMLVgxEmxCwm5e2
SGmUNgSsVtQgNtqGLM1BSnV34pTkSBAw71EEpoNiL0oQW/xeLHjIcuQjPWIguOZJ0c3N0hcm48yo
iMBy1g6k+fVAMQuXTkTxmSj174bokZOJEDYVaAvNtdV2L0xrvTVBtyEvW6l2Us58w9l1ap6mvvGE
C3nDfsw+ZZoTG2MTA2Mng2B/AWQ5p64yrPXhec862fGGHDXVm1Xk57R1XMnXgU5W/JTFYHEO4Z1g
AQUjLWLtNJIpo6/fbcs6A0+oiNdx2woUSSzrCGHUlIvoFH31wXUQnrHHTPpoGK3Yi1W6cqc1V3hQ
Pk+g3AfypZifqdxyCmJNxMlAJXcsykQKE8JjF1kN14bn7lgjv5wN4LdPQM5JXe1SkIZY+7vw33uO
pOOUhYIORFjSXxEQ307EnaiudDmD6JrRaRy0pbU5n1azv5+Vzl9mwg1FSm5oDkjWHPD7b+puvX6e
UbcXDKAZpbGTwUTXASm0/+2LtMo2WCLjzuODHvXkw7+rR4kZpokY+8MP+Wg2UC2Zkxzr36TfEoyj
4HPFrcdJU+lAn6tnL5Bbfh9AcPojfuB4gmg1pNgH4PqDk7TvgKC04ZAfVxR7Cf26GxaEpB10OE9Z
BxbL90/q2pJkEqMqUABfj98fnq27du1Q+jZ8iOvdOnI7YLxqNc7ZJdnUJVg/wYk4BWiQAWOIkCY+
nf4nFSWaKnNxHmKKojJnL9K5rDGQCODcGdTXuG66MrzwvsDo+MUqFgpnRO6QO5AVMeUKoDGfD59I
mwH3WUKxONo6vfgEKyf4F6OXoqGTUzOBuuyQStU7MsCQKSM/yKyl9WL00ZV+uDLnZv5XvL5Bbbr/
mu7W48TaZzU7KESiQT5eKIOu9VCvOVChpheXPuQtbu3g/R/kcx8uiG1sOGXacU0iuf2aecl21BmX
2SIrfNb3lFXy7J4/Xm/D8zrP+rImiLb3SluccbrshTRLWueOeQ3d6yz87BwJL0iNs8Zvf/KciwVn
cMzWMOfx/H7wFCm873VcdchUsQQRbp59QSbhQzxlxEKDjk799V4P4uG3pY79r9YIe65XYqxXlJsD
k2vvyy09+5tVU4vX6lidXjPlUgzT1FJ454IaeW5PasOlGfFj9i9HThWCEw87Y+a6edmHFIaTEPEF
OzHCKfajlOZcDpNIpbADkYKFQqXDhWg7DyFHPPPxtuCVobrURWjPjPt2y2DeLTbW3WbdomEAELGy
Q0oC1vdGM/fkjPNGCLj6ESpm0F5ZiBsAT/CY+2NTSYr1RudiJnG3W28JxuZyDqGbT3AluHaABgdY
7fk+yIA11angwBg4yodBlIw6jGQFnmllJGknX7M3T7d6jaN1Rsb/MnuCPnE9vbc2jjmGxftdnEF4
QTVI4D0ovmWC55WhzK+6xd9sJebYcpDjdxLuUe3RZzb2gWAEcFQJs96UW9ihZDOWz6JgK+MP7fPg
Qpnnv/qkMvVUqTjTSRpDAyb+erI68XNjnTme6gElU3rLMtD62ogfJ0Rx00s5Bljl2p5qIPhY+ZX8
UZ/b7iZyjlngXZlJDTzcXbuvAo8j857i9pwl1PNEl95c5A5+q0lI0CllTGJ1ZpXfZako76UVcOEr
dde2h0QON8gBcrdTS8J4nCft1Nm4RthbdKAU+7p5qFYfD2GDG1bFZPTCUlBET67qpXQkTQO7AG16
l1rR4OvMnC++hUjrma9o1yrGPFAyu6Fxou1NnDDNNtS6ic+F0jECkOkh9phlz9P/q26b65fbR5PC
s/rVj7busckSTKey4tWqJqczSXXs0hhUJqs2G62Jd6akWS8a9YBlUyqnC3pF9kl6tI+2KorJrSsL
cQzintVzlM+fCvwQIH1/dWtqZvrW+QKcj2h41jH7QVH9wljXSIcBWg9JiPWkw0/ISuR0pr/ZAJiY
y31bd803Dly4Tuj2BFBjUbJ/hQMj1yumtWUIKxlp+V2PclcqAgdCdov3hNt/9lUdaBRJuY20aHQ/
LrbcICPFhxE/Anh1YjNf4Cb4zcA9neXjfeNbuhb1DgvZbeMn7+IM3I4d8sX3bQe1lj21xfelRiE8
0b3Pfb+gUO6Hrh97q7qmKXt5eRURwibUQLKrqo7mnMCKvBST7nRxZs/9cptTh5pC1WS9AAUp3JP+
0OQy4jWM6C0FSLz9ye1vV/WU6DBmlRPTf96j+wgIB8Xsb9DdIARUgP3wX8G5gqP0Z6FxYkdV918b
SUPhLxh1P3sl9SHuRqn6ec47ZdSkhfgbiUDTWL4hRmcmLWSKuPpG+Q9V3IABMeXZ7+OiBzDICBzB
ffYq6CzYkX/vruPAJluqQfEtR6DsIzmCVdBmlwoz9HxLo7EHfdyCFlOsaTt3UJZHzTazOUgkpKhw
EJaLwTiPEmmiDPV7Rj6blu9SZUVeD01+4XK5WydMSiwsJm/oOoYddndt2VlhBxdDvsJDxlObhf15
rDEdMJfRjNgJIc6XWx8IMxmPpWcVmL2oaCufGMT/cMK1268BzVvZqRpsxIPjJrBr1cU4ZVNLV2zS
ItmRQHnwDZAuHFPX80qKlreKton7TS5wwp/jXCZ2JnE1uJF6NhbHEXc/BoJgKtUCAVJfWgizJ0Cs
F3fRXHBwa2nkXuPvFYkWM4Q1e4ilGmPZBTHKSuYDXbyQ14/hPIHIAB2sM+I4Oi9sZ8zY09KcbiZy
ipaE4YOFuUp3wOJZhArmoEBSTxYi6NJz73jH2MpmeA5/Zafq23AbMnxH6uucZ/NbloqpbeAVYJrV
8qn2jrs1qoE+kHBknPUxy5bw7hydQ5Mu4U1PuQDbQaGbGPJ1J28Sirul3XKKuI7JHptu7nx809i7
Jk1/CfgdmXTyRVIm3pq1ecw2eHDK6hK8SdpGVh0FAnPcVkFKfS415WQl4jC2Fk5mEVQ3kUbQ2Z+M
GJ9KCsIUzR2S4slmqwbDXKPj9wsPm9oTGCDukkKGNudduiB7xxOR19pM54DLWGyQWqpgIkT2BObY
KGXV/Oc8IfvKhKRleDwAhPzXNNrkOkKytYcVWnVCTUUGIcbbp37yBOSDMhLWBvLB6iDOtEGGpNIj
FRcVySpJVDODDOJc8A5CR1/4L5zdNYh81GE/BopUvu0C/HyqQCe0FD4bugGPsC15YYfltOVd9amy
3Cr59Kb1mOjideu2zuOEKPXgivSevyOdNUfGJFfhEw3DPsNDeGfUNqrU3RAGoCIKTvY7/REkdHi5
W/RyBOi8p5vqqasmm8M/WNfgnWDCXEmla34gQaOy+7tyYAyVHeklG0w7NYU0TxZKF2NuQ3uCcxto
+0xlbD7cG2hPFTSDyVYQOzCeR7FUtm6LIYpU/1IXo+4M40L6V0BWmzmYEstunmYNPwgiJ8EugbTj
JZ1oaegip6SmRNyCiIS2sb2idui+aMEdiqkmFX4GCfApFeFNftVn0+8JvVrJPdm/6FC6Pn7uY0Y2
U7Jw5Fy7sZ0pI4GA7wSVPAOrfu0JSfvVY8O4OWHFnsfRh4ABVH1n35QNB3Aqerm558N0Sb97NUN9
NxYbSizboXfSLR5njZX3nppKgxhaBXUT6QUnidQGx/rdCmYllPJhDarWQlviZFjX7RZw3/GgmiQJ
IMK3+QyA2udf0GwtWT7KDCm3q15aCuVEr6xh4/UPvik5czlHofYqUaNsHzHR5IPE8oKrRAorcr1P
qXDV4GbjctcwHhmAAdBpy/pDxG7T1x81CTPl2FasuThJhGHaVqiHLmQbBZ1Tf9ZtagCogHlENGnc
UZiOG6CJT7MUrRDNh2BD/rfaiEbmaT2bCK3/m5j0avtgrEOd/OTD3VHZ/6ceT26LcdT7Rxf82GEV
qmxEHnRLdY7rtbEf601K7ObUCxFERxFk1zetdsoj5L1MpNVktsyjz1nfxJoHqTU5R5461Y7TYHyY
ij82mf78lZRF2feg8UtgcJ84dW4ooReFLCVxOnXtJoMWJNDljSTPk1vc6i6uZtubTQgSOLrn4D9f
kP2yUeCfX4IZFvZC3CA+yiOaZSv00y7U6odMEyi2qRpKTGQ5KTBkxlthrmBnbVXR/nv1cgWkzVbP
IjtHsoaN21FTOuFiXvkKtRsghylitFjiVXHqyp4S5MTvBUtiOOfny0Xtr5XymdvXl54SdUTQL9IA
x3v9p9lxl/z4gzvuJAAnEzcdZPwo8ZPP4zkqyVoiWxq34isy5wMItLF4K6ueHqI5KXUwXdiEgr4q
plpw7sCUYKUklJbh/gxiitMYnaYXzoj+cO+HMCRjtrefI6k1Kb0xJf6fOl5MeIU6I1kyojS72P2S
IbNFOt5mKDpJ0pCsJRz1FlypcPMwMssHL4tgLNXDM8upR0bxY4AhGFyvWUXbRJnOt9lUDSI2SuVR
uxCqeI6NqJ1MX53YY6ubA1e3JKsPeTmhHnEl0pxVCk+mClPJF4j8sgL9NwfaJyWSZ5jCxjPK6gX1
01IqpMYlPrp1VkhF9Qayq8CvDK9fYPpmCsrBf+tZ/tvKxRTvAMck87JvdogD90YVQ7bcFGGEvOtO
gv5oiMQPd/BQqI1PJqNGu2y5RjKKfHYZ6PQxqWFx+nCtTNdXidYxN1jv0LXWSyhdEVvzi7HKYp/c
7s7oXoOxwnvM6bkcRSYvbBi5XinrXHmwdsFXR6dX6py4+n6LSqsARKg1MJqFYzArF97Jyvf+iB+f
Z3c4Lsn4RgAePhXGe8xZrC6gdFot28ULQPD5s0iU/Vi4CZf7cqUlyvSKgbpmItXaomOf6f6xVNht
GYUwrhu7A2dUrKAYt8V9h3tNIQWLU0xckL2C6t07t0bTDh08Y2drZGFPipjbLUWQtqPgEu0PJzUk
SFDeTAdbbWn906T33e/LOQtVQr0Mjj02CrQflEcE9FRlVfe42u1MnhbcH3VltKHQSoszOuhayqnt
CR41n5iNSdc53XBegmNbf8YvwqDLR4VwTAlaYWNniWd3a0mhH5tlAuoc0FvkvXHcKiy+xv4w3fhy
uVZptNv2L+PdPQe7P4GbwCGYOrOZjn4jZbslgLGxEVIhp+CdSIJr1LGF/+pEwcToGXaEVa1rhn+o
bmXojCO7nGAhdkc3bB9hNQHr8vofQ74Nc32eExqmkwvRFzbJVkyB4T/bNhxB1opQRT7yfY6Sxh1x
o9g31b2vV+KO6RoV21noUoL74fkuAsfRNhW7SQnoIANl2EaB1htSDFGHVnjtgTBaqANHEeqgU6jW
4r1Gs9tEVv1sR/9vc6USPHv8IBNQlpS88GTf1i83Vwz1xqSrQo7PuiwXauaZwH+yNxk27ecfYxxi
bHxQzCPd/S6xpOEF97VDMLh3RLpk1EGavNIL1yMDZ7i93n9ImJS/RZbTFIXWTcPpBGHiVUr0IRa7
+ydNkYz2sxT6NTru5BWgBtXNwSClHieCL2uZOvfj55JPFJ/HmUuwx88wxnhZSukxpHmRZmB3S8YY
WTqd5uf8M32qBlEkKFtRinrAT/VAhz/gPGzFtwrWrEhqCggb45Q0mEIxxrRuNe/usZv8VrYO8/oS
r8oOpLLilULWxIsa2HN0ycdb3u6Ssrdd2fHxR70ZTxC/2H5FKEgeYQxSvh3LnTeynrHbcVwvIMIL
x3jZD0rq3bD128eyPdVzrkSNbEUv/vdkMMgo2yOI2G0aDq/kDwxohnF56pT6nS0ilAYQm1Kzcsgy
9cSeGegyefg4AceAeTxi8oQdEOcUui8p6dmHCgdWFLQMou14oB5C/URXDVP3SGedNDoVDtFqixJb
uU34oGMVw90lwwHIoTnboO8PHS/1j9Jg8Yn6k4U58Z9xFAuDH7J0eQUjHjFN/G4Tx3+E2aspW7Iq
lFYpz9qHkb8/NDm8tXE30JpygDsr7TWRM5pojlqdt+9OASg1nBOvz+peE+uKf1rlhEEGRKEuT4bW
4NOlV5ivIMfNuXUMZPqGXoSl+jmB0bVK1Q6A3vjZBdkZMwMiYeu6YGnMDic4g0auCb6FmFWugjNW
VS5SK492va4xD00Tja6P5XrzbgjbfN+nV1icS6AgjEF4ts1j2OxbDyt1TvbcLoXyg4KvWMaKOiAn
+/D/GbR022B3dJz3zBiM/yCi5dGeawqMKAl6QLUOdqERS3zMFS8h3NP2UQiDtxe1kYTMu5petMwX
2wcwCJucQMOMrHU6jTvU6RDEfcT/XI71A6+PDRRMyMSJsYDghLXc1jWehNvK5c1tyGubes4Hg42+
F4e4n4o7iKSCxF5GxbwhnqINIyHDlE2dikn+j2to1rTX8ZdF/HuQ3QCgOUCnMJkflGsGj2LIO11s
IypIjr8IRFf3sOUXOO+0kIV1b7bh+V9lMZErJpWlC5oi2LEhax7Kbnyf0kI0ub+or6/ReoO3ItIi
YeusoxxxY9grvF4OdBGL08ZBbYhkRMEfW5VQY+B/gw4NdlnlOCqYvJuCVtY4gR238jlT29ZmZAeu
QXhC9pnapYUxrgq3d056t+larN+9WBiD8j0+rE0j8Q2tbQ2aGyRVFXOHkM8anzMb0iTs0tnFelay
dpfAnkdj6qDxK7aYYlR8yqG67Ige4Jm5O9yvaXGHI6qiiNPRUBZIJkUIwM9nhEQ5ehDYPNJUsydV
VNfvIk/G3alpL414bKkDnrU2xpP7s0jNQW896b9KbCjHK5W8r2XQVObyA0PDccC+Im2u/nDYVtAI
B1hMLmcta1JMJAkBHc7tSzsmnXLDILMR+VpZAOryZEpGbNBT6ZzIDCInvAZuvE+RMkjeb+0FolAb
Z6uOfWsdY4hLTlHJjfZjwfnoVcADSMVc14wYzHlx+EU9/Nztsn4UGeQY5HcV7noddQjggWvyOcQn
5bojIQJqI2kTxBKjhr8KsCLbpBAUuLcc91bpKmoPNdBcUiqjLM0vrLL89QJCP2FUvxEnpJBVHMAi
M55O1mt2+XkmGD4LJcj3gpUcc6V7LuzH58nujPxTLcy5IlJkPdfiumFqtNv+kyD8UxLlSgpyViiu
h9uB0deKRO47SabkP5lncbprbXqKI3+qX3Zp86tmaUwcf5wHmI7/MEjWM7GFCUXqvoTFDtUDQgz4
Un0E8Qa+UKnPQngAaHshcx85JVrfLpC6W1ra0rMfJEW9x+xWu047qV/AtGtLd2geAx4elg0LU5p5
XFjJ23cOsTi5OUlGp+ho2vDxbvb3DeeoZ7nsVc7al1N3DuTQPU/JciD/dHbXIc/Tlpj1cvSb7gfE
CFyL2lkiq2LD5PXUMdtiaiG05KNMadXQENhpQGIzPM12r0E3AGizYI5+00k1Ja4gkxrOrxYH6SwI
aU2JDYfN654Ux6N0Q+DIEN8Ru2itNnohjyGJK9cqY3pDAMUeMsfv2+g4UaOCqW4/z1XVbiHwYM6H
0tmpc4ZIJruddWp0MK9XfoZaZbCo4MWnLN/hbHzq3tvT33rKxTEUyqR97QLCAjTSF44Vno1UNKio
mCL5gH166bHXgs1Lx0GkEqx7rXyZ8BNTwLs34/KJZ4JR2g6dMipOCpgVmp8frJ0F3zrvkIyWob9o
4vQaLjjvA237zAWR2tKeGX4zzZudvU1Tx+YxEwPJ8+BIbxckYQYFzv9lG9tK3FBUb6MZzw9K7rEw
PycDAmeqfdlv5Kfau5wWF4cRcKNIV37pddI8u8eU0uq6dara08C1ljdYBiIAf6l0dwF5eOPliXXj
vlYYiOuAmwwycsLOwnwJRjHA0duBUQQ5nwRNHo1gaVjBxE6PKcktzqDqpSh5/CdeR7bWos7OnDfY
3nkWW5j0ha7NQkbwAdQcU0IrHeCh+bHnWDs9ZUcmHCqcNrxxAZzPkce6ncpmGmu3tHQ2QqmuTEf3
bx22nlcw4pvdaQ6+Gsq1E5gx21Vo919HRQJ1nTXVsRvn/N/mDT+x6JrbLBMGrKojs8xVHXjQrKRa
vyRfDOIE0Nt6lOzeUWHPzhYC8Mx9V/YKXBC5JdfUSVB+MMVVM4O/SG6zFYAlZBQ41bfpQlHEKEbu
phqADjREpbBxfPjqzORKXY7EJu2LQUFPfMUZNpz8SLOinB0MdAcM7QKe+bKCA3y5ycPC0MTiOWDY
mif9Be9ZS5836xe8uoV5HcyiAVfPkmT6QD8gDj8XUms1ngUrICMPYHAVHTdO2t/tKCGiNdkODCgW
uJjw1pyBQTmU5paXi43Of3VUR8HS4l6hKrGVxGgfAGn7E1bft2fQX9Hoarw2oolKOrIJGITke6WX
vsXrW5ywXV6vl7DKNFvicJ1Loz3mzG9LKSpqX4IE3aUK2O/qUc5vlNH5VFFkQcgRUr1D4w4WA8c/
3lZTQZ1dbHQJ94sawGHGlmGfuePOqjINvuvu/1EA312sMk+Trt84rkQzsqOPkq8KHqu2FEiUimCv
/prmWuxLo1oBQrC1yw8DIXau76ZF2HJyzMPtLsoq4Rr1XYoUXqBJcwTFLznkYT+kMzQNsnuGIZe9
8IkJdOR3hSY6dz+9zRoIacQsRertgTB0DIiseBzY6r2SokkwW1Cb6OOtjMy5y3ysmgeYKHsFA+Zr
LUpNSzuqVn/35dMIql46gFyUJPt45fPN1oHV3ZWR74fv/ToBrEswy7YQTDG8yUMmQc9SWn5smU6J
v4nTwJ7WJrw1iI1Tqv1WRSD9VF5dCKdIS6uxIVXFSL2lvqYdSB6DVOV5cOFewPNY48jFGLwp/vyL
7LEbMseq7ZOJ8jLGPEooyI2nGU4TVnUPbKhyX/Iy44vKz1BwaRW03z4ZK1Z/Fm5ttTpqSnjS5kel
UQpb4QNf4dSP53DtrOuf+AO0wS/em2pbDsoymRwVCUqk9MsNPoadGSp9q/rqkuLcV2NLX/1tJWQ1
Mccc4EppbSU6QYozrZNta0CeGOiPwLGUHXlASkc5Do1kTdgBJPY9M/6FuaNaix5VqS++fadroHyQ
Pi9L9ifNoCn7fIz5wKqS4rreaN2HBKMRGsszJ/55ZdWEOn/8Gqi7cLZYKRzQFagQ0VcOHPn2b1IB
MHu9zEC466rOvdM8uyUCsYAAfZM3xHi8x6s5C5hEC5XxHK12ZtBH4T7AsAGnRd0D+FASqk0xc3N9
n7dr0pSucMnVyKoYm4VYfb0WduGWPvfBPLDss3da/NNpm5cxYot3jtNCR5du/kU1E/uOtIPHvUZa
vL35RNW/2j1rYrxbu5s8MS3SsWJHlB//ztNOpXcvo8QZ3SpLc6CZ1W1t7QKUbSEtVDBgOzeRBSfb
GI6QTB9FKf9CDcHPT6IK59+6CazTcavLLBsxTGOqcZvwFyeaGZoqiTlVcOoCw0u5RbRUoaJQq2ZW
MjMasX2kLNEgMz71ktb7+IkizVJM86xuq+tYnkS5MZK7XHAdmH8awy+5ft1D8mbqCu5zC2732dbz
8hjF1XVli+DWctvRg88x9eoiRvj4S2TtgtPpWQql/kJy9F+OIdL/fuANE/RGCqwjzHRz56HIGQDC
i0I1ZXtoohyUnT8yGNsoo2u1dxJzCJgAZsiKXVWU91wOF7RylRtSOrrbV29pyO3UlnDNKJxX8pi3
laH6ujkYH6wX7ERS230z8PEhdp2VyqJ9oZhkMZMKADpFQEU7K4DsREX71KU8ag6pBAqZMf1fWSDO
83Cbw9bJTNTuB2ed7ncYYDXgntHyKrQxVpgXJfYTzNvoHZtadZsYNhuOJfxkSKPFB/NO2bxuhOLj
hfl2ufNUWqyn0A9DHMj+b3C3tccraxNLQI/ikQbW0ayhKtpId//+wOC6a6TyKUs8JArtABLbiyqQ
QTuddsS8T5309zJGjVu/gA02Jro/cOfT7YnMe359DHNSLfDI6yIHjN1rRXtQcFR82mPedVEikHcc
i/lVxNpt5/vntkM/StnQXS8nrAgSs7aXGbKWKMVtP6f6qZOO2uMjWLdBRPK2hOThxR5vjUm39c30
qJEVjJtIerdIx9iAMbZW8BFHcnNib1Jd1I++O41gB6VgSofU4O1jg+80mxilcwnCA/yrqUPu6VHr
c0drksnXC7htgYlEgwomhS9XFy4TYAeJrpgABtl8Xs7NknsmFiEfq56Yn6pVkK2usJonmnXooAHB
j1sbCdAJm4xmeEA1t84RYd2Dw9fNlT95rhPSdPe8csmsGQ9HfKUBtXsqnrXJ2SwKatNsEBdoR5HL
M8oC8o/D6EOIcybNtB8/SsFd65LSU5Dsx0ruGomDMVjKwB4V6THikiXU1utKxF4Ph7mFdvYn/MtK
aH1C+uRR6jBkodA/Ic87Vs1hx0CFcilAkFda6oONlqTtexrgcJNqDzdNkkx3ZgHi0rZq4eqrK2Uh
ZirO2NJzNJn1a2dDLyxRhVWlGod6di+zxY4iZsyq5Bj39FDTgR83ejpWH2BRmeelx+XwH5T0nSqc
cbrxM80E/PbfewkCEvJGSg3qSG0jqSoaqIJCJo2fKJO8UuOmRAJyjesYfnmfogDmnMtsq3aV1V+O
GU98ZRU/XBK0snWYka8eEfaqgYpf6qtuFKe+WpCYNm0SfYkSibIEU7XfPBjM9XmIbzw90ArNERFf
XHELpNqn8oUO/fQS2xNbBjK908Z5h0RepmW/mQm0TsDCYJZ3qKZxNlGQQ+m9NQzkvg83ssRpiIAS
xWGKZUl9DPXNsMCQVpGhIux86ihWK8zY3Q28JigEk4DsgulE2xk4DnevnBSnO9PsBlt+CmL/9KnO
9/JKI2c1/K+0awk6ny2cc3Fcgh96NNkLCjEaBVRyEvw31EHHa3uEoi878ix80NaSyjJ9vaptQJ3M
9XrIl0DICbgxT360RL12sGhoUSP6pdP+AvOYTu3lQ9RxZcRBPbsYmVbob/HTEIUEmEwEgJcwlfa8
j7xkSEfyElKPVExinK8XEoghHDQGb5VZ2UIm7DKnKYBaGWCwpfZ9FshnU6Y/x1v9tdc7ZY8pqaH8
YHuWOYFYvA4NSuFlR9SgGdD9SJh7/OsPxClhAjUo87HNjGVWHfaBhrspor99U5Fz703S+T7bJ3nF
rE3GMG2toW6BqtW9itwPdOInuTxAetucZFoC4w02i8CUVnuQxwrG8hHoFRPGlG3yF53wfS4/T/Uv
vJAqtzb4lMiHRyt/cZbWaVV0/nxJLtLPKAYnr9Al/lRzQf2u9ZefWGVQzli14HMtz0F92f4BxDks
5ox+ADtD9GMQ2cKMOGqh1a+oAgzoixhHt/A9wAFLS4lgjJeDSAZFdnxcumJmQ2g97+Jh3pF1CTQ/
sDbbQ/9tXn539rqSgCONFhBfmVpwkpqx/1SkRSdPj+3Qu1nIug8FQTL11IdU2W+J3dhLRJS8NJfe
iKAddpdcpV4n/0/e5pMhykYlSpbptxUlTq3hjbkEGYb2hu95GrRvFIYwUc+HSosY/JZGlaMgn1/a
0KS+JA9HQ8oieGoHM06S8YJT7Q0vKLuwO+ZXQxbPbJySoLIeLhnv2C0GKltYAqOMqcA8t33dJJQm
0jtnedRRXC8fa7AkM/Cn3ZNJe6Wo0rwVwL1hrZQSrjHER5x7C1uIp+SQB9jOy+3f6OQMiBzVRXo5
LJy0dJ4yQVx+SF6Mo2gfj2ZglhEl0CXIz0zIEghZrzd3NaohyOUJMV+bSvE3mcTYt+WG9meJMmA+
W4LOM6tszbAhey4ZGn7y1fdENWJvU1qLIlUmlEc0qj6iWGGvBry4y74hutnEHuecKDanw4gWCE2m
HKcN8WOM+QT5wRfnTRKj7Z/7sG+48GJChV6sDpa0+r9qtdY95DYRH8ME6cSMGbklR87Tr7JeEwHr
M1PzBU8uzATQSRgTHSRY//wxu44jztN+CZJjkUDKABsXMlTvuiS81E3uC8niwWxiY/KGEAv942ih
iSfASvt4ww4lN9rb2fln46OEdwrCLrbg9soQvvOeeWBt9t7o+FvhLfdTeQ7YQXMABmHodAHKdRZF
eDjx503nl2+lhUthb50ttrPLVHVLPZvRSVa4+07qK1SOYRFVdnYAlchGn85O/XUCi0JUhRdwOOBa
SWzAlT3KmNyy0RYtRZEEPBE+OvCkKWhEy+oLAO3q0Cbg32QtV2tz5nBBSSqn3+DN7km/rMQG1mol
jYnVhge91j900ko2Nv8WiwcaT2oSmuVMuGsQiXbE49xtBPZMnvVEzItXL3RrONMFtdTTTtMWIBid
9r7mL7kK3F8AHSKOxrPHayA/KnL7tpvSaENXYWuUrex3msZQ0UrUwA51z35zexZLVZ8sGhNMnyy+
b9FJPxt0m4fXCB+E5wtm+W/RCQvafn6rCW2UIWARJKpQDF/b/4jpoEWTW7itEV/73EB5x0VG2nhy
gM9KxdctVma/5IaK8jj5EWA4JlOTUeI7fFSvrnGIaVRadqsC1AewMTi+LNpNpKY2BiWwnz0VAFs5
onvzjNj56M2FZli5tFEp0VKzOehv2FQDR6HZ8M/O7MH6WtAA/AfqSUkzXMCaumVn7DageJdyPLnx
tbJeDaNy2k55A961ub4n9Vp13uB7XIEnBBlDuHp99RC6p+pGlGdttoNs2YK5yre7uUYYrpOxkHEg
WLxETrZEpGgP0MhpLVWVOtFW1tjf9LZheYo9JG1vof6vjDgA2ZDxebejpBrLrPjvLFMkPjmVganR
o+LdCteW24X+ltflu7WqndzfHKCddOGtmCANcJZHCw6ssFroQjeTed+v3IBiKXeQamqyicJlJoMJ
skSHeHxnWCrv4p0gAGB+s5bcxmj0gV/J6s2a8OqnJIJh8CzLngnD5NSJA9koH/mvGPMJoAR6BAO3
qmKQDXARyWy5vCNXqgKs8ovcVG4otdH9rMAuYQzZmfsp86v4ILV4KSv8o8FOkas+vhZuTLNeL90u
hMifs9fIgcXgf57Ix0OZxSweC1oXjnO3ubGBPfgDN5CoGciST/xfvBH9pV4HJuUlJEZz70pnO94R
Ss0Fc/7qqWPJBw5pYHBFzLKU/E1nfxwPv+ZDf33iBc7TV1izYq1AeJlImBf3i3uGmT/MqaSZn6OQ
I/0o8OS2mxoE7WeMk+4vKT+zd4qA0g8/fz1TFBkvncEdU9jrUe7xh5RwOlsYtf4Zw10JwWohwO+C
A21mFQDLDewgysxyUDxrKKtzuP98e/BgXqG0rYiOV6DxrNd2pycsn+SCYXbhES1SEXREnWzA0cwQ
EV4T25H4mFwTQQ9efmGDGVVMo0D4lfifhQeJMOYWLqLIzftzcvb17TSapJmgu/CyZRNOFN35s8aK
F6OhqD7CttrhM3St80zD5Gb/80kG1gY5A00N6ebLyyfTD2eDpb0NUdRuic+H3qZi9YkWO5tF9sh5
nBG/n/IAhVG4W226hKEEJ2KnCcl2g8D1dgQiP6v7P+ZfJd9yffzH508B77vgQZaEbLbUKbUaNqMF
SzXChAwIrnn7poVJyA8g+RalEiF9rxL4I2qKsHUpCE6QKzBqBWSIjJxz9+q0BBdzCI9084IgMG+V
s1v97JWBbZEcPIyFRsLygmehybgpgvNlHqJgJ8jBYEGARU+jX7eKixs04FoDSKLOfaXbVqjKoLC4
xFTZrehia6p47zmcyY03C6nLgmf8/fVzBZ5abaR8fLeWzn/tW8FUCaDSCOIv2LKA9mn6YBhilaKs
PVeav9C2zM1xWliPNsJDNlGFEDf91uzSjCCQeX1e8Wgk+eJQA1YhJGG6W5EVBCsYLSbKacDA9Viq
a5BRd/WAyglyQV78IKBv8TEb/IlHvGEe0cF0VTG29gc+sufPE0wPVpX7ab7jhh5t0zvqQ8YpVPM8
9ldUM/DX052ZPkULrv3+y34XT9dF3zjHnkLaRI4zmgP3uMyvhk7PLHrw05VwI4cnLVM1nlVxMO2f
NxRQ3vM1hqL6pyMIM65fgwr1x3QydqnoBxtQmua9d4p5Vo3an2WqGbG907DZlTcTDi6tmCXhoVih
SYN9t832IiHZ2cSnqFgPf3aDAm70IvVN5mGMj4eKqNEM4ktulEzov0FTdQiFzdnkwy5LlsSSyL6z
Lm7jSaBjDt1MWz5ZeBtqT9KNeCa0pymrvDxdtejbtuSBeDuhuBV1MewZRH1GOE4dCOWwxHNr5cKw
VbGgfBf9VBNfzX3jsvkUMTZ8p3Bp3JkOZ9yHW7v3KZ1y+uePk1p/sLaZHY2mNykJNuOzTM0klRT7
wekmtJIdYg1v0H7pLkQb2gbcOibDPgpayTp4Eb1IrULPUw1Ex7fodqb+8ZnFar+P59F/pGykdn+8
ximgaydUGvQxV5WyQzaBcA0qrI6MHptC+QeBEs5RUfrdpQVoxjfbW/uzTBkEXkj2e+X/oiBGhK54
NcrY2fjCSxEBbcbYD/xOWam9tykbPiRSuccwx9FogWQ6SuAxluNVc9sKQ4BLspaH/4fbInpVbyZc
BPZ1NU7THtSgBzirUqMhmR3xXxnlBVm6th7CjcVmO3JOqga6fVEHenf0HLkYzvejLqQm8mfP6NLG
hwsGKEbzMJymjEnQIsFD6VGz7ByeQnhsBNgP9p0tgQZtXo1A65dbe8BbP3/vWgTpxWYXMcvZUpl7
GgYR5X6PJPQHp9oulbd2ieww8sZuiUp/ZNvXgxZmM1tWIXfJkJv9JD4gkTUuI4r9JWUIUKJytiiq
EILrcujOLCP82QS24T8ECGxmL71+QzJqF643FM0jdczPtUk9vvqtDvgrdON45WZMwCbSLf30Qoya
sYUdLe0z9T/4MNBhJmrMFZJWBnFRAzLqryeeq5PoNpJOfmPMsMC1hYS3N0A6oyiCd4mrkHC6rCGO
n1U6XH1gUkjyT35cRBrLxAEBO+vlHbQFZn1mfiSyFWUKDjMA21Xuf6RYruBhC2wu2E4AY4FcVfa3
IjhyiM0i3r9SnGpyWRWW8BBMzhyJIWK781j8D/sKSTw23dbkWlGUxpvhfpTyArtF/mLviXF1ym4a
4OumM3aWV2e5K/a3zPXDz1B5F3bha1du+H+HfkMX2cf4xvM7hVKceSyRpiNW9cSu26DXQP2T1123
HbbyP407k6saxyn1fUK6NVJXYCT28AwHDcvmbJd4aE3youOy1gB1aJe3MXQ2yRxs4NshuHTrSYe8
zMZhpuqV0HaYOCa+zSpguh2fvVzK1ZWAr6HctWhL/w4MOv6C+vcN+C/kUw10VexzjwXbwKxumFZx
6lHrSnI2plGkqr2HjToGAn7+xQU8xU5Jr1SG8IFtQTw4ZFBvxRgtSPtGpmSW92ilBcYWAd+lwtz0
kCi5f5wHf7RUlCKNq2R6OiV3E0lcJcfqYdSURQtK80WXRNRVsCsn1mSQ4T6JEHkz190BVft9aDat
2HtRGlpnKkDSN+PFdAO77TmmwkFqrXv37aTXEdyWeFVem9wNJNIN0Pl1EiW0e6z4J3RByDZ+awh9
kwZ+0OcJ7Elq9vocCZ0BUB84eSF/h0ph2vTeczH4BRQ9gUh5p+9Ee/2OuLuKPqoo+gtWRq4p8XEn
0ItCiSFfby9784dIHv7NklSANG4BS4+2e1ldBcFL5QNv9lNUyZiO1DqTzSsXkSDwUk9Hb6WDZ7yU
SWTtTqMqun0HX0C+hLemmbIngt23s66C9+qn5LXbrGvJv5nEz+Uv1nfe72UojQm9op7nP7gOkixm
OKd3YjHSNnMo4HneTBmpUAWrhXXTz+55Lm1HHpAvWT0IGah3tXcCtdLBwZ/83iks+OAMkMcP/Al0
HXnhDn7RaNc2QOiv9di0oanR0nXnKNmmfi4uGy2T2O45IpTzmUz/V+tXyl2z+m6oAYEEzuEkLWFJ
UtEzJfObGcxxVnJI360Ud1YRwd4OpHdcjokI/2LgVGXYvKRLqqUe7m9aA9sa93AmzBnDi51DhOCy
Su2duo1qXdN61VW/LMfTvrfx8iZPsAp/PC5CNXPP2lj3Ul8voYXtsGmNbzdSqKRIMpOZCRVDfA/5
Bv+T+4IRDaPx/KtF6cNGyCRfUEWUQeBjzsM4BPJKdil2a+gO/7hvsSy4vMbJANqKjmHMQ3n57ZCy
OFYjEqNYX/+Vyi73IYIgINt6m5VFBY4Vse85/4PE8nzLIe7IvxrwFWiuvUbu0rUO9XApFPcdShxu
qcZd1UKu8JwAJrcVzEzZGpXiosDBuAotu5VFDrPEBrGamihJj57U0rNxfs5rRCWEeFC2uPwYhcX4
gqg+Akgy7yYuEd5DR22w8Tn7QznIMx7J3/qu3b2o2CdikUWcoPIUJk3cY2sQ4/gu9CTF2xTV8zxX
XRtlKeuwTOpJwc3xttwn0M4hw9fSEmg0aRPcNODx0+EyyOhX3KuhdKIvU8A+GIKJdmNdHr5Etdg2
vCB8u2DfFxmH9VEGYHMEsNl/+95e+OZlWwDWe108WISHp81tT3t8y/xhz0A0GZRH1xYD7BmCMnMM
vRUKREwSQPf2CG2hWhVEdS47/BNv1RM3am3SxZvJ7lIJZgR3BWkNeIK7nUxCj0+kaVcs4hglXYfP
INpGUvE/gFO4ohieuq0plVO3EJJnYMDDKQPjxFeN+OHq9cUSLxdueOKgXmV0lxhOLd84DDuG5SwI
OPh3mOjYGwpf5dXy5i3Mqzcq0OtEE+96o2rBmkiyUpeO4U2kTSnQvbyJLo9V3T4jtERU8gPmHMNj
YnXK42xDLKxsJK2LUcSJBUuYzR7FlMOkDBtQDmuM+LqnUEnWvgs5jkz6s3hIWvL0I0g+SfweIc5T
MypRDURbto6zad5w9TISC5qvfQTULQXYLqh8b//gSwWRNkDZVkqil48a1D8bRwoRnBx3ovTiYqar
5g6WcboA+sD82e0iaKyDYKcK3oGncXhqtXX4d/hiuOt9EHum8HdO/aVsL1afhGUq5wMsXjqt7SBY
AMH3dDXNwxJinStJT9g6kHSUGQqr6nnYOO8C8PKeX3+JdB9onobkq6xW/DRtvD4+lMl8WZn1YAvm
yBAPmOJbqYFOMaLQJHIrq4RSlz3t1Yp1e6Nmi4E61hlMxMuNnc3oIQWar7DqKlFBF3acr45Teo8v
op3bydo8GLDAOWgTiW8GrAr3kcPXIOgpQnhMm99A6CMGuNQVDXt7Lv3XAHzKF6kbjXbtA7ctt+IG
mDWo0SJCwfEUSelteCJBCYF/ZGKAIoAQtxF+KZapqapULuAX85uGy5+h8DIoSFsPz64yaxkq3IM+
Fi17nWs7KE5+tIQnrvTNnZ2sfz5B3aIoss/8YqYooo7Ti1h0c3tzP6cnQvY1TxOBqV8JtZrLpwVh
gq9aXf6ZzG1aZIxrIZkxmgpZKnR75FaVxkA4snWPqLvG8bUQUIn7GTljWpujM7EquACqQlojvdf+
wgGRvoExV+ChQIzgDlE0XW/1LLOxczi+4NKmwBytNDOglK9bL3zU31nZGgQ/SdeNS0ooUeHrRiBm
aDM2fbUveTnVK+K4+YfQhR9Cv5oun1pyabk1hqn4N+CE1uiz9wHh4HD3/38kpg/JqIDD+S6khtmu
77UoOEiH/VKd7yAI/VTwIbWZUml3vnqk1lPJg5PJBv5piYhDEUKEX1MfGtJoc1L1pFhBNTD+7eNo
bV2FzDnJydAWyydmoo/m72Ur8eIyoqOceefKpFVNb8UNc1xMxvCJiuwmst6AcE4SxLIsMYWXCMuL
p5VrGmmZxTLAWqg9IETMeI6bd5T5Mulmu+wmfmYijaGlQoxYOv/ePSAP2z6+JezT9YhL1jP74EYL
WUmLFOpra73ktJkFV24SGgY49Agns5zMFM+ICbRAEsStiH94XhESI+mFZF2ygracS7fRhV/Yu5Y6
S+v6I2KEx6uBnDojMm9SL9vlKbO8Qie186G7jDkKnncdObnNzHm5xZmSXbI33rVFnAk2f4RpOwZI
YWSTlAOEQ5k6tSem7PBmvpDD739y16MT+6vwBZtcjwoiaTx0xb641CKV/jW99HI8WWTibYTxnoOs
FuzlCljDbHQEs6AnOPKKqKvDgTHvYkK+8KNumB/8B5vn5a2wxm4gvxdTPWZ01pAn/IdxMeC4+0PM
cLo18gApHMCavsDywhPD3E0RHcJg1MfsHKdLqG8IiHvb2xeEx/Y2nDj5kZT1/DN8EnmNZQ4RhXd7
kkK5feTUKXM6PJ+Mn9rWIKEQmJZeYF2KO8OEmJuYGYaGL7I4khq+oP2Ku5tqqsLW6Qvb89ND18OW
ElMeUuO0WMImcBz9sxQXa1YkvMLv1U4FUfYwyyQLapMT4UEcDeAQ1ceRKV/RiMaZvgYmWDodL9uK
M8mwC9AbQH+0L1HwvXZO+p2cMN8pVFT0nhJ/Ic9JQOTr+j+ygLcaW2PhCcqSjPhWfjFoJprYHGLi
DLSRH1DZQAJlY65m58M1c1u4wg8LD9HoFReUF9oNlR8LcGqEVf1T52hQOpieHTYHxcerDdegG5wS
nT8AxRTOvESQAT6Sjiy8qEF0LEaRDJ1Hq/3TJYP+ZczXeXqKK4lC0z1DJ3Go89xjQaulKlh9YKvs
5/wJQBD670mgqDMBTgJ8KTGwVKob+pL+3jNXwxhEjbJSi11/MIntnKWU1yxo6Y2oxKpBiJQqXnhf
ZKkgmcO2AXxY2n3m68TSOGf++3gglSKju1oxattasO9oEpR2DKEbeklifOe9A8NEGNRkom100vrJ
prM3D318GUGOKsfLnLcA28Uane3zkSsgosYYZqhHWas5hYEmO4e/5XqM6x7heZe4ZIpVJPwPuw7N
WinjrfBE8+PsXSTzDGzvbs+GcFse4yHVo7JcFNJOOi+P5Rtrvz6I4HrzMvxk+qouH/hZ9YMrVfM9
nru1iQxiE/XSR4v8pv2k6ZUIGL7rAvgEckSI7piXWrKfQ3wwYGBeL5d0Um02/aCr7/+GYdPNC3hF
sog1d4SGKCu1YOpdHzafhoxSi7LlLffMOAVIrK3Qx6An8CKgynaa+ptctl7Qvj3xyoyehWdy/XWq
L99/rmAXMurcQIJ0HoKChOCnpokp5bp/v4qg2b5zV5tWnuq6a93ZV38N/vUUh64vtIJiVahaO+J4
1cuhcjtPGkuAbqhXBcPV/qu7Vf2on28Nim9NWOPAEsEJVK5DYZo3QJGIeLjbsSl2B1W/iE7rQjec
G0vczVEDUHRyIJb92K5P7lj7SF+KSmvhjbYAyHAGrZjWPtkq2YaNRSt0GRisQegKGhgM7mJOwp+u
HwHb/iHNN3ShwI4hOiDiNodIRthvopuNWQNiqEONLKifIH5hM0itFCuPLELlFbY+CnXBMsQZ/ck3
2KETSbkYTsl+llzLswnR7HAlvFdprYM1z0++MJxRYoDIlv6LWXCb37oLZqwWvjDEn1Fz6v8eTRrO
kvPy65VUupWd/Yv7kynk6INZa549To8wl9GeQFbKNu3DZ8V3x1lK7106VBq9W0WlVIs+hLhllxM1
vcyot9+ygqowL+uz5ALEFtEI21SP2Yi2peqSAQ8fHTm2ubaROTon4JE1hxJBHgoLYW6pghogP31+
E/K3OySi9TAlHzv6U5k6OBpzVdk+oYTEzubrzZ67RBkuBOTF8WwDn/jnR/uKuSpq4AWCuFg4Fvht
Miq594TVYQ9ecZqknyANeQvTjp7rWXpl+guR9hg8ESeBstHEwOO1DZEihIz8XJRtqPcE0h4pLaJ+
+kHPEkJTp1lBXQ0Zg89S+3GZT+KYp7UquigxjHyutf6PIFFv9bTnibrbOvAlV4vf7LBeX7n2WQqj
h2yrSTnj2uTGPtuFjIB/a2mdG/iHPaCh54pjbOSIP1SZYB5VXA4MjCX7ZaoeSaYyBfpNfH/OEB4V
qzr9XjKZdSQPy5W+xEeqBlS+t5ETPWEUSI5NeNgoNbhF6Tf/40hOi6RH64daafE+xhTv0rPpM85U
y4peOqwRjdWts5cmHFpoLPxCVUm6N3IzQj3UfrOHvFinnLKJvj74M5emHtw5FKqB9g0hXs4BKecM
NlS+KXsW8iDzZLJ9QOVlmz9PXqz5LwkIfGRipyxDLmVLvryryDtCUBiZlD/QoSHx/EG3u1CjDEAH
7odvVdN8j5XdsnuKjlwaLTbNqr7tRshoe+l79eTbeOBTCGqILSgw/el4QyTzm0xsqnDMRCGEfqrS
uYdJUbS+5jQ9QPUkIjWw2nVX6Z7d54ICBIJ9d0bXQesRHOqIzSogK180/Idl0aHiBL4eNosCnlKL
IdNFyCusajP1hwM6Oez4aqqpWRp8K/DR8mxAwJRwFXLeYYT8zFv6RxckSKfqDk5L5eKmSTztemRz
pYm782zawANL6DzamxtgjN18YHC0+ILCrRUXdTCzWOY3wGUjNL9yQpvN1uM+SXnLe1KjCeGGok/z
HIUvBjoh24bwJyQs9nNbKBbv33aIxtrtHru8ky6K6f381SeENaQZbExmCCRqFNp41d5Rn39gGw/Q
z40A6sKHkoTfGQ2wutU+wTnqZGa0gS5EbxPlHnRJHfJJUoEN8fzkVomxuL24mpPzITFGAcvwCSTh
EUVzauF61ZW+YfaTWU0K6Mh0rjCz06/pPpSCvo1+8iniMy8kuZn1ujSP8bwlR8P6BkW4+9yY43CA
k98sI62h0RibbYAoQ5AJDXHFO8rZuRE6n0IQrEg7DdgX38+EI/OZOBDnGzo2Q0aXA5cUfge0vhOf
l43npBsORxjwnkLrOldpzqIbWuzm3XEJfQqPM194OX/ykFIU+tsSJ6yNQnzaWjaLgUB0NhWgGpy+
1P4tgKN+E1VaPMLBMj+xLpCbsv8CgUgNMRh5AFAuXa5K4gKk9KbH/Okn37FsILgydm+LkIsZFNa4
aX/9fyMp+jGchu3kZgrQ/E3uaw6+uTR/kNvRrp+BRI95nh0nh1pwVjA0XOwc2kJmis/0PfeeU0IM
S8HFB0tNjiUFc+Rkdo+PaZyaua674EMFL+h6Oy30jbMIp/i5jOhNYDf/nDy24TpM9g72tfcGdHLq
cw1ONaG62JHLjWewUXSAKGUje7T3+BMZZw+3UxFF0HvVYpt7mDPhXvACnL0KjNhlf621vSZ6bdfX
i/4T9XjouY300QCNMFkH4nK5HmwA1Dhr+C1RfpHeEAMnHVOyzAngU7ZACJqsbqtXAhMLKSc37p9Y
I4GcmWSbuvxW9eQ/JRCDRGZ4cKj/JHIW+axHqyxLdpoK+qldpA0YNISv2S0y6oBmyy4JHWnzWFwu
I+atBbzt+VM+l/fxvW4CNJwVeXUxXwzWDvQgZBXkkO/elJivE2aOc7b28f2bMcjRbgMMd/M8lVO2
NWHkTfJ2PQfbYK+qEI1P7pi90D/9bdTXAdjudniP/2/1BuoWI1wiA8oSJD9HMfjdQ/oWyIEqY9J+
CwRT0naQtMoGAvX0kfJ3q3xam6yYSHACAcArXhOOOh9pUsMg0YNfkcO11Due2DWZ7saDLAO+4y8h
WX61kAArHr6awdSmLM+lRqeNOhiDnZMOopIdtb/VlSCHd471/XIdmkOYRZqsAOF3x0SnJxcNeC4x
7rnuf1KRBEcAy6IUgvCPD3Kbv45szF2u/jy5XmHe0lYsI/keuDAMSXB9DLQ9fwy4rC1YL29O/kuM
gKy+6Nul3wAcuLIj8767EzpTYzb6lNIwiK7/Csj3d40dYWU6+NI79k3dufqAAzN1N9bxqCk+x/vD
kQhc9QNU2ZVEcMtRwewkyP5Mugk2go2/rHLDgiF7mtE8jIBQWp+5q8+SNn3xhc2mU3Jw8ruADaGe
fNKcm7GFHa6KUeidVMSUqs8ZLMovdCL55KfVNIzYAM5hraDrSfBjMWiCDQ/2eohWJqmE1NrUep5J
fkGQRmbscZOucKslutPFT00hRaWKLazzRgkVgxHRPhFTMU94oK0YxtBl7MS1t1SmBP2Nw4yremfL
Y+zfShBPk0xp46FL823f6+b23JUrpNDY1t2BDlx0uSvy8AxdrN5Qpk6XiKrAHdGCrCx3gf2lZRGC
fgQAQkHxaN3+E60MqONmktYMv8+mrA7UJOX7ITbgqCIcjl3WXjkKtDgySLBI/bTiVpVoC/6l/O3p
E95g/YEccda1WaWztEyLe0wxCmkzMpH3slUkcwgECP3quiVIGR50TwmUrqQ6dEhw6qIBzgbEYkly
joJWueCylmazEhyFyrxOaXg1Mcw+C7R1gD4KLT2+baZYvXCyRwArSFGhM568figirSnKwa9hDUEh
NHZ6N6Ylha5WevizNfVhX6GASDbCeMn0URXc1kwQZn6dCoGjhwJSeLjfj9lIj+p99jdm6WM3saDz
7JnsphKE7a7LQadr33DZCHyVgxfqRcXoALaW9+riEJ3Y8LRBTEqjDU4bh0s6CqyZ8B7iKRzXtYAy
9z4iGrfhJnG7YPrDt0C7MtQu2RgG2VJVRDOZy5VFS7voNavY0G3lQ904WwsVU6+PjqWqIUyyQfDy
rsxaPcph4Ar4DmZExaxhhjrgOM2RCWOLqrRV7hKloski6Vla51DqYZFos1HUntuTK1RoB/UL2FyS
E43Y+Mj8CDua3PhsNBFTPOT1ZdCTjuwti6ctBnYmfLIwlb3q+MXTaXfOLDn9idSrKHudLX+qdlCJ
nRN4EOzOFaLQt1JyxnklRpt14yfCNjD1E+fhTYf0DaG6OHVS/qRx/9Qfr7/5jLWHviEjEtG4WK2y
4+DrkmNxADnGIkhzlmEnqcTL3MMORmrahXREP8FEooH3L4TsHa4YbSLLCgdNtTZjmBbQ7wUq2mAj
b3V58zeJaZeZJVk+9+q4sAUae7K3mUw229w1A1ZpGGw//AEPBhwOA53gmUT1PIhzcz0ce2yKSyjH
wbuwzwNNK3ni6vcjGNcEXCliv1h4PjPNhhvR5fQ5wCUTdDUG/OTnoxRU953vAGacniojSprtTxjV
njfhkJjvOMYdiUb40+40m/FyivX3puyY5X3DfTxkTUGoxrprfh4MIjGgLMFOzJ6MmNC3psI990ri
3I8OavbD16EJ8o4s43cStjLqcrlnUigbGQwJzkCcCrT4fQOy+KuvRPV2tcX+WeyYSDWta2p+s/JK
b8LALMKsBsKBdiQhab1oS8qAx3gN7PBkHUH9EYAEf3hC9xdELvrDeERv/euynqDdjrVyDt8cl6aK
M2P3orvNcsk4hqT2aN5TwvLNkCVfpo67nJ4eh8kWS9YKwN7BHnLZcXYOGhkOuuWyHoBX15ZWHKlo
CO1r3DCNOf8GLxTqvFAvu5MqXKRemUI9QlL+4VIaaEFWYMmwso6f9vnDsu6KHadXP8kG4thlBPnt
RUY1qmfdo4EvedrRhoJr51QPwoFO0WFakGctBW2YRJUFrpsGP4Cq3GoBSO9O1LkuzmOc+YpZsZOc
4jItIB9vlsfukaiklgk1NduPQjoyG5sJlyL44+OIE43CMp9pWEpWxc8TLS3VGXqwnB98VCOZR7qV
hEOPMMWsqwGzk00BOsb23UUXJFREOoweKuVlU1p9YA4/8nSIhVlPxGu6AiufVAx6mr/odqy0DvjZ
xjtJ2DoTRwPea4n+akfqK+5BP9O1PnDgRY5Tsz1mBuFSNpZr7OOmXaDzZRLdCC4JJwPw+yLwS5Rp
aUxRzRdStOejARVg/zVCenjI//HQ5B+qdhh7YSiH7ezSDrARsLhLtKCI+60UsZ3b6Q+FyDZfBAhU
yU3BlqxrcXJnXO+NqS0xppTYs6Gsbq8yTRh39SBgeVhjMopRPtYY04ZZVaJJdz2AMNxuzs6V2L3d
Dgx2bf3hH5/ry71lJAIaHiz045cwXwUysV3rr/VDl9cc+HvV+9La42xsErNZMgY8sHAMQY1VFMvu
jrx/wclmFbqwtY4C9H79u/twJXrKEF0LSMaIJHtQbWndjVzSg0KPrD82WQc8ELWRFPYPP3Dby9q3
BYEtsgRRQELdJAgPph82zt31ypTqPQ35CBYdN2krjP5xtf2y9cPSFqrOZz9T8xrEqyOjQXMDtabb
orlnIUwsDNph6fWqALhJLYu+UDxSxSS8oL/rBpLtygVgvcANfZ8Z7JmCwRp+JrOPfVCM/vblSGvu
YlAJhdVRCd4rQfLvJ4NfGB5O9iCdxJNd8TFmBHDYF85wo/ffD+//tGjWACLsRfRr+eJ3ElPdpPrU
Z4q1u0sU9CVbTIB3VoQx8vhQiCCcZ1509hG8AoBNbI0495sRxClEBjALBD0e56oO2967j8EFGom6
VZs3VLrywO6zE/79zlwR5PF7/DyaIDj1C/r1arwNWQ35ipt4zEYO8dNwHZG7zQhRymUi8+ljIB8a
I/9jL0bgOFtqbGhQoR9DhKx22FQq+ifGUrM1Ciyz3Wtd2UqJUjCwxxbe1LxA/0jHIMsI/tjDhhqf
pnhOeRXu71ph4HNBcpk7GWLr360LoHthivqlO7XnUdHv+SqeiehPlrKJ22FTWKGRZ1lPPWtv/3dB
g//jE7EDj3LaG01p+DL0/TlKtZ2AldFuA3HE2V4z02atuLGdRUTBAVS3ATB5C0jv0UHtHs5fY2XF
SSlkXgvl8ENoFkZytUJwTFrlM+ZrLBenRzXnrc+NT6m2vs60hrwyt/QPZr8En5YMSQ/B2AR0MVIH
PKmHZTApxcV9obO+VxfAGEL11RWsJfV+k7lim4/pS6aVHALOReBSuvf+9OcJJ6I/EVmy6pxfCUTg
m2CVpoLl2xynViocEHckruLPc4ugNl5Cx2kxakm+phRqnEsoK2b2PDUUs0ZQM3eHD8ONfARRYSZR
V+wBKj2xnMEEMDcEHtzqu4ATGioTzrylUBx590Ypb563X48PD1Zd2E4HcMah3iXGb8m/PTzCEEfT
mzVfnSFv+exsIQh8Ej1qqAoOtVsA+aXi3D/e+XKCMNIk2nBoprQndRjyyZmkn4U+/dFTQlsuoj2l
59SjFaYG5NqWaM7BRewD8GooDbpjveXXMH5ctFVTMqQFCZTRYjDtZLCQStLW5J6+reuuc0y7PFMO
BhP7kdVk1CJwGjdNAaBcvy/Gfpo7qV+KPJGzcPpgu+IAFcleWgV0DW4y+D/U30yPdhRUx4Chpgtj
sKApdB1kQBMKOvNaWBdrbSu0e3qcFwC+np2EuSEGTehYdGlljzkIXZsPyVv7z8GKl4ZP6xuxEfH4
s+VCKgF5VEC19CvTTaZJvja6+0veJlr7JTTKl24/HX+KXdcl/L2qhRc/3QcVuveTRkzTC2lbJcMU
5YB2KfkDUcVCQzYtsutWxzc58nvBQMzw+8xWBtwSY/jTGzZEY3uaj1F8qKKO5LvgFS3dlGyqWzGC
jfRa5iNVfQf53yQAw8zEKd++stIoIvhYGsK/tC30hrZS+lgjNEY2RVv0eSqGPyhRwCjw/jVQPALA
gF5PVMMGdlN/MUa3pLzGAT4Ryjr4RJ/cYeKxuqM4iJBt2ndPvSNiLhyGOnXcjgfEdWlbh5SDI48U
lh+hiYHEQOoyfG1P1Bxn882nAJUSwpQzAwgOegwf9aawSHJ8Md+GWxEXMBa8U5wPOxSf6CN0FD2V
aqYEZeaYXtWZStCCIhe/RpX2Z6F+4pLY5/nvj/SM/W5UZCzDhJFqbtjeLdr1CKeHDltkLD8p7ZXY
pSbHuNwyszBS3V5RN/DuKnyZbkOODZ6CM2B+25a21M/iSF6l5uRayJ6hOko3Pf+dSjm13sNByeRp
xoQDMoFE5+HnZ5Lf9jKKBYqAkK8W8RA/Fz/PAwzr+biNltCdMyIxh/ULcqEi7ZomMSBniOQTN9hS
tzdceadFbsVMcwIgO9+M4p8k5essdsCj6CJxRNTGeuOXzjBulVF44GPgIU1rXh+VBQp5VUie/As+
ZKPtdp/MoHtd+8n7g6ZT1pBQE4rB1JYL3S3DYpgtUEOoSH5kWzhz/eCiG/o7OP9Bmfz44uPJctTY
s5kdsPAitkETRS0DxgAepT3k/fRfPg8fuaTDmlU6bwWYVEOVWCsZy2yHeajF6yDrxQH33HUjp8ty
bWjuv09FKu/hvMRstIhsJsVAz8NJoShR3weTNP7xzBiTqIrsCRrcbQCvfOrITFXbLNWO/DfD3Apa
KV+QErlRIADNydf3lM0H/0xzQNnx1RC/8dUKh9PGDnGnVaAAGKEQRUM+CinjYp1BekVL1BD9xnY0
EqVfGqsD5rDRkqSEocYmGUEIGN5jKVjoYsyHmBxKAAwKC+yGj+t58k+33bvGUQqCGvBVaxkM8hFl
6qUjrIW+LdZJmo9O6B3pqD6ADjd3NCe+fDBZNvUP/SyqUfeQJvHxrQnbVZqEuC1zHKU7uzylyG/G
c0jqqS72AFf68/p1psaC1nr76d7UfgXpUwcwL0+1ymlmt0zapDsw5MPjN00oS8Xx05CPaVv8QGDZ
rFLJdjOZsPPcso8ZLxwaRA5W75T4L8npzw6XmTnWDJUcuMTXrh8lXexmJYLYAGLa0FsyQ4ZLqHsZ
C/soPqkadNRW0yaN4ktphsIorTdYMeTvkNU837CkMAa8V5xCwqOkWURRcYo2jpbuhsIVv2Sv4L85
HqrCWFOSWaOMdE1U3dvxe5x2YbhGJBElOj1QnCgNIoy9A7IGGU+qAI7A1GGsurWTEi11fBDAn25j
ElMtWor5/xoD8llbT75myT/o73nUXmDmlqWJAZwUZDJANsP0YNCYmbBSf2tKKIBCPOpe/UB0I1Fj
07oiJCYvLFbSEep1AOKvP43GWAysAQtpZGShb/p7PlYZuu6a8yM1Kfe5CYT5xyzpYseaJja0eYhB
1+JYbnlH10IagtBwEORklYQtHqoaSFILlrH8Fk2Z0l19sh5ccNwSmWy+Yt+IZiB/xkZhoP3H9rSX
Ar3RzAB6fx0o+Qe1cxEn49lkV4R/kMtBmCmml+p4CEESnyFqxVY4UTnHrrp7XclQxlfLJMlrxMQf
2LQYmFWzGM4xg20Qre3MeRwPYFlhVX6pvXjRatE5FjUJYWCLxCYbJjnGTiHQR5S+rOxjai5Uzxye
sD0XbQNB5nwqubd5F3SyyHG56gs6lQOC4v09nIvTAjI5JkVRcLgu7UBDQ2nDqlDLhY/oNfrEZ0Qe
xAdjhWANNBMT1ULlGP/pSdWWlqfLU1UmoJDs/jooKzqyqnST0LOoGie6kZKqFiddgBiGUT0vsKpM
aon+wk03sUFUAYTCc8SRYvAXedY028b8S5CDB8KlR6N6HaeNVePQu9+lPqIHWBUcToP1/3wLbgu8
9X6nLVJJ/r7rZ3vck5BuoUXaktvu+xkEKwYV/BPJGZtJKdSasZd4Vrgi3R2hRtJw9UHZVZHH1OJL
Aa0QgWlQrHe/fFPWIk0dYONF4J3z0V4tGuS+56XhE+2TloTqSjO/2AFxAPEOajBzUls8n+ZygCDt
nzHeJcQhVI/7dVrMt0iZgL3U5cU9ftTuJ5PRe9Z2eLEWieNGSSZnSzubxVjmJgfi6oF0PvkW23bT
ZRCTZNdeAZ1qqzcsSf68+VTHBUail7g5WXMZxK0C1ElUixCchqgkufDyFZdYwHY2mPvys5zSmzRS
l12Tcv6gAgx0N1KC4RRqN/I+fmOj8bo4y+ArDYwXTo5dSVDaw1s/uQFdbofQ4gv2MLnF7Tz2EiPn
taITlroUXhanefeKAyoApRht8QOVVXP0UlsgDQFHtUEjMzTYQ1SEQR0AygtH6n5InBgGNTATadNa
qEe0rIT9h6r/rtOdqvEo3MS82fipND4VXm72NHk9/J3RIiDvMfvm4DDAq1nHeCez9FihqCJk7DNd
Hcj3quV75nlyNTv8wvh4ILqKWYR5Jfh6/OdH5ExmPnWkf9JcKFLxI1+wazy6xQqJOzGhgmXyfp3Z
uvVIajY5GWJZkERude4jSancSESgdla6NTNjrFCWzJZHBK2hdZw0RXCPE/TE/NN7YlssoG2+laG1
NLZqQDzHhDbKX/umFmbsn4KgxlZKexDoNqHZvoUJDXZ0VjKPKNpw8O0TgBl/PutZApiN1VTwTz7S
K6DUUNJ5S+SFX853TCkj/To1ipIHBWiBrTr57Ga9sgmQqzUmIJpCBqHBzGBFO1Y9iqkk7Hub7/v7
HbvkRiWgwCrWIhexeoKQRIVSlXQznmYe4rlFo66JSqTuSwqdaNwx3HTM8+kldkVEqQYalLL5cEGV
9ua1tF6O9Fk39lWpdhmJYKwc8v/HbykjkVHmgKTW1wzEyDXdYxlPXh82QT1QebP51fftCsN9W3lc
7Xao4/ZbFqjcN7B6CSMEiIMfQRO1TMyD7DElNXyPyuvIV41UKo+EdVKsafqdg0UaaSLHS86J20HY
r9sWhEF0j+A4A8GAXtGybD8Y6YeROqNd74vcV42pG5YNfKXT305T7U0XyI4T+eoZZK2PeevwuKjS
7+ni1J9F69WsbsSZMK5Y/yBgeGBBoAz+WNrcurzr/lnnWkjYOTe/QTuTf10zY6KPM6rtcEFBvQ8U
vSETmG3/EqGerKibwnxrLzuVvDW9xL+EmOL7MCBlLcm9HUKwIsIrIInVuh7t06zV1DGVyTtrV+PT
9bxaXdi7eZXG3LB5bdnW1JmZPoHTGbJmB+DMaFNI+jy8F8w6v2/M42dw/qtO9jtQLGJi4vEMDD+t
DN+X37BDmNflDVQ7ivrfw3DbnRZeC4rC0rbGSzrE9s0n0IVdGuZePVSfY8uNXzvmf9ye+quWKhX3
h/NMms+Q8F0Wa1lCMtRgqUR80Dk5ar+smklFjnE2w+qMGWNodBQbrdhDd2aKWqZe4xWOAkapjSiB
uXhXhJz79bx2e42bnS/4BpRw0Ud5Ttoweikhc/wRk2W5S/SERJrdUYAKMwqWgpAbK2Fm02FIVfEW
ujpO70EeTEjmgqJhGFl26TRtHHkhjYLXiMVnsw8z+Tw0/MdHqeWblnqKS5bqawO2Y5cRKpX0eX8/
s6SJJBoMPmXYD0U2T0bQjyYMHmaPPvrzFB2+7KL5lij2sCJTsp1Ep8hgvBMo9GWoYWojX9uITxGW
E4t7NKDJam5Db4+NXarr7xt5HnJz5R+u6vJJuVQT12vRpaX6KBc91SFTx1J+uLYWnC0Ev8OK5faY
7O8uEeVjimhPZY+8t+FVKPYH+39g2M1RrY009VjDMUZ/vIT76F1qO6XgRIUJTbyTfDIUx4p0HhZM
RuEIra7huq0Ic28ujciUgBAvhWraWKiLPdD2Pm1LJpFmot4vK+LzbIIWYQZgpz1Q4K8Ysbnztfrw
QRU0b83KhH7WCECLEhs/zQrKU/7pD92q6egM6Xm3OB9eVuqO7Ke2opzYCLYD3oN3j3Q7X4IAE+2x
1m+ipbSUS/u1/58FHu4Fkd9d3eA/OhPwt0Dk5HdcIiN509nx3WTZekFJZF8vAK6tnvra/aVJoc0E
JHbotn6TuWVNa+5aZDoZ1TDdynb4MZ1bY/ceBDOM4eBS8rFaY1HA/YQ5X50gEacuP4Vh/+0We440
z8KU6abO/lD6DgpuUb9/tkICDtJMrod6CdSbjm0JDSdyUw+X82xDro41LDsITtBlAiPt64/yLnXU
dWNIz6Tvur9DCs2EnRqOqHXDOKRvutvl1nE7CyWU1apYlTr5EFuHCET1PKQemUAoEqevz/EFk0fQ
ONdkY9ek3T4IvYi57yRqG4woKVMam6ac6UDS/npaMiH+0thc+4dZEKUDNlist0afJjDbFHJRzmOI
tNl3tMJSjcoEiF13DwkxM1R9wWOm9rBhxa9AosJ0h70+aRixjtHDjUytL3q/HDRM14RGyjHObtr8
Lh23PtX5AUaxn/BAgwFMlKADSry7KVkHC+9Gw/FHFxI5u63pq58pOdXjNNOPBvtcJdaTTOIM3ITw
VzwmV2xnh+vXW6HV0dCoEwwMp2IWgFDny/kGU7gC4syQMWwjIzD7mmADKQOMErQ0hLmOq/Yex14F
RkEQ6h5etN5EimC/0JtU0tUc3PR/ONYPj3IgKZDus7mhIxYJz7xHG63ID2SWwIBkpeQ8itb2q7R0
2PFiCjtXpF9iNGo5UkCRD9PHuw3hxkpkXc3XxbazdCPQhU73OOBY0C3MO6q947Q9jqY4uoy+blUc
GUjH2+k3Ztif5XxQMuWmXd8ookk28wrsmwPo9YdlT+DCVcaZGdWkoI09jAV8VWJmiP8R2FNAk5dV
I0U60cT+7U32jIeV0jUYEvr4EhUV1AiEgZyOjjbWv1SSJU4yMiYBLWMn+H/VnFW627mJOJ1BwYsO
Y8pH9zRJHjnZsSZE+ZydQcTJDRSeYG22imytD/pNlF/BUgMu0L3iNMVL4W6x7AGe8Fs1Ma4ZQ0VB
3IffrvVNUoTgl3gbXDQ9y6L190JKwG+qUv0tmm9nTayeProgD1KfpxoUrYtPYEIDLzYAQ+UQ2t0Y
+dKZZ+6/nbHqCsbk6ZkEHEKRF7vNkJhc7sLFL5guoF6zHvkRyyYFVRoN+ITtPNtesnQ4TDV/vOsW
6OMr/H7XQhDDGHuq224MqpCvJ1SE5sVYZcUf+dKzIu0hc+g3OuBdfany1yoOBZQST0ym8csICPHU
jNmUg9Drjn2+QWdSIWV24BIjB7N7rbtSld/qciiNVTKbhPa0eEv9Nds5L9+p3ivJE0F20q3dRDmd
bR1r5MuSG6gCuEYpr9s85UAfsu20/hMaE3Z2YeaRaMukELpU3sBXcTNgFQ1grB9JSJs9q9iseo5j
NKI1AAiaMaYnbQMPZHh6jo8yHYJ42Q9rDD7lulLOiot768cI16Bitt3RcAJPVqNZ9PIMF3g3O1+K
tOHycWSEMdN9IyGn3Z0Gk8viva9xs/+cG5hlu1rwQD/xG4/Ux0my2RZg4sm/xkMvDgzk5CdOMI0j
U6xb/3n0SFFoBRgoctnuaAVir1UBfqiaLy3gXToMAWRUFBVRy+MVkyCd7vu6Byu8T1b32Hov/5ir
vihXPpg8g60Nk+BPsaqkD8qXOmc1VAY5GJH19y/+u05zsNr06UQu69OIjBpGMCbNyiM9LhIUmosy
0TSIOZynL432fu53gCnTyVEQnUmq2EstPN0rOBAkIOAcluGHkdbnARER1wknetYfeR2cyDDfSzAR
W2Fb280RncVLc5wS6iDuTc6UrNrLbNLvHgKQ41n5qCVUnquTsGAOhbjlxIar8sl6oFSPSsk/y6/I
uoSoVIdmcgAGa5+NCWEsGrT9pbYnLxIR6FZHd9WRa4UbGBnLlZtgqzmbR5o7Ah3K7h5mDTKrUxCa
NDT1XLCX6IvQe/pzj7iGxK2dZbNNGptIPcuQR4Pbc3I3jDsUeif/ADhuABGVg7p97sU8uZETtun0
C6imB6cd+ejb1mu7kFtm+z2+/CPrxedQg/zQ8zafCBE7t8JLd14aIp7b3rG7nzLV/dArCYCLPYEI
xfYr0WmFXrjupBRVMDpP4qgrEa+f82c9nM+7XVTU5ZL58rIExBIfRDd3GFzUZyxBpmkUAsmm8ltD
IhDAIkAMwHQJc3CqSo1Ir6UC0Dz8mBY1h9T0N0iuBF4kGhd6QuFKOy0xlEfmcpOMGmbF0JTzlcth
rQu92M1blbaK7YEgqDwF1PCTbI2EKesSakQ5DunxWkigdRwc18eIY+QsXuHx5Tfb2QYt5kiBUnMx
T6+5hJ3ASQlLIZl8CMb6EvNFGghwINKMR2eYFSE/jAPWV6Gd4cMZb5PnNMNrDmJX6PxkrV3IOXNZ
m9Rr0ih09DmiRttG07DbozTTg6u/06O4KinHizHc6UCDpXQsxUOMVXGktVYwP7pC2sFHaNNiMqn9
HyQL+jhVRP+RhJDf/UfDCMCr9OMk2qyNI1+wG2ox/8DBpszxeMGCccVXbo94P744fvZfLwEyP9Cw
Im/KIIJLNCCJk7MHGk0pYhiMmddyWjh8PKDf6wPIXd/staNEc+gI6B/qgMityw0bNAsFQs6HwodW
C/hTxOmUheXPA0RBR4lKGWvUsD15IyjNlQ1jMBH3B/NDjRUDl0Ns//aJvwLhhyJTu/1J5sJD4OQj
4RSDRbmQyqGWYpVv0moS6g4S/aAKPzmmeJC40IWl/QC9f5JeNMEPsx4J0t5kUAorBV3QKUfNsR5T
c3Kf9wd7cRMKlXupbd+OCHhMKa5joqWNxJO7OopyskbB0VA48HDt1RrLBHbAclNp6f2uDOLRuJRf
8CNBAVjdYFZnTnpQB9gQ9Yzi2xvDduh4ZnEooI0EKHysPXIobjng6KOvofsL1CGmPhc/I2i9X4/m
UFNHXNKiJkWYFrgiuOmonoKDtd9IyQy0BnN73PIEam2hvcxd18+/RIpECtNvH3jTtX8byDn14k5T
VD5CdlLDNIbSq49m4/JUgbY/zuiuzy6o9cNvyg7jIrPJ5s35+j8OZh4jBR7i9EaBVfnKHe2lUBiT
eHFgpUV4qNYjDZ1grM1q7PSl/EG6QW2swzF7qjDXDmMY14TfjnnemwjJ2DPAVVoB6mgH8i+S+4wc
y4bRuLdT+IpxaNB3zgjzikhs3ts/i2cuqlAIi0oBRsb4/962SbHVHKlpTaAyVXFkGjC6S6rycZE1
D4asndwdBvlgqTqvcq1/JD/JNOMJV08YObLLGqfsopiAYojWovD2ioj3J14UPhMe6OnKmJtqdBUr
mKEIoU0tmOiUrdABja2/gUMIii0NOfKHGfZZgvPw1CAARvOvtLAWOhd3TDiUp0KUnnwVlEenRDK+
u/JtbcdWWBQoCFULOwEaly/Siwfei7si78HggSHDOMKkETka2mBGKQTX5Rn8izyG2zMR3WbWQmj4
i8vXOCbT3kyw+OiDc0T/wYgw+fIYtanHa7KqiM6GiqhjCowIdUdxRHAcjsVeRC11zdoU3pKP18hk
hwocHwQ1jKyRs94qYNXc7AV3JEmJaJUjPh8VclpngoIf5eMdSGdOhc30vl3xHnWB9rawShyVpTnN
LdWbTo0sWzC++12qAgzY+jXLLwpTmNQyjZEAE+sdXwYspbckL3kBFfFJ+qAHTmmtex83g7O7weVL
Hj+BT2v7S84DUNuEYVGV5uoZKOwmf+HbbjJq6K2BtsIqhvk//LFJh9tqyE/VIITIEpK97TqeTHgK
hjzeRnXNjAbRhIpyZDX4025xle0Pkq6TDEJyt5oy7H1xZJprnohLmb0uzb3uJXvMUgcE361L9uGz
o5vlpwwKNxOtvpkzU1R24MhKMU9dA1zaySxX51W2r5qXlpcO977J14NcneFHADIRpMSdFk+nnwVq
jMHXqRTwZZ3lUnoGOsIg9u4NaH3lgxqkroLgWwQC8kPt6Lq43v8nUzxUZtOdvvSgtf/zqygyjtoB
NH+OE4pskBP3xgIySHpuH0kJSc3NBTzzY7stltaWdLl/EdICw/Y4E8W5MHjDjYcqkVuDesdl8mr9
uH25t66zXNi28YjuFI5WJfA4Yuez+5f3ygGqzlwVPRtjg/9720BX4AjrfEmpBTO1ETC/aTRqvOBv
2trKeyZ3KhCbTYmmc2iwetQqRpsQv0LwJLEKknNhQF5pag5yG3qmPcqRNEmLLveaYKaQQy1sWClS
nZ1Na4z1KdAKUjsxcdNmtRB0ZtwQNzZUaxYMwqmk6MCKFMnwEfZEW2hVc21hCMeQhbF568TVmBhq
qNy4yFRLwd+AJHwmERzUa5ZDMUR7hY9Uicpe8UR7uyvgFUkEkuQfHjfpoiLB7fvcXByVcia0XIrI
L8rZ2CfXHIV+5EHfY9uojiuCyIPuHpNiH8xZtNyPylLqGo+ANUvXICVBGns71dL3cbA9qLyWJRTK
3PkvAljV/BgjmdMoh2b5bbVIQq9qE23TbbLqB3O1vUISaKZ25MzZh6oCiY6o53nsTEsRE60yLxog
9ZCV+lLDXNaxCBljc693R7TZEBmPIz79VJtFSrOLDDfllP9AW5A20s0T+3HuXMLVHjYVbl/5RRKo
A+VIPEy82bnB+hrnlPKCiNTfVy/Pu7Q2G2btp0xxIOVt7rp8Wy0Oc12q4w9zoKyR4NW1Qztczo3l
3BRp0/e2RkrUEOOm7mdJ946kCVCTFPShpCxb5cGR4SedR5NS7RBA6kP8n5Hx4NGtZQvibBXjc9l4
+GucnXDFbG/U8CgCPxDBY2KHoPUBif7FFgUfDSWbPA/fo/H01F8XCgDJV0+5ltZx67++RmNuKwgB
LnJ57N0gabZpgl6I+QgrrrsnxbbWpTLicONvgA+VgTLKd7KYdIfF1gkEtXRkaQ7hLNZPILhH99vg
3k2AOMMOkYAaNXSgnSvoLI6qalhXUCMKkjbkLn/ZIW3V63yIv/KueDWaTVIqQCWKmPcebu/BptH0
2AHIj3Qc5rpaWHqtbr96yj8eb2T20x50ctYsP6ioytpci8jXIWxfjX+30mkXwVPiK5x7G67jANUV
6VflyjGFYPYUuALBFhTCb/zUtowl7xfcT8WbtYTRzT5uPeim0CXHJdDE9rUkoEmVYWECbD2uobQa
C3HuRFVP2wvRBrCXcEnac1OELZHyz3kydPF2MPwO3dY34glB3/wj0PIOQrsBicmm87haMLuNss5g
IDz11ClmU/gIJJWaJvrsVaRpI/0wQXL9lD4sxkozu/Me3DTi+Rrm/jbeAuIGaU7iMk+k7CnWEGZu
QMB02wjJfFcHlhhfWmtC3MF4hxSZ4NV/ohH/8k0Ef/tvHr7HtHHQB4/ZB/nTZ0XtqwMpQqKTtmIs
TXUFmVUBFVAOa+tgFqSrsazayiGG1pk1Fg40oOMt0j5hR8HnduTPohzn+EydrXvvKFKvRJYSa5IU
NwIDSzrMW5elRb4wDWtHcIIfl3muysHYgzkEc+VTcmagvgjXr1SW83eDVm//76SizxAKyTf9tFXc
t8ZQS3vjHBVJ+gOxJMV6wB4TM/TowIRR8x40QJqM3mAIfsdUByyiauBvZrTTSzlWBLgp90Co5MvT
fx56vyU7oHjBd85FCdtOgablw7d5jiIVEcEG56IUeLoIP/t5aBjwUy7X+vPWPVAv5aFk60iQEaMo
b+rsYcCx67Ju89AFxYrqGoGNEtdWF6G6YsOVROuOwCUd+v4VRlQbVmezgUJbNBKmSsor3sMIrsI8
HWuka/vZCxt7srHs8E6VIhUQkPBsnPo0qKnnFfW3pa84Q1MIGKp1WOLuk4PbGSDGLQnnxwKBWiTm
ocZ/jd5Swmsn339fV/bQVmtcYDZBh2xuDd7nVSPo4f3gxKPqa128AKFtLeZ7tZshT/bKfQA63bdm
ldDJn0HDNqfO8U2Dj11rlOMO0wW3LTG0OeR6NPKogXUIAoOkl4ff16j68IRGydh97040tNWNhc5z
L0nOyqQVjjt0h+S/mzAi5WhWt8Cp2noV8nHZiP3AkGz2oGE4VWklcxu1OZiMz8sZ0ICTgZ5y2OL6
t0K7XRJr0iRQg0tt7ASva/S+1RvCsbPYkifRVSImxAqQpkTgW78OkUPP0dBPLObz5pGROg5VPwLn
FmKES6btdaCtm/E6DFAbWEBvtypzH5zivkNx1Hzjq2NOJXwrccOC0nbGbna1IfuE9Lg6DWRoJjsf
G/AXCNqxiyLj4Kv5ZozZNX8xRsL5y5GwhqirSN0PFIP6FnYpRbaRVKnZod4ZhrZQ+PbDlzzTP8DH
ClnkECcS98PAGzI3G/26VO3V1/vZbGSUJGIwfSIH0QlYGo4n18DKcP6PCIAwnQwi293kV9gi2/BB
yAoff4N/sJqIRuVhGeptBpLcyAfPNhL8Pypkn81Z2c0sDh+0Ntb3lyWb7ytT8TwmxJo3Q3atgDvO
i1Hu8KLgsycNyIwsHc3wkV/zmWPE3s8HPOGNX/GJbMkTyNwdOGvZFu2qYW812fYSkl6n94+00r/W
iinbz4iaR9B4hvfpHkvdSzcFCDUT7/Eq7lDPcz7aJyY4X83yRfF9IBXaiSgS/r8Gp0/azQojH+7d
uB2RTj3hYsStsByJNiG1/FOOzNPk81AszyQzxS8VxKPTZOJhPCuUCEbrMtwmx861R8+n6MgD6fFB
UikLFhV7urPdlZnCCkrJAdH/LJ+dGNNtSoIO9pvpzEr5C/uC+HcRMUq9MyHO7o9CZqdHB8jUQVCa
TpSpIAIr5+9ANcNY7iUxjxB2OnU2LYyWnT27wJRuDM80KrepLehOTYuu2vokAGQMi0xuorDsEr47
t2+D/sVlYBrOZJYOcXluzF1KhpkD6E6eGjFXGM+HndQd0/z9TxLJNCu7WOSEzs7X0VUdtSgcfKMz
29NO/40l9eV4DM7CNJFdnLFXFJplNZ67VxyJmqdzIHc8jdSt1tbOe/3xmyChvWKcq726AitZC76r
e8JNxuZ2r/w6Dyi1JqPIhaSCmV/ez6XMGRnirfECbz+AICePeh2EJQkNYsPslV6nLTmeWxpCt1Wf
KdshWShlI2ElxaAZ5fCuYHf39eXMCwJFo6tiK1SIIKszHhxuK4+r8BAGBgEV6YuXiUuFzm91LwzW
2wDocgNV5UGOIq6MdeW3WEevgMnvvPAQmWwi6G10GRrpPUPS5ljC94oPPLApPzcP1EctAWQK1IVy
4InHw+iHFfjA/mVboOHTYAaAJ24IkEkccZhBHkYHRGZZay9SYxqsrcRUKWEiamNJ2XiXzywlr5fm
pLV8FxK84M3mZzWd7Pfplf/KIDJSf2kEeNehyWcNmDqpYquw9s/wXpNVEJ2/3+QU+twT/1KTpQky
y6olkiV08hXV41AZNfxN8ynSgigJytv7x776i3xZ1GxUuGgVnPgCLQ8slnqkWwvk76+MoRkXlsx9
rh0SkKTXmkYXUfLrt/LGReas6GBhHAZ1x4yzIuUWn1T7JExrPUFyuzdAqoBcRuyk3bhrfprb+eGH
r16SmBxaAW49zWnpn9MeH99xKplsN7ab9eDc6uKFI0t4DO2/3cFiUFtlopjthgVLNExiIZtnfq55
aWq7cFmL4jp6Njv2HGxYhJd1o3fm5qFXUrDS3uUCwk3tG4qhKt7RcxNin7OAVni3djim6KMslAYq
L8capzXqR8ZWhCn4ewgSIaa3q2B+wVpqP1UmeBX8Ft/pmwmBs0TQsWUvmPngG/crsdYzDH0roL4x
D16ZXqDYqhlKCBh0iUOU6equJBCSU4j5AW2bkzE2UmnNEe4s/fkhbCBNlNFF+1x/8BGekwAEJBZz
0idVzmDF0NMU+q9DIYIbhppGez5UxC2mbR/JFkYr4hgyd8LgvWKcVroSHz2M6VIBWtXQI77KE+kU
1G00SjjR+1v8/FDG8trCKAKfNBGK6ZeltgUVMk+X64FXM5svo+ytdcDgQ843Utmn46rwOfJ4skUa
M0nR+4THP0Bm2nModED8KpRmTTo9Zdz6x0IY03xhQ3oEfXKuID07kblT4eJTNYF+91E28cjEkgtq
odhmsbxLlen6lWgwsmqGju6NViAq0Ns5Yw3CtIcrzxBjrILZ/UfcY1Wt+vSEtvPlLvyqjIJVYO5C
7G/XNbcQYqp1xTM5ac1QhnzEjXHK/sbe10oXfnSjOcRe6Jcgy+RE1fkc+BlsRCtUpt0KTA/YR5UB
jUJd/FUfzx/nXhJvQz5cB6MRdr7OJ1mzlU+5fExsDNxZYt0SuVgNQ7qbAWsI5GkJOaky2CuMmVEq
iLmLzFChoSFPafwQ2ZUiKLEkrjZQzX21Iri+3pGB3s87UufaNl3tvOuvoKQGBAPE+vXxlG8DTYRP
fh706HNTCT0H4hkKg7OLPyL/OqdERl964RyL041YyMDjnjqY5OrWgW9PoH1jVlOw+gVZhMZKYFMG
ZerRo1z7IsooUvsoYlEAMQ/lmGkVICDG0j2N7xValPVwaYjcRyomVYrocAmdaeQWa0OHVKl5j0NA
DCgWV2jhTf0eQ+FDTkGC+mp3zuqzoL2HSJeR6KGMPy562WkIOH1rqdu/vZDoWGhmmOoePt51rnbu
qc4IDgHcR6cUbmJu2rNobt6jaSuOORW3MTjCBfmG3crkQJF/5/ig699f2N/BfjOfKPDzcCjF5+7N
Xhu1y0HPOAt+HiPKF4CWq+8QMQ4M3GWIFe1aTfmS7x8iTWfKpNAjDr7l9Uem/9/m/AX41PjbgU0N
6uDhxibI0cByUS/hrlVoTgTXgerfeXIhCY7fB/NsS51VGTM1koNHlMhWUaXyq4gik6zjH1ga0msY
Jvo2P+ZR9pshD+8OUFOb8jnLLOWogCKHpcHjI0vhCqdnCwfW7uGqPPBRrpfza3umvTI27VmjB5E4
n/sEPWXdDmkpUAeMzr4Ss+cZqoFVN6ecytzkVP31DmlVri8f79HYtFOf3eYc3PvsW037uBCBXiNh
2SHhmlkrKSzLvuhXZw0XGGkgeA1gcIQ0nrG99O+J0WuUttXUpkaqjAmExdNVTeIwAJKO7cresp2v
LpkGamwDbqS5yoMk3vXHyigJrdu39zlKElC3/h/T/ZNZ3W63MmsCpTE6Rn0lD9azLWP8O26sLfVV
gqhPUDefDd1o2hf5EiaYHWb1AVbB+MM2Yu/oydSoj/269p3R51v+g/IXw+6aF5hRWkHEllylbYu0
a90y7A1VhIEhHstUDx1kStfQT3A4VkXgPlIgmLlfwcjFJXAhOcrVOeDOVioW+3wzN2H4D9GWTbvB
Bz7rBf33DIX7IcvM0C9mNG9q9YFXJRR3pFNOtWdcweEOGkRrnfnw/S2W9KupLS8MtLfEEli/ZZiQ
jddeoJYb02HtvgrdVPIKotZ1vpcKUXxB8H84a1HCn6g81BUfAPbTdpExHQBVJyz7maRMQKbA9ZPl
NRc0DBBSSsIxJRnCkqKI8sqn/+TnP4iwToF8IcQigxJli+/m2Qe4HQLhGqc8yA+w2C/zEMFkEvyN
37xPqlkgNDVmiqVdSBmbzArrSnDY4oG3i1JvUXzPdnQ83IDPclSL5dchAIEgZ/gnolCz4JNHW8zS
kvQdnSNkv1n60xVBaOPLYSk3FcJQlAsfWxtWDpZhucwyw0JYb5wFFZ8VfMs2g74IBAM6fLwRX1Vn
7Wugve0tECTtREDOfGLKIh0KM8tcXqfef7m2Ob3fC3gGHRmnbdkEarRlfOcWyZc6kilOwygazUav
FFqKRlSHNvlJTzJ/e5ccRcWMCKtYuszPxsqKBPEifcFZKbeNXd/gN2lPszF4EFnWkIIlp1J/161V
AFi4rOtE4BnzlIT0I1RgX1CQuItWs2I+Hs7WoVKg19qVpeUbyi1c2PunYN0HYULTsUo/7bzJwRCA
js64uV0PJMqa9LyfE4QRJixKft4vCflThNmDQkkiqHGujBcbWICFx4/xla2c5Rh2ZTvFtVEiwaOJ
8fNnULJDMQdDoAWJyGFbEGOAHfUpCvCE9kdrJ3pRQj6Wbb5QV/7BSgDwV0IR1wZ1ndYMTnzEYnqf
p/OZMOJSGjkLUg0Z6at68UmKVLfG5kqCYa7NIVGXHvHoBQlqQ6tnTvDgwXLVYNEeKgN/smUpCsYE
TkQOG7cceOUzjOydqvXZo8CaNqgYuouX1oadqpZAMkLuRE65pRruv3KaTJpGFcKkD6ZCuKCKDmDx
MTUc7y76IYn17geEVG73Ok9oZJfeSyUsYNOPBsy9C3l54/aPDh5NV4BdoZg9p+hDrIaCToP/Ba4n
ABkAWsaHirpSv93IiXgbzfVGL4Jl77qtwk95uAarX4mY7RXD1Z8YNNPMFWNSapdCQa2Gem2mj8GL
KB5OZ6ucI+a6ZkwuwKzdyreSipAcGmkeJFqbpkF03TRV4QqvAP9forfDgM/teGK+I6d3STI4byrd
V2weOk/1xvV0jaq9In6F8+KFscKCnS7Ww8r7QEsKSvZorbEiUNtFFM9v0eWycFKSdt+YFbsQYDgR
fodP83RniLInscegqrNv7hAL6q7HoXwC5480cdNSRYDRsoFmbNWIulhK1OveVF0XvXobt+/ldJEs
r1hyQqNrhStmCFLSaoyMn05BveEaccfstjb4uUIHkkK3/MTr3Ug/QG6iiBg/MUarczmTTw3Y3Cua
wYIATSm02GzaSnftyO4EunFLv39YlT3ysFNhDfIJA2nPqyKqze4RxiFzQLTlC4pE511PRR3b6NG2
RYrowQmO90e++8n8s5Fd1mPrAPLp9+ELj/40tbH0O8mOi8Csu1tm7MykbL9KoCoVDRKWyGrPELvN
vT0xRPZaoWtZuPmGdUZUWqIRnMrCJVCdM9nwqrgNdVexIQG5Sa/vYLqdyicSOB6q0921Iuj4G/78
+IV8yYBx0l3Wd+Beb3HGO3cehthQd01So9VNzxWJcNRoQFmElceKTo8aiGys8weYl0P3MDyT4kTc
Y/MVoqQKgu6Puyh/YgiK6783xSqq7uaYASXxurLpFH+JBSUUt/P49iKFuYQE/9t9TbQYTZFrWQfv
Ia4FdnEiiPvrxm6j2cTV3RDVcyEvCrjRAl97dj3Dwfgm/Gux469A70tnK2uIeI3aBv0bEVANmCjH
FP7H/iwYOFLOruEgQVl64nlbAJn61hr/DsL6VlO54NbEpBd5Ei8GAjnFYqLV3prZYZdb+8pV838C
69pGwqJF21hX25ZKrqokP4xtrtKmJC6CA+1hSqJNfYSs72NiGHWEkZvYhMgoaQm90GmSB/eLCPMX
jjvy7h4B/MJT/sByqFze5GmRlfXbGRuzXb3HLbJAUdCn72Y07SGNamkGUotoI9oXkIGyz6f1Z5MQ
oO4uOkE5uC7fFo4A7UDCPcCesF4JGqn5oJkDCrapGnhdF/rbPg9rtQAeCnqCwWW20N/cSrMRKTx/
/nMGfT6TNCJyRFbxqa3jpme9zpX/g4cjrvchWEHtG2qiMmywb0A5wt3SHC7WxhzyQgs20gOgqRXU
fCaXTmpy/QW8ijECo2+ArWJJSKSyVxEF2Xp8YFkCs08vOgi19Xm0yCZKNckIgRBr2hi1qgrAPoQI
cMYHbCwx/BYvupYSNI0QFyzZQVKSuFdedTKvWNpPyl6ieT1c176zurEprut4H9nFHMl1yWNnQB4+
xi+rr1A1VhxsZjRm+iQ7351ll0vQIoXqF+SMJbwcbcv6y/VhwB7TcHoLyEnkOg97ZVsT194OewpT
2TIQWzr5K0PDH1sNOgoWRM6OMtiaPfTGdl5X7G0gB/HfcoH9JshW3YiVxkyYa5cbfmnYtB1iJcS/
icaCU+CfL/WtFpgIcIHpD2k+OIxd7xEll0pRm+FUO3hl7VrtnTn7tNCErnFtvR4hsdNUjOdjCeit
/Xx0dc6S1PUxggc02W81vyrzjc1VB7vRwZbhBBsHq3+CKw+pd13e44ccCXtDK63BMsgkRvNAEOlw
7GLYqgr4ZMex4i0sn/HVHJzszKXaxAu1FPrxIqm1/KgbTpQXzp1tQ2vjyVgiFEtRPfiVy4Cj2WY8
ERCIKADy90WA5Dzon+ebNT3mv9uWkw7Crpm9W9RAN4PUGrI9JQ03MEabbh1aZqnp8d1NltqPUROj
VSQ+E+3ppFI83NVR4l7IceBRX9EmjeXfdLP2lwt5OKBtz6+J0u6CHvtxXdauiPKSsr+rzGOwpAPS
9Hy2qFR9z/AVhn9CA1uF6/J1zaCYHJhRL7WzCAWrN4ixyoGjH6UI8OZ6Do/DRXsPbJJ/fzO1QcXH
dJduwg912wIzb2ztWeCLy/4t4I7Ca4vD5dHVrrQcymJ2IB3As64mNuCRLp3t4bfxdETnvvKzpLsb
A7XYUISu0J38gnT1Eb9IHM58+ZAs0TN9ESbyMJ/nCIf2qZqTre926sCLexwcRbVxug9ENhlm8gx/
o2928zKPvylhsA43Nz9MzpuOg9pGUDitlUgwk6k/1SZRUia2cxWYSaBb/3vG5OJjPc85A6+epnXi
G64c6NeTJzWHQP7NbzqLCr6/CXhWvXYlKQgIz6ZFgsVNmgyVB0nEozIv4//iG/0w9urrm+Gep2i6
m0bj3jbjHiSfU17G5c2DR9E60EtVIFpR6XhXjL4xXjqDPLJBdiaR/1+GbgBPVpIdFA/NUCg7ySeJ
fzKyKyercMndAqTBkQmT7VCsUS/hIQk1VpeGxmLPJ2Ld79NxMWzyVYcXHwCVZwxQ3hi5Vl4USeyQ
hvw94OucRktqk8htDiq8oVyPbW6oWjTu0sWbexk55+GY8Myxniy9CpuYPI4Iue0Y1OGQ/5CMCocR
OdvPM7RmH1AB4zUjC8AccHXtzh5now1f0yy64EEMNzhfywcRFrmGn8lQiRjt0jzUTmKFD80VGVow
wtEZL7LPrCXqvy2ElicsUnqx/VxOFz0eIHvoR+kS1Sn2baJnbGuDCjbb+Q/uGFOcwLO+9E1plEnL
sZEglQaoN6iTbHM2CWbhloFStc2BbqDhK1l9Ng1JEV+xShxbXO0MNiJH6mHqm2tZ3XYvjJ77Qyi6
Pd94iYM3pKGiydCZpAQLr2NR+v3ysL8x7VkMUZTxt519b3JtqHgjByY5KV51AKpz1es0EfIdNbQ1
qDzBk6GCF1EGsrEVNO396+p55TfSrHGYmbihHEvUiv8GMHRGhvm6914nVxlktk1qRDypnWNjls2I
IMR+Q/gaE1hJBdIkEZX7hLtOLl+ow1GwC4fLBYY+geN2KZEL5iuew1fAPlBaNhSYzinjloN+DRfa
ZmQFdtYfn32ZnCUXV936pMjBlft+1ILrGYKTUaKRvrPjOE0MfJdSrhnXgYfjuWgOVsTqPhP9JgnW
FI4lqmHxYJXgAwsBvS/6HLLZG/ZjIrNQ6j+PSRoXTLzbT9gP+aekWeFvsDFNofymn4tSaB/+hmy3
w889X7BINHs4gq6ZrK3X+t0eFFSoh27/xa4IvpNCfFhTcHTu//fX9vzfhRHJ+FEdgu8rD/VasD4n
c4x85UqA/Qa/S0KZ1x9h2bgZc7iEHtXCI94V9AxA4gRNBsYn2mkiJcx5l988qCCvfuf1tx+/gYDP
PwkJjg+mR+DNQCCTC2+hr/hKBxJdysdZmOW4H7d64h/6B/lYSEeDNTzr5lJrtPV9x1oJ7KNkKjSY
5K7GWmcysZeUD7PaoCB6xFytL5ZPL81QnW8ioT1xWf2nOpBPG3FH7vIXW2DMNIt5iPQa1jJO1jUC
E2mw/q/6oQIP2trEz4+TgCTzdZqu3SSeFDB7i21BxBYZqZOT5y7mua13Ypn61sX31FPOlwR8LlTU
iX8prAq4d2lsGgHp5Eo6QDnHPS4isXURkXFxpGxrxEJSMKtGCWBADllmirUNeZjHaT1flbwqPNox
vCT3pUWUlPPEXARZN6w4oZcoSNiHlhTTL5r0zRwpCVvgUFy79l3kWtbSskRiUWud5o+2pcUCT/w2
Il/fLvMLp4RlZnMviX3JI9Q0JZdcZgwpMJcaC1JHCe48X4cUL/Ose11sGekYQspePEDSmGXJ60IQ
x3gWOXnvUI9r+iUWn2jJG2mdjuK7UIDOdLrykt4TU0JtJuslA8EYtWTd8T4dSEAGG3UvEmVdOtGF
GAlFU2oozKd/77At7njsYeV19D723x1gbCYzM7sqJaPXewPxZTv54j0VpAPb2cjO+pITkwQ3zU2S
N10pxQwDHW/gW/Lw9GL0yDKU/7BPkkP0nc5CdkWr22E09wq1vWJpZCg5EXPHbVGb5B4TNGz4VIaq
90kc6DjEbhjKahbDyKUqsFMiBjGPckp0OLhKz0dDlxlzSqUldS4V8+9OiAqc7SoQY6bhsatOUT/8
UVStJ4EMFlpUvtzisNn9tWwlWAZuUYi1WrcJ9U12ubPthoHNR1FSCkzMUmwESIBsfV8tY2opvq0H
aEHHuIa8Tt517YEsvXT7AhyhzDTUV6qEv9yqGAzbRAAKQMLPJ4sl/OJUqER7K4aluPcCQUEfTrxb
fnPMqgpeLyBB+RRytF8oKICFXkX+1jfp1V7++cHURitbj0GACjxraHOxXU4YiLrSiHN3qkGhBdkJ
RkUN2O8uGDWv14f1pxeBHOxHqwf1YuVCQ5+GywARa4B7AepUpMsy7VB2riolKlGlMt/n9oqrlvrP
nr4Hfdv6idg11dYMLNQjZLNyX+15glLta9VKZFK0YqQwn8S4HShNuUlFpzQrOwIsDAN5sa2BRvqR
7jFc1a2SytbyHKRkd5i7vq2fgkpA3O1QMt33QzHT0IAEhNbNJVKVueUofjKc5aRewJv2OezgpaTe
AvtT6e4gpi3E+EqieeNcuic40LcWnBFYSWxP3Eu8sxvodX7ReQqtPeGjrMBQm9aEHbo9VQDyMN44
VSInyXI/ZJCaYrA5eDzZtywVFi4wNdlCAb+sPLTCM4fzQl4Kdmzikui7DNau4VsUD9SXgMkGKdaF
QKz+99S/x4octUqyDdZbk/f/p0vW+RBORItV+CGeBtzToOKw2FbDEF6SS5AD0OHM74o+ge1WnkQD
/94zPYy/JRQDFg+0odnsK6Z4+eoF17Wa7S2vHd8u1a0QmTbZ9HmEUQAHjYGIkUkPMcv9XwEZgJC+
GOcLGCKrPwF6XDJVpAXarmLa1znimniXQMukt00RUmw0MgBhICnVJQ7BorrATFIWjexYLtN9nKWO
nFLvafOHSmO42PY9kFRK4WRwBu8OFytLhst78LIU8i4Duh2oopvmdg1k/CaD4HI70k+tuGjyxSwA
6Jiojs+rMhWNYVgvPsIsAZgMt8vPZO1eiCAAzOlWKHHr6zz7Jh9ELDhiPgbpZviwI7J0dgc5NVuO
APIchV4BIQWV/qrHJKETLd1MhMlU19cP2RhmcBiNeY7dCfIeDXcsILIHu/AuKpi6WgHRtt5FZb24
sEQS7JDFS3t+5OAKkonBKuIg64tYHIesAkUr0PsforhnQq9aPWND4B/r69BL3b2Ee6kZbNjECMZS
gtUke7jTJvhEx+R/ByIvTDm2F/vFnJYCceiNGf4ar+Hc6G9qgV1O1Xagg+MG7IjygM+1VJC7HA3d
iViJ/vy9PoEaGbTDo+liBHg+nwcJu2xrShnbzgV48m+qaiWG75W/iwNr4mss32Y6MRE4LPs+B2Jq
qe8kEiOpfEAWw0t5AL6tYOMxZJIOwOkVBf0xv9s4vbnGieJ5Oa0DTqv9MPu3Le9+iG74SaYMzttG
7CHbaHa1TFG3tHQP0SbxJ8HZJZjio8wJks42JhtKsprBJbGZaxn2Iiw6JrgSsJ/m+Bhs1VUFhaGA
b/LEjZCEMeA2ElSKrskodzuSadsWE4wevo1INTQODEnDi4oWMA69REtmmFd1pB15baYxUWlNRspc
b+7GbPb5+WMfR8Nlh0sBix9LIh/tkApeiNYoCBJjtELosBOwGhmOo7x+NcQSjmLFwdQkIHMcQJlA
9DSBa3Hi5sCU0zzL/s4ApB64AlgmWibM/+659wajp/YBE5n7XL1hOmxEOIcEJhhnnDZ9yQ7ftFtI
aLgj4kERuYyzVhyQQkpHFe1Tdo2HyeqAU+8O80YkrEI2uni61PaVVVFwGxHBuas5hwdTCrbkwt4b
f/3Ld7yqCy6CVV9O7C80jIsZakxrYtTXsGTd8PvXE44+FM4UMnKiKX70hcQZT191rVk7KZHVQ9qc
cnlYXS5mYFPdwOSbzYQWc3a5LvFkthrX7QpBjl8brW78RY/T/gozK8BXU2ZbjWqlqS/vXa75t/3c
ia+EXKBR96qznFsD9t/j46vwm0L97zIoRRM10ueYmRoJqVA554e6hc25R9QwJQElp+eD3jcATrLJ
fOeNmntiqaK1Wdz03KRuGmoVPGQYy2+ZyqYg5SBcmZsl8U0hrc4rtR+41kdjuTd7KX4Hj6e8AVZT
GLyOULasyFqXsgRx7Plz9WGns/yyOw3zvY6O5A6xyr4usZpA/03qQTQ73AOGI1/2W2D6QfELwQSY
Jd4Ke5AuVvbI+VuHsxMmSuXj8CbRAzsayLx2Fmg7RiNO55j/7GYi6HLYAKUMGZPTx8dofQijyW3F
cB+EcWPUGbKWZ2hJDHaQJ2APCO6Zab3bWqudfFK6F/HLPYfUaP6wNwfRkTjlNvTcmtn3YG3m1pBd
bLvA471t7Sye54EDaxMzodkmUHcUtTCgTarMf8GWQOFn334pIVcK7yqG1k1ujUCDkBqsLnyu53iv
cuaykb4FKna5L6VYqKvi9B2xNy6dh2if1r2rqGUri590fUVGlPT0jcKVl73dxVyep2j3Lh9va9Uq
Mi5iUMTgRhwjfKiINjtj9oA/hjZgidRVO0j+emOUsZqfp5FnxQW8tD0ltCwBujaJzO4DLMUsBiDp
7WTqZC/RzznqZ7sfiQ6E78DHpzR/BFB4GmEf0U97gbyu0xIdhFDIvTNRcmHcsp1KMz0lvNr9x2xU
c/tnLA0C2sRKY9i6yHRAIM7Egof9q84tUDQ/JTd4KGVUwKpeDuN/a3AHcOVfn6N+eGy9PcwTXOa8
mMnl6FcRfppl/acNDrWiZH3Bujc1Sm5BP5DORflagpo8WWdaEAYQb1xiHy9PR3+wAKJd6Y40/DKp
wCWXnx/7lqEet2kRWm0gufkH4p02QbyTkzm4/DJi0B/DAVehdeWp1KIHjX142bg3nWN9F+4DC+OM
alIQyXuWLUfpln+WLnLLiIevMQmUH94i1GNnc32xMsEx26pCJ4xa9lqx6CvNvO69AMWKRgGGZ75H
C/1I+t3dF7c0V/a2GJULn7n32bDjHoko1tb2jiIdRhaIK8Hehv9p58QjSiLfN+LNuvtuZXe4s4Pg
zwKvliwMXslLmqKbnsDaX4PXhMgwc2CIiB+uekQUjX/OCOlQoja1PiFfDistS1JNk864yomF08Ss
xOUhMqYlHUho19HNMoWQ4wFliOYlqUQlg/W5JlVm1CeCuRTirWzNlnz+sy8Hwv+zOCnUVrXhP0rS
+y8DqeLkkKKtQ4/CvOA3ZGhmDVBxEOBe3qBNfep9MCKQkUgGbWiRWMebrmRESY0Mz/aW9VXtmbVK
s0VH+bzLkD8N6aCtvzK5TlzyttEMx1omaVkm0XhVi0QVkgsgoUQG0ujrBt4pjTtUxttR2gknOvYv
JIoDtCE8JUA2qxhhSLNN9o3dIvPo/1WRjEjK7SpqWF1FLQDNTsrnx7smFstfWbj8qzVmPf4jaVJe
8EsLd5y24rP8RvYosvVmjbBtZgQzQD2ZeUquEq37OxOTQgWfgpLYigOct0hIuHjhUPL8SHXdaqiV
IIDdoFfNQ1v29zmwhpyTzMTObu91fOrD2RQf+QQhjzf573vNafcGKiofENbwG7BuQVT5g+aPLFgk
HGcQld/z/3aP5w48LiqSDfAwAir8XZw8Rr0Jd8SgHh7xzr2U4HGpuKLbpML/DkuV83rwZpqp1m7r
rFth7MjCPsmLsVffQC8R1XWO1BhMgXKmsDEj0DfxogEKnn0X77Ds8mZTkG9aHsRKnYlxEYndn/qV
l/BlhWiUR+6SK34RZyLvV/2I3bLtISdys5fstLLYUNzeuC+7A7HAdHROCW1HcvVGvD45493jIzM/
du+oDaHGAZWrGYiMN+YLaZ2wIeNSmBkZTViI9+GR6A34BaveFOZo7qrh9CVbKZRhZ3DKY0jjhNd9
Hn+psizecSa+INN/6cJ+DG/K+Dlvlrr2985vJqWGLIFZhy5rS0X0nRWFup1XIlfOTfETuKFm5Vwt
cyybyyztzrGyWWJ4vnZosB8Q7CNxDXcEL5rhtH91183qAuu2BHT5GhwSpa33eI27Wcq7UdYTgYll
zqK/fl//f6M5XG4lrGgqXCrvDEnqHIMdj7jUbuBvkODvuZTKcA3OlKdUFjJlfr6KGmOMyJ8rDPRK
mZXZDpIJfBGqgGpr7pjqAMhOq9pfrBB4bl0ocgUuQJImunABO4P+izSmtEf90ubMxdJfrFlKgWq7
bXAxfM+e78RlEr4RadRF/8sndLZzobN4WkLoKRABE2le3TZ1mpXEJMVGN1rZysN2qBq/eyDYzfKF
xi3IDLPn3b5Hza9QjwFrZ9aSzHxgvpiT7ILNDq2A6r51EIP691BWLEdi/QnIf+dcgItjS4vyrEk5
jJd8ykQHbO2NYFZq7zfZ9dl99vD7LNz3Q13X6Dx+giDzO7uklUrvX0p0egsA1km1wvFmiMKtbR7w
olj69wBYaHiw9lDEKnBZexsHsfxvAaFxzEXt3tvNK6ZSPdrU0Eumn5d4XIJH4g+TcRDzHvtH9RS/
7ILwwbjio31GuTYU7djXee8eRPSrTuzFOa6tH0cmVmwlIrLeQQOBEsWxeup4zaFiQ/t1Sqrb5rGo
nXF87eCjC690TfD4K9r2quzI1xzfpaWjcAosIA6CHUOr7xVc7SexVXWwCiLzPurnfhGotjqYuUKM
jMO3fJkiw4/XeuBDGdtA0QqnRmond6LYY8PPaudRgvDcOW2oE0U/1DyJrAB2+G9yRWwn4X8jW9Yz
g15DxCmPHD+NX39UOQmR+OtuGyjnIMiP5mqpgrnJdxDLNigd/GAjU1mmxm77VGJAH3DjZ4+XHU2k
N20Gw1VmZjBZotwBwjZyDkQdYW250nk1oUKdRMyl5hd/CA3ogVZp7NWb+OlDMHEx+G9ZDxgWGaXC
1MPLqFhTMi+qBQZZGMIEC4JZRXZ+BwuxhrxMyDC6TlFqRo6pomuMj5suUaCZTrT2/ATgO2SPJLi4
OD254qYsaMqBuqw9XOkmIfpi7sjRkmW/XLycmuKSdJnrB2smRIik1uTHPl3R9wlu8j7Tkurnglxb
8/HGqBZLuAsmyzeErlVVtwwoU4nelO9nLHtlZWFRtBZBGJ9y4YS4LkwPdwrLzh7JC6zeHQcQTG8f
Me3opMxpXBKZcoVz7sRPfEkSZ3WzUt3A89KKkbzpfnFZ6yuL09b47Ja5Qk/YvYC0dWhEtbkOxsPW
/GFquVafV23ZbLWGacNix6A0HLxFasLgTsJ57WiCi9SNEPVpp9DX+kHZekEMs9w9sH9toel8x/t4
Lf7rCE2oP+f5iDdwgLszgoEQZLU76QeCCcKWXdiHinuo3uV5kkcYy3PPqHbtBZujJd4gMPmli5Kp
GMiPQ5FBa4MlKFqEN/sbov9wMIoVV4oSiywmlVWz75gYDY5zK2CbWc63EwbjPe3dyJRPDOkU+2eA
0/2t1hwEgdK3BG7k27COX5/vKqmSBada+RsF3DsY/NXIKBWDill8VPi4xsAHrWTTNHW49FpKWVi/
XSdZuIGUOlmMbopTlDbN4Ee/YCxdPC65VEJ6d6sVsCsPsIqclc1rVxDDpdHZ6h+vU4K9gQXOirvm
9E0/Yf/c363XcjYylQ5t1UBIBRHTBv+cBgjhobo/C0Ww+TpCNK7Nf7TDXC2Uru8nlPGQHWdeWwxN
0IQl9I9xL1XP/l0d3puoIuvjJZoA9gMM0n4MwmWNqkjBuiIeKPcDJijh0asYyM92fjLh8x7hPuBs
MFcotkmMbsX9M+JCTdl/+gLj5TOpIUxXVge/Y1O9ArqG3XB9skGNV3xirVMIuTiw6wBn+91VeecW
WJqzfEYZv8M96Ie/xcxuR8jsIrXTXLKmQI4K97vVHK8wWz6hueTd4nxtpS+St43ufWjA//rYbuRY
4dO7Y3T8Y0R2eDZqXtFyMPhkt0vrs0BnNtBbSYF/8dCYAfeHYcGB4eq6mMXDJzfvZzqLsKnKyOaK
qXwUobQz3ORQVk3SPJVXO8je92RVYDArm2dWI9rGKrdnPZXcIHQCM7PkY0oQcwu6scDs7v7XSX50
ygoRJR3xB1JIVdvxjCE9Ef7JrbdNfbxNBQHiJVzQ+t4SuxhVypA4igTeTYQjxY/UNlMG7pQY80FO
L1v5fOE2GpNxM4vE9kDRjdX5stPqoFzorYI/Tt6CRLRhhlGBAz5JTOfFEGxufNfc/c/03ue8StvA
YBtlkNpvWlcE/bRch/YgAZffFHf/eXXniFSDW5ojsGS6bnf0lEsnMYmq0q8RHSisKby/Ua9Ok47e
Ez8Smi97ZlsQmlEshx52NQDgGc0dxRGZ6Kbx3CSlLZDoAVpmg2XPpHAK7vGef2WdhPY3U0ad/gmR
7eDZZbKU2ZRhAQY5lpa5zJ0PJ7xfH7GkJcAnlFTl+vLwvyf1TD2B5HZP1dijvlqO2esPioZLGRc6
V2Va5EFN4MqS4+eV+fgT5BWkNBkupY9awgKaoE/R53XrmQBzEeLIOYqQ7OakPDiP3xBUwUPKhyfQ
N8gsSt58OhVPX4LSLo1gifLuMprHv4fyWwB8wPQCNRmUXv3UaynF6jCO9rXdvG1CmlwXeevSM78B
G47HDHPi8qP28xUAP6TA89FrKbvcJ2EVwDa4PPU0+L2CXHhhctCAwNwuD4XRPC+rifflGf5XhWpb
YK4Jo2iNrZguNGQqI1IyN2AiZeioPBW2ZCGDRZOW/Jmk18+gsQ29crNOZBwv31oyN1rtdpySbOst
QG3Ig21hmBBG2CfG90Mv2cVAE+Wg6sKQsh2ZrRUBLclbcI5bP02vdBlkMZeTwVE20U6v/QFtIW+8
Im99FHQLDgKyPEv+LoxeVSZK/n8NKM7EzLaFfc4Jxo5OsXGluRcrl4vzqsF9wy4R0VR5V5OVIv4i
20LASjfoONXz6teKlr8BBM4PEIrysSZdrPb8NGtUFqGmC2DdIICt1vYdKtrNs9bp4Hiucx8zCNtg
x/f6qQZXGyZxlD2KTgRtwW30pNgk381xuDUjjUAov0y+37OkoDEDNu4bQkD+dL/8uFDtpCZsksu5
bnzoxWL7/KuRLb8hL8YBS5rNjU7TGJvCkaYGulgXhlkndR1/HVHQWrKonbJLgcuEfbhd32yGYr7Q
wLvyWaOkhb3Avp5fFFOTK2FmKw3hfqL+UB2bH6XNpHbRA/1HuIVTN8afLUhfcqQAZmiqHWQ8Ot5Q
jjuMDrcDmqQI2QhdlTYvrKKHFcC16rN6v/hKasKUTK1WGs7XjqZDMRRUDs0nUMNbzezsTL7/1KM/
YRQfbjtSVT8BI75FP6FUElgpjjkIazTMaY+d9nVFdtWKt6eNEaXVa93TtDkFMsbGmTAUvaDlempu
JiahWqGQRHAoICn9ultyaqlnVtOgpkmF0sh0dbrHkpAb5aVmcitmsap0C1qAYZl+KZXofWKTHWiS
MTQU3EuP6gLIJWwNaJ5fy8KnWpL4couhso7DKUSaFopWrVO5sTpdtFvMcrLQwK/U8m/PUV+uBBYy
Sf8sIJlbV+PbYaHBl/BxqAo+HG38wgli2Ke3mV+jy4yvFb9coJqkwJXOFUQhNBKjjgXPjnSl6E9n
tfTQzMZ9FvomXZ3cU4AFBeWIrP5oe6g9Ub4NKE7rFQFHQmQsjalgAE91dBJNe0SdUw5ArF5YPxxB
/e41fuwA5EmD647B4SkeASLWyBruLBVRRXYchZmdpsaC1WyLc6MtJ3ZTCYEk3JxeJH6fXzZub9Ua
ZWWq7E5kW0v3fKE+xUUzQrNPsm6RHrVu+vlnYa9lslxoJRG63GzKF22lNqAsYSe02PQD39bNDExr
OCkW5pI5/Mt4Azdwlszvlh+qBXNwgFqeEYq20zqMA6RUlM667nHP0T7zxLo2kTo8QBCJL/wSvA5P
cPkZOtUeiF5fMvv2GxytlNLOU1jWqrho5CtpD24uzBVL80sS6F4dIWlCHjzDgTxIYvV9Mg3D/Flr
3bkrVvRo2v3ooHbUzK1oq7IdxYn5FYzT+B3XUUuJcfrxvNFCKCYrstLt554l8t015a30qlxev/M/
DbCZ6aaioAdktp/xF0QUfEaFrRwrgdiVzHvSeJLjBUtNqLjbF0WgEawRg/2Hrm9K0qloF3k4uaLu
qWcnx/jo9JxYsHTPCvKJYMjotFkarZXvJLvjYZRkNiqGDz2D+uA4OlOjvu/5G3h9NCfcW5ofHqX3
5VEw0sW8ylWBr2dsUZ2NrxX6+fYGOVFa7EO3QzNzmbmvsHhBYW485yEMa/eu6QG6rxO+BI833swu
rFP5oljZZRMTRjnc3MrPRt1qk35BmkAts39FRsnWcT0rMGAH97s+JgigRu6BjTf5F3TEnl5X+COF
JhdusGp+55OT23pBfl+sMKkecJ5mhURi06BKQkB94+V64kOulKTYJbyF3PX7ikP2rrH63g3IU6Eg
ZUp//JpFil3AEOXHzrElzXCHNuFdBKKs74hC81ZaPUXrzrPBsvEKoFxBvG4Achjfwhq1zz+/CQga
WrrN4ohg/d3lhE9c3FCE3X0ZDeV/BG4Khl7eZzq4h6zISzLiSyZK2J+u/bM+uH5Gf4ooX9wfc9Ix
pwH052AodHuTZ/JPkXnCAmiOw0Gzl52MZYq7IU9ZMbYRn5KJptYpjpVxyViwrQmSEW41upZ/MeSB
1Uw/KMKarfZh9UqdBJxr9sE8SCUSxYMG2fSiH4Vbccuxc5RV0b7xnGV3i9U8zwe+ugtCrWJMSoKf
0v61LozqLz29g7BCE7XjcsMVWPufD73FOQtSBEW3Fo8MM++8gCEUDcvKaCIq7byHsikyIh30Nbpu
YaOjuoP4oYVIQxXW6tEmebOrDpPp//CzMmgOXRmMN1XgIYtltmAYg2GVSS+cOfn5Sw5K17hu8JSV
Mls8OBkxUD4TR5PldI+rgahOqm2jiWiZ/K/klAXte17uU3DzZRbvxcHgEbS56+A36vQn0RUFUWm9
t6zJsRdAis/+cRaN7DzVDqLPEFGwGEWfb1sgTB/dIOiUddDOoEPj7lJChq/RD8LTwd8QgLTDzLFC
0OKzbU8PQrJnSdBn4uqNzHsh1bpl6HLeKoXdT/3q416gnmnOV/DrWXKP31xGVBXsBW2sPIXjS7/O
zP7HblKXERljBwscOtlwqcFTHedBrP3R/vZ0Ew3HwpP5jVL8habMYfRPvuCVxchrCRA/kodp3kU3
61Al2Wikoy2RbuTfhODP0l2S6MmClamPFGnT1DdgkNWRzQYJ6PGG0F3UaiGJ1lqZK8WIcC9q0AQH
5B2B533pDIZTIcKiRQgwfzxldJzTuYaVI9WY5vbkNDnEihht51X3sdWgftF0jvJNM/Z7VvF7Ch5O
hy6w94b4sF9xGUmr900r5C3NV0XhQ0DJjYAEsGpTRf9KpHJalMcMXJ2FEocbo76Gy32y2qOOmutS
a71t1jCLPvSN7+SeDLyFOd5fM7sgzdizH4Dd29ZZ+C0XUjNcVxssn5ANrcn3S0PTLBpSkCLXhf+5
AVjnQe0NIS4HxbUPIKTpQc13WG6J5DsaWEkTdxsm20N3PP6mLOFNozQzsFzdvk0w6raqAR+AwnUj
At7u2pg/ReR11rwYTD7P0EBQLVZHeDKM7gHScCdOcrH88eM7BzEuOPbgFsiEb1EXvW6KIdtSP+6f
4rThwaOlY5fH/I9Wh4OEI+2FENRUZrbBE+OfdQGiUuPqmfV5SxgQxmStBi0q0JDgOwJ0iU7AnkrJ
o42kOYKNLpMttLa9wNWS9OEeyAYw4qXtuefpAhkWS3gev8ds/o37ljLsQKFS+YzNfxkX3X6ptsm2
SqmFOLQY2yZ1HYcUeFHXrENowxdtuuYneB1Tx89Z2U92iOS14fdlDuijkN08csx2qJVVYAX3UXS4
Pvrwm+w6oO3yJXqtvNBN9z455w9jy7h3nr9LIhLiNtoXc6/jTkjBWS1f9WUwJ3m2J7H8EvWfFqfU
ODKRMsMKO/MxIT+hIFxkeINGNf/WruZCtH2bwg/CA4SKUrgXiPl4dui506JFIQkH3L8cruubI7Zf
HaK7GCDZCYyLQyu4menNURqg2A+ybWb9rp+/WOIU93wJ0MDB4FgOamqQt2r+Pd664vnouJVoSUyG
lpxC7DYFnnznsEcGupBZPlhkvntizM+sVcYv/Lb0UWrhNI7OXPSeCWr7ZGhv5dphK5QEtFMhEc2J
qVcK4PACVNpd9VFQHK2OFDmO0jEsYiGUY9sMSRvjTBiBS6dot/4wHwEk6K7kzzVaK8VFNw4S7Kl1
zj6OId5Hm9h4OnOMEw7RIbYqLTQzjJQO/Yet/Q/KhuIPf9YrQIipJdh4NuMIAMa6dimG/mrSs1yQ
JAWJ6oaP5Zc4KK9nIxkJ0AALTGqnlFuit0g2bW1atrmGN2soC2qxZXr2Fnvv/ZiP4t35zD0u/zhr
SuGkGJy2lWIS5S5wCIHRXCLdQKAgUmKQ1Oqev/30noPR1zPldyl2uTm6ILz58GHIg7cbcU3+weXE
sntrrIF5g3jLYEi2esA5nQp41ToM9CpxoovtDpTjTEINP2mRhGQ5xeEXJzexx2ARWR/BD1nvdp8f
kIG922bpPDlNLCxQcfGf+OSwgQftWW/oqQbs2vaJnKP0KPUYsR9/GU2AxhdJPbzGPfXkNOukMcYQ
iu1MN4cBwsyU4MiKdibLrCIedcsCcyZfaq9Ef2YYV3J/0eGy3wem7UpucnL6ikpfk4opYaZA8co7
acTjwfnuLsbSEVw420Ly1/3qcbnwsdFzbt5xYwoS24QnY4QaCthEoiLdWoBYN7GnoNQkJWHyJ+fV
tUeLn9yxk9/I/OaIMH7+5LzJ/y5nS4aGqo8PIrDEDoo/wwcGzUg6e64JaVZJHFggviOgf5hlmjFr
oAfO6YkIPBdfNk5LYBzWcljl30cQBp6JJiDn/jMV1PPDjQasj1o268C5h1CzFyYm5mPLsDpWsfl4
gD9Qi3GQPysxwNLDZZiTU7kr8I5Lgq09DWPh8yDzu47N1vJ0BE0dYI1aqD9FCytNSFF4vskI4Q3Z
lPRp+yCUdpt4Ony0MOY52c4vzKuUQBVyNcNsSYa/bCRFD4a/GECglQOK/kRS822nSnrzbbPwYGRP
sxO2OoXNZ9RurLRPMJyd873QkmYnGf3tsH6jxSzboK87HWpl8zTlWuCD+6IWr+1cY9NGwhGNXWrG
lVtNiALYB5ShJC4W4ZlaMaRhOxBjaGP2WYPpWTsspwogYGCxMZpC3CZSJswm/fuIsfkXASw7vE+x
Q0mQfdRnTs8gS7XSECGyVIF64NGPQEqLX0ErXDMoCi+sbA9oTWZoBa5jcb7/gW1tU/iCBWQEGRnZ
kZVk3KOxzUucYB8pLKb9vBxTcFrKM15z6uavczCWs2gAdkwBJBeN8ocawca/tsGMFFU0l6CzjLco
5NVRVNI1qwISc4yF7wXtAeRRxddtXJMz0304+Ri3hsnYOGi0sG4fzE7t+CjWuABfEBeHpLxxOXLE
/h7u9N0BRDBh1HVCo7Wkhl7hCJrboc2RGoWNrasuE3CDoIT88FKO3am+2IuLwaBAqrJ3OnR09DUj
GxK7lNpOdQNsArD89pR2v4Ek+pkFJ/mA6xzERV47LowYO9iKGGt1+UqFKMftp13chMo6jmUVxCZP
Xn1VdsdVLRWMuYSQsASlnFYGF1cz2vxwKhqIVWyZA0ltG460IVbeCwmvD+VCCoquTH7sHDWJnjzf
iaXY7D9vqBbK32IpbutwcJ9JQtMFPgooF1vWg1QXv3GYDUzuWwXftj1DxMc+Aeway+ZGn3ALmX0J
3Lf6pAKygejN0ik8wCYqfigFJuZgIgPlVTuKkWXX22XhSronrSFMGzAgTQEDF0AowMzQ338/N4Nk
HK82auI2+o2Vz0411qxCC/6V9tvUzJjHm90a6oeScI+ssN1kskJspW+3q5RpbPBlixGa8WAAztHi
lk/+MljFp+g4/9xj8uJ0ErT6hCHEhlOs6vwyNVEIB9Tl/xTVP1Gn2DxkQFutsnPxmWtZ6SyNBy62
FMrj7F1xfnCkSkAQ/3a7MIbRhgyuAhBr3pN/qyOjbTRFp21d7IIyYCNXGArQx3SfKMSv9MF5yMrs
74bcPBCCilSD1ySuxEU8DmMSJRSsGnGphGBoV7Q1c70j6sQAaVXu29dQbbXQQ0asBHetO/m1Nj22
me5cWW03T4LM0bgWuf6p0Wv8NAXRwzuui++07wn8HCmYkhaE+bZNFEZxQ0TH5c7SRYfgVn+mMFEY
4Sw+irAVXI0uSgtjTBOnTKHgHtlx/lHBLPyNw6ZDWw3r/YAGGJ+EOK+AYba4eq0EKvl/5w9w1GjI
9csVij44pDIXgUfYDXUcbhjpo4gKcq/xtS+UUlYtpGiJ45aqOjy/F8K9hlksNH27Djc7yRGExCLF
pACpQs8S0yN7mT78D03edCflkbyUHLSBjI2qYJZBvNlaIUuQ+p5on+3zrEy6SRiAhLikkHkkF9dF
TMdOaKhyaoKRVa81Dg6G08PSf2r8pjvmZjpsa9e45mwAzIdRUw920PThI5hnIqiAGjn1HAErPFqx
JDW3kNLeUSlrd7snl0L2qU0oGgKbw+Tu+/8ssZXhu+HFpUP3pr0zN72IOF12OGmp/Wg9/6UGH2z3
QyI5bEYZdetejnqGf816K2eOcJH3csRJnbu/gMHjxol1yyOfHrxA3jclyDJ1uIk/SyXvqkic2x+a
3MPDCMHyRp7ej4pJOAZVmBcGGh0zBANzxZmREMUVMjXtAgVUDM0gyLbsg37vJEfXm3ybDHDa96S9
hf6OF4lLnoW0DjdJ9Tn0nscsK4tk2db8iwNqoHHFDdPIEXo7/t3H6xJVlw6g5OFkQBBO2i+SwGHX
Iy1m+F8+sIVVHR5s0g7EvRpXrj65RyBDKjxk/KaKXCcOz/SFWFO4dgnz/PkoO6P33E8sVk13H+gZ
hb/C2wuUnFu6FzYxdQO7KYru9Xh46tHLjQIg7PPdkAsO9MJHS0SL59o4FTnt3QCWBv8sTK7GM2YX
DBadj4m/Q3naPPHcx8FbCxIyVVThGpyAzu4shmzk79DxIDINtwhxTg+HNPJvFtS4kwY3OpM6Xlxo
6NqdZzKP4Wwu3FyeBSeHII6Nvcu7dgN2v/8/6GHxHXRanLlTGwmYc6Gn4n7DcfKkRu4HtgsaKyFC
q4tQlPfATWD6/5k7jF9F31R/yIvNMWgYTp9DIotIWIs+7w6SPCkoJ91tAl1kDx/58QW9TDotcuay
IWqeeZKYBTdUw1LQNFLOo7ft2uaN7npB/6qGbgnl6C7HL6gIV5eDgDS00XVwvOiV1Fj7iOU5pb3x
C9/0hS3nuN/XIPLRjfVjFqlxC9GhSeW7mymu+EVN4zKpmXe/rLEHm0HKA2Z/GN1E5nyz3b6iv7K8
s5TFVf3mtILr3pcdRXFye+Zv2XwUsjCIRikq1ZjCx0XbkJvQXXvwDoPbLXduW+nDzC0urEVqq1Pg
bQ1UypNWxwYsmVPIwBY3DsxS9qYoIoQkkkMw5IAkKAm4ZJYWbHEnUnsaVPgxivbqi+htHXsXWDa9
Sqg6/j78UIRaw/8jx9vmpEaEJnoxOyrYFLM0dVEOMGdPp05rYIGV+8+rQkI4v8c8Q74mOkR9tkzI
iuGJgT6+NsaV99Y38tkwMaHBH8wOD+AVBZXlWMgjUYx7D+fVpbR6cSFE8V5NXcX4c1i5ZvbODoRM
6ERMMhKOCPpQob0lF89RMDvmtIOOQH2VoJhueAtJveJldVybX/sqGQI2bZVfuxRy81LLXSz11owS
Cq/ve4f/Tg4dmTXLqwmC+u76QXVseY9Z6aPFvsa9RksJTS/H+qprXKmp4SIznyafEH+grUydcfAq
uYsaK9vsusxBLxaTx1TYD3aRbSv58rmfQlj85o6jSAUobTP/E/mgV1ABXfHpdHXFPYBLr9Yz1WGB
CgLupfmg6+GZD/p6BOQaX9PQrJd+GMtm7iFhI8mxqCWnrX3hv6FPkhlYMNjczH4DT2BkRK1s/1LI
xQCiApzIMZ0ySiUa1+mkSv/pICJQWXlkYJW1tm5tNKcDx5H4N+pr5/lQRbV2Itl0WI5fNadPc4AG
HUCKOtW6qjmsR2ZM3ElCqkvVPOUa5CX6B4kJ1/y4NyIyw8ZuQbS0yCBUqs2mbFybOPbW78EM+MxG
J7ObMfiMqBJRZbA3gRESA4d4MRo/+i6+7nyaeJ8ApJjOqzXkotmFHt1MgFvFBkQXCnJjxkitr/YK
ucIF9l6Rd8baOyXaaMlea46UkOp5QluYOCqsntumFo+xfoj+Wx8T5AO4ayZ2cL/b5F25k9G18uNO
NEdfPp3ozdy7pfrYW7QrRneCXGBgt5HtIRw8WwPyFR4U/MJPUQ+fvGhejjPYunVZknHv9eg+yWW8
RSBrHpxbea97sh5Y6KukX7ZmGDdd4ogs/dsioeu7iwz7nK88SwwAG07/5zO6YQTe94qTCRBI/hKX
5ae2kYIEkqdqUTG1ziKgGtNSuFBNLxXcRpfmpfbHomeQh0DLLLVey9u7Rq0TdH1cRotQM5IJNgJ8
s3HQ3PrKLWwcItHVPexB4Lc1/Zslc8lWteteCmPmuWlVrCi47qstiNV7cvARyFdnSFMdJNtWlJ4D
Di/zWkTVOBlIQ/surEqBBnOMcUA01mpKKeoK7tZX176TdIWYPQ2HsoE3ilqmbkiuMm2ijDv0uVGp
xm9dqBeNKdnloRNLt70IjDR4nIqGfF9TnDF/OKYNSVhwUZIUINAjT07GCGKx6ZRtXZu45RDa8olI
t/zKmpeX5AexKdAgJoEaptlNXbUYZYmHycvQGR3PLtG1la3ZrMc/p3FF/PUCd++8ss14Ae0wRRZ/
IZTmveYCaPNmb8YMHVmbcbO1ys+ZJXpPJ25hyliAsi11FW7tc4inMcNXvysc8FbNT5FCXynv2YJ4
1Iv3pCQVXAHPmRgxTSM7yf5ycv5sEAUkbpuCGSSAnKSkv8pzwCoiQSjdUfHeGb2rdgAZ8KyADyl+
wWaJaCl0ARJ08yFMlHXQmHkQ3p6UqLIM+bLcL3AkBtSkgs4Epgp04oTrwzWUHtObcn1XytR09OB1
V8l7ke2Je5/vdEN9KrzKHPyYgyyfjnjT0D/ngnl39/TCjtI3JxDi890J33+gAnPM4ARpBxfrEJDS
GqB1qESsGjTKYs6xSBygI6P+OTI/VWzjHaGeuMz0rCO1Ke8Ox/xka5ir5QM+I6QU30VxIgETc9fo
GTTtSVaxR57+ae4mIOpn9L9CYDobG7tSYqICIyyTb2T34L0nzwnaUXeuC9GnHLBGSMCu9ym6E8ow
/RKV8nI3QSVgdJNvPQn3a6n2u3G9rl5vLb1edQ6nLllhtL/lA7WVt+uiuAG/9RmXrKAVBJWKIA9K
FaOJ3gDJOUN1CHuoiZC9kdYOtknT2uF5bXWymILILpUyEWH5WGho8QV28qeeSfhxX+VQNNSojyrj
+2aylAarbVZZBhOqEqQdh+clSxPzsZytV2yDcxm2r3LlN+zg27E6iVKUC6l/WMhRNBfRibSgmuSN
v9HSaIfExUR5BkL2wtcXLnyrqlK7AekKtrC3lpmHQbkqmJ4mY/PRiFpmwICEqklmZRt/+52M3HAh
4seA9p39SH8BoxHtXpOWZIPNEhtnQy0aI8tyq41e4WfcFXBREPDeJEgefXRvwDMLhkPBM/GA8QkC
+R2fxRQK1iOm/ESjH13EqU3FHQFqHP/wwdg4+UZkA5QUAzJKDnn2fo2qV7s+JdzytwJxqWXMAAsh
oacBc0FGW0JE9O2NJePv7B+zN7yNcfiHVwe4+YI9YqughjMpl58ov6YcSBunMqJQwQpwFAG2wEvD
pOCy2iI3n8FqmJoKFm4mT3aYYv+kuk7jgp58u8PLHRyvMJgNk3SMjBvpMSjs8c5FoeFxuMz8xkck
Py5GEdbprt30icq47kbxX3vgJBejn8XuNaH11ICHWD5TWYfRMsaqEavm9IUmOy7ozCXB/RNz+0tX
HXwhSqf/A0kniGYXqSv5kNhX7GeDKCEARPFNh84ZXeHFPHB4t6IFsO+lZRIQiT6eiNTd0QGYcv4N
FNHWv1jfFjSBWEn2iECkPc56wtKEz0dXx2EUPgo+l1R1eiNit/bW/8QgLJG+Vaec2VzxvEtQuHfn
jDNz0QL42bIuBaSM/L+4ZV3dSwWyjQQxeFoU7GIWk6tJw7WlI20cq9aZvvHCfzS0y+N79sLAtt+M
So2WDfY5wJbX++/XsGXxsJTXuoxETeUscoGgY5BmIjc0DH7o8hkWi36r7zRcanI4XfNzjsSN9iVL
TFr1fYnoGHGmsm/CMWjen/nkpEsubIMc8uiopns7p8u0CsB3vN3szN8xwdh6Y3sE2ibprQVPpbrF
x1joy3Fr5TfKGoV67HcGjiCboT9DdxGCZf2uj4TrHrypXl8PYozlaUeqor2F3G/7zzro5FJXpQPv
4Sj5LmJzsCX3ofqtTzIZu4a8EiJzW+22jNzPPZMp0aa8iRN2QHlc5oXpkpzfSINv2zH5tR0h5a9U
1K8goeaKHrTvy6WI0kPT3Zij+7vLeUHhQFqVfm3/aRCTks/qxPhJb3d/jarsxb6n3IVaaT3aEQTa
8vWcOH/pkGGiQoWZSnlUojZjOyX16Y4sP+4UIGDdponSAPaJtJluOJGgvTmFYL5N/8G6dXMqvEgu
mJYrN4yXlZpFdRQFAOBpYwpFB35DPc8FeBoI1z9E7+Edd4e2Yyv9VjeT5VVussCpRv1O8FblI7yz
/vCq4aMGxaiARc3CA2icMGkUSeGAgivS7ux5N6KPdyeif7ObcWV5gaKoJJGpBCBL80Y7DpHuK9dr
6zDeAJ5w4e2X4oDX4S4sC/wnFQkXTtmd4pcDc4FrSzmpGHOTkx3IDtRxyyYanzMgekR1XYO7Wqig
hvHEuO2O6+zaa1zHFnvHmhdHzk6TvGpZGbme8Y5qnzHROV8msBfDKkk+OFtYc98I/ZkbZZnj4f/4
AzNPw/h5Z9xK5Xm9f0JqJ06VDeIQomP48eCnHM3wCxamVmOeYLRcbC07i/Qycfo9ggHQ+FVEnPDf
wNb/HbYqDuqcLqssYEzg93nz1YbRTCk++QquOUp4TY2EhUtfzN8WuGxqFHd/8u7lPTmUCF2Yoatx
ShlH+kyk+PiELrm8JvRqSszKqh91KBfvcL4Ic5PlDNIdp2uxAXCTPmCkrd5/vnYUrVe0WcB171TB
r6TbpTzUOqrP/vcuZv6xkcVZRdste6VVhV/SnOyxTokoP/JIg0jcvjA3ujT5WnPVtMsTW7BU4Rbj
ingu39psapEEoXzElBOXKddsmbmS87mb65ACxX8cJLuPm4E7DgjeYz8W7skw5pBuBTV/5SYAiz+8
3wQvcPYr7qfB/QOdmSdIwy9S3LpjHxvxHBIlNknCVZusjxRXwDqZ+YjX6wbf6kd0DN35ujXWi4NJ
IBepiHkUxiTUCvUtVDOwRyfv5NVHEFdb/8GK1+oJXNPCHzrp8PIhoqGnDtEJMTLI7YVr9+hbqv7Q
B2Bx8UBX8sIL1223gBfxo+7xTVbtkWteWj2A/SrYiDCnfLrEYk38FNH+ZYVMRbZvWDMt1uD3xvUk
cClOk5abEgBqPJfLWu1e+jtsVd01a2q0siZ+F0a4R8MpfmpH1+paflYPMOc4miVl/XpZEjjRuR/9
tmnKaUhjImS8hP+ejH/V4+yanI8YHyw1osfIZV9vSUi6tvioSLdKSqK0RSujfLLgudLArCoKELOV
q3dLL/jrVNEitBRqXOHhowUfaXMX2uDJjPafo5OIqYay1w5RkXfhvH3YB7Xj00M3tzJO2cXos9Gx
zPUS1HKLq7J6XKWOgJm1w83g3Dw8n7nOjXBlr6dj4k4LMQ7EZvoGsp4Aaa1qI2LyBJ6CT0ffezhA
wacYKrjuNxJJYSuwQAvur4oPrEtg8JeG92E3FBybsnfRwlmEePqruYz4xz/ASs5wS4diJb5CswkH
xXwkNK7GZogH29iExeZhRxfd4VxAQDCrgyX/5879KGmnLPSKXkdQ8YxXqPlkWlZ1TIaYxcsFcYGl
G+iEfsWkjtdwy0ilGbQJ8cZJilI5WKKzaLatPt0VX3miXoptnlPOGX3c1uMd2LGPy3/u+yH6UTNZ
rI7fFaRIYBIeEnuMLr5gl8VUWiqx+YKaD1x8DshQ4k1fvChqvN7nxzTkL5iZ2oW9Mjr6XKQUynf5
UvCmjeQ806VYKBjxIGW7bVu3IjgFFXIQEEImm/tiFZaYJzWtUlpC4JtevUYrIdnLM3MyTc1+TTXt
oo+06CnMfKW2eMxhAVR7izzt9zZlokkSEmK6zPlmClvSj/1P1KMj6UjUfDaWH6LuTPyPh272PhVZ
8ae+kCGbm/XzLHN3FtMlMB7o5SW8JBDkb/qi1rcYRSuUCN/RO8QEld+WkxnyY2zv0tHRpjjhE/E8
zsaXQdR41RqpoWedBfQc6e/zNmjXVpDvkvHOtbtlRPK+p/SFn2IrxxbbqKwP8Fz5dDAFqKfrrFa4
My1o1ApeT4996VAY+kCrdHha8T4+Rq03rRMZt7wzpma8LvyHqKnGjHLTBnu+j5YVhKzNQEm/ldA5
7bWM121xUYvfk20WMYaxhSeBAITDTWs1FAqYqwoK4D+y17seoNzFEOavdutfJtQQpZdPiIg6OVyL
4sFmxadhX1+Weiz9Syy7rseX/N0djbdOqtMeIcLC/yqvz0QsAxeuwAVwe8LzkoTuoWMfR5m0PYho
w9tgLhUu0KUEl9LoA/3cG/MGPGuk6tzJuPKW8pyzt9e2CkBt+97ia6/aemAIJkVJwfYbs4Mb/0cw
aXtTFAvLKDq5CEs05gDkuxNaWMEIfi70ayzYh5WOAcUQESdGUNW60VVhNXaOs5PHXrf9rA9VK1Zd
u+bKXZHtTSq/hi8yz/Nh1lDJcViv3+7TbV9VEHzps0j91LDQ5ML5G0+M9G1j/HoMGU0242gNimgX
ZpGovxnDhbwen5vP1I7pIbTn7ePofOCb08C1g3DFMYhub6EktIxedl/v46/jMN5Ffrl2ClJKgCjq
lW/sVDaJoFyjQxhIwSV61x+5sHbmsZfRpAVTiLc4aIVlMdodLUkJOsGOZJEM0tUkyyJaCrdbnQZy
sokRsm5wLth1NZVbtQp3MrUpzrJ54G2ZBP5zIHeWRo/27nly/8MBDWo3tT5LkwdKZtwqQYAERFCL
n4c7Gu/wY8hAfW3yBj4xc6aI36OiMcr1/cI7txyn0rU8lCfUlORKuWjWX5w18TZXyaPyIgKP/95R
oDhG86SEcbW80OxZLqLeBk+DEzI5vZa8ftQG7T2bIkomUnvIfSfjr4Bin5gQQ2LaN1jRJmL72iVD
yYqKBccHFX9eOU4xA+VakZz7fj4vhKYwns4QwfryXLEqsVnP1t9zKFsCugb/NPKH+dhjFmm56Ppv
e7QNh+rfpjrjhL3qCslpl04oNjSRjoU+QsOvykcTbftQ3/cGhDvo3W2E35nwi+2XMqdt6kGjux6g
2gAIu44g4c7swXeuZDNBHyf7je9vOs/7J6+h/3GMp73ylziAQOe+y8F4pg2rRQ0+AT4L259i/Ne4
7m9Fkz5kr2EYDByKiE3QRbnYwC6q21Jga+B4+TG0clUPAgJpui8+SGeKTMxYAF38gmePqMa9FST5
uHklWuYQMa/GLomJPUz2izMDKV0Uh8n2LcDiH5FN39FtJ1cgDlUzg9BPlWa8MfrTR1GA8rFRFNSL
aNc7eoJ+V6NleklCFf2XLgOmLpiF0yabNKCNoxnquMKz+DSWa6tvxVqg2hpsGIpXp8tdpj9F/JVt
fiSlRZMl9huKSdOvOLdQUE6O2zQc5Kxz6zKC4RtRcZmc4nC//p4kWIU+nMBMpG9Km3PIsJdMSpfb
XWS+oS+N4e9PfvJQboz1Nhe6T99TYxN1Ex5UgaqlJSUX4enaw+NTIo6exXLblUEOS1LNqn9oQLae
AacW4NTL1AlKz6isLbts+HBjncrIDnl9MjVFvCJjdePt5xX1LYoKEhMzLhWyiYojuWwvz2v4rzA5
vnmqkjqX2AQCYg2ckPuKFOfc55GusprPywiJsb8D3sdvcLoRnH9A8gCOF9ZhYoieNQrDkwdy5aEQ
D1cc111zL/Ofn9Wpw4CPErSz7H0CZBVp1wLqI7EAObsce2GbB+fa2dDk/wDR0xzcSdzWezEvNUnm
DW8ast7SF3iYEG4XGTNuDs8fDIPeSotWvMq0YXmI1vYZAb7IF4FunP8Bxa5kAhmKVpkeos8iDznP
W91npduEr79XqMOLz+523UHau8ejDlm2bh5rnaELYBk4n7cKU52+0K1N9uDU64jJMIJb/9DiqZ81
A3vugvu+ura8AC6Wij6cc72C3z6VKk5KyzximnAvWEkzza/5MC3qFNtmTdtdrJpEIWkdpQqBSHgZ
a6XidBYfigUZW3WBIPY/r6I83VHgMNbN/Nhokzsj0SWzPvaCJk4wSuRUNDwThuespGugVLbcefLH
Ahqh1Coh7r6A4u9otBZHV2Vs5op6pWMzWYhn78ZMr84MZAHqOsaHQ05Kr1pQIOkOs3PszE/PoqWK
lSex/ch3pw3Z85pd5k4USli/9O8dZo4D2JCyQeztvb5S8GZD9gis4V8ikJ9SDTiKzKBIQ6auJ+Ad
RYwUlY4Ml7Fu0bAUWlv6mnfiRI//VsIpavHkc3GWmDFlYUsvLLalxNhQYPJtKMp1iuUSPB9MbCOe
5UntScZw6+klc55a+inc1zCmMUNAWAiWmUluz/B4ooyjFFtIP5enW6+fG/NBp/pDUUNTp3ik8ypo
LWn74hpg5sGDNWws6sd8M1z7N7MCpLNNsC1Reon8iPuo3XzQ4nes+Cfaks1FAaBKqYL6HNfV/hLH
3uFKp4n7ZfW2BdPXDbBRFcxB8TeWGevUqMAXMlG/qtxrgTsL8+kz7t4AJs8ith7KAnC26vRQDdm9
ZrKUaIWDm3exeHtqVzBLUhlsyP1TSctK7uGk6NioNLPmxrDYyIva2II3k6AouOTqKiwLWJo6EcvV
dIqZhbSlN7lAxLFaLBQOCcydUiv/uUHH7zTPqrJb7wKnVZDUhvms2Uofq7Aqg9uuIi9T6ZOzgqvD
iBS4+RMnsihMI1fF85ZtdueCscMFobRRf99QQgN/fYBiaPLL/YK7WCPqOY5WY6/xTDzsYCVTFXEW
sp5PhuVOoY6stCd68+mjPcTx+Q1ft1aZyP2LkOz8gVNNhKHmK4KNxJGQbzK7euaMOR3WUo+i7i6N
967xXYonE3GMkNFnLu5PsOeiAFmhraOQUfFnB5jQbvgPK6YHPItktqPmArhEwyYrIahpel3Fx7Gj
xIe0Zw61aEz5utxsHD+C+fTveJe6wqcuxrWucJbECYx3sYFY5LJMI3hAmreZObXZj6n2BVpe+VTR
bdG1IrK/oKNpQ2es8iTbUZIwps+nENjX0ge6gcb8ACOu07cDxveCo6q5dd4E2cCWJrv/pqSWMAXf
DFPzJevJ1KvYxHde3gRUrNNlzZrpQSfEKYykSZQSrU3zxmvv/kypKuevZBzOStDh4ykeqeJC029F
ox87R2e79pCvGeB9trHf1nhSAzxEuuDY1ofvarq3GihiWMTpialv9CwOoj2teSAOMkrjSUX+IncW
mWD1ldc37e21CNPmSHkp1aGqcmS42Hdn7LxfO3k54P3x8BrezqLCp7bk68DG5iGKiI8NikwFHItL
ayPdDOciRbBOCKjft4y9Gq1RNkl/v64pYvZnwfGHdazaXNfZ1cyD7rsInmjNgbD1MbR8xZnRYgRE
ZIDX4ZI1dngBPI+/To/nEHIQCcSCER9XHZZL1p2QPW9/mnGqsKAO+Prhh+njAkbV6C0bCXFKVpOi
DAz1ZlAxEJPe2CSZaVXVfLcNkunbky2jhYmnmIZKOKUXfqQY2dsBnrhK2vVkzPrzvMNCOFD8i156
vG0HT1tXOApkCJdIGaPMARtiRiEwPmaeUj+rOUPmT5vmoVwJ5TTBfLZGDRwM8nQRpDohqzE/5uyF
WdG5d7RiPQJJ7M/BiHX+WDk61AdLofFJ9B68D9rgeYeRhAwij/leoVm76bz6b3SmVjIepVyZkWLn
6ggv7bh2+Rb3GQsqvdMVTxN3TvgQB57a2vQF6V/rkkL4IezpDsZ3FlwyODkCNHSYc/GI6yktAUsf
Le6ndivf4omrvBUE/JzseGYRDmPrnnVGWXapatyy+NsWLzxBrM9HLNQT75+QdGcFfwpFdUDvs6lo
xV2cxtVb5CHdB7URp2rjuV0GzG78DmTowbBM8n2KJZtHkIqMoKFMJX5HGPGTaZ0nc9JkazNf16Wi
H7WaHl5XZpPOsStMOjMRAPsOoxy9bp1bdixGdYGeZZH5vu4ZYHsRY4AZIxFdaccKdCVBbGAdw3kV
lmm77SYHc7ykK86sW70tM85sfW1fpLxttBch77RNAFg+Tm4JGhrc5kovCKBlpIHahxJxkE+GpdOB
+OOSWPuim6vafrNytV9bWOtfC5V/Vo10WUWfL7jGchPUWyurmLss+a0Q6TpJEx8NdF0y+yJrPtxS
t9Dirzi8VtlNKWMKH4PwunBaDqnRd2fbGFPpogYPvEkER718yeCvfiZNKpjIB1m2AYCylhUE7j9l
nKU8ol1ckxTcbhYfV+k/I90aDGfHhdaSaCDLxcz9ez2fU7E7FghgMuopQgOUYfqkCWDynh7QXcvS
UG2sxljOj8vjcVZPUBz2OsN0RNzLxKQfUL11quxy+4aMzomUDS11/UXBjUW/E3b6cY361y16Hth9
V8hCQYdMnylFFD9NoIjpLNKDqskY5MOtT2wAiWVekyEh3mWzOvxSzrNSrl35WSWBC/w/A7TIWwim
eDNC0V6sNRa2rrjTJUa+/KVeOSYaeGmO8GrurJ0KCWB97cIzf8m+oIAB/5j50t+AM33vj5vmD68D
HXjTFOoRllS7XxVkKu1Kd6MRxfLVHGjNiMITBGv5Bm15KU7uGUHbqZDexmW9vK1Tp3JwTPiLw1sb
s89XCAow06RsJuWxDCKJ+KKNZ+VHi5P8V3gHXQ2j0I3LHwQDjZDh7HcBBDRmjZqkyX8g8kBRxalg
R1K2OcCrxF8LnCt0CoMNrzK8gdGGtZUW5fM5ox8ORkyKJb7Gu5e3tKjWfjeNfHRMA8utkJWjtssQ
YTyFpc9jloGmH5M0WErYHHiPO23WDygibVr6FSDum0OdvXJDc+d31F2x+EGJK5Kn5bOGYusBRIbp
BdTCpk+/tY7ljt3CxLf+nCu7G6tGxpzfYy6hE51gpzYsCo1WO1IhurZhwRaAblZqOnqjoZCRqeN3
VP2dSWaSd3zdbwptZQhkaOScr0xtBK1Qo8D6If/rtstN+7Z1Ux+OFTQUxUKG83aiA4Ec4GBmttdo
cRamLcfeJxWBGb0wosQJMo03e+POLeB3NsopOP2a8BrfRyt9uyRUGFj1/s8C8NX+Ilg3kf2djr04
Wo6D8tMJtNfbHLbb5trGDFexLKokkBQgBQrVdbxWx3yTQCXxjyrzWh0jPbCC57tGhhS37m4tnAqv
dmA97hw4zUWPNwNcXbATsD6g6CTUIunR0meJ0VfaEidXMoJr2UuhZk6Igb5Yw8DqUNI2xVcmlR/L
8SXyVlYdrcOuQFefPzGrTAPmA7LMOSV8l3Vkk3d88SuksT4DLgQ2D7BS/P3/B0W7EPaqa3Egdp5v
4QUYHTzosm34pcKUQfC/QyHbPNJgSSfTWf1TEI2SNPc8jk6h8UoU/AlU/ECwkl3b6ZNf1hew7Ay+
MLYsAr2OVG8CrrGF0KT9J0+cIHddsJRKtVngsR1h/X8TC+qG3zQ6hzc3hkw3+//204+v7lQRbr6K
yFKozdkQJ2o+75VsGzUhjxct6xvfJc/hugMfw/CmoDmpX5JdicCtypUHopbjw4JY4yiIXq5FRuMj
pB4PLzr/SAJvy7HWgXIteNwXg8iwW72jvvBxIeiKN9DDs9t9rQWdg0gY5c3rGxRwXeWlREptthsb
S0AciQhXVxQgPi73qnyGi9UbpxcmISjA2nVPnwzAps9pbPXcbh6FGM6a02pAXnVVC4dFg7fjc8pU
TIqGX+Et/FKBub1ovyxnVG/CDYOLOXMpLi2EOO3pgVGMCZBMBokvx36KqNuy/9v95OKLUGhDsFli
BxwG5ZpNn8g4WGUjDJXME6qIj0jsICI/QOjuLiQGj/vcxk7YbzRxvncQ34VCaKyxZxKDCehsdf2q
EPQffNFG28EBut8cMmTTtIou0Id36BPWwLLpeU/4KUcSIbVi1uvTfESfhLRkI3S6KyyGyWlq0//n
7muSFj+BuagIixD+ajuhvQEhiot+NaNWzRg7hKvodVAyWWjrJgb8l9eWhlySB0ABrtFGarb6W/M7
2ICMjiaCO8bA5E+jjc+4zcYQCn8/yudp6Yc95GwtbtHmBKLWL0ew1IGFLTuKrp655PfRsxZHh43s
WZdsnGInnHAFjXgkdN5mV9bnamXB0xvzw/JFYOg2b4CI/Fh/6deZPM8zPKZILBnYUXiitG/ow3eC
JB+N4guKhiErvQvxgG/x5syMAzyryeKqfSLR3Y5+BJ+ADdv0gpU91oRF9mHT/ji0YM9MmJAS4JOM
oafw/Ksqf0olHJTMKm+GLAdTffwyGFuIJiIa+MXxNjy+ezgfyu0DB1lY38aOdt0zU466/eFmN1tc
+Nh4v42+l3//IaPz6cQay3Fg4n8yJQWP6YXWMSAmNt1E1mTJH7bqPhp/JDaTZbfFdg596LtYeI6y
KTMlkVScZlKOrQPgHIzVeqYTE39NkEOaEtFNck9FtJaD6CBm5r8f96Wm9xGLv8Fe/Lr6UJ+RJPWO
MTRirX+d+QJd2YRLp87Rq14UB8x2lE9yshw2HQw3q+nNYCWX+U98O8YheCuZs9HT7k/W5SEovCuF
XBJ9zzj4fEZX/b0Oj+T5MxKGTao/JAlKP6GVXRd4TmhYUQKLxdKPdbnV73sGtT9JNiCFLXRaj5tL
ZtwqeJto98mUbDCg/K6VuE2RAmjUO35W+B5ArJo9iMZ9/LpPRJwH7NHFZcUZB0+SG3qI95xMADnR
JeknTSXxa+PkBLfCG8RSI5v2pmyzJ0cG7GN+9gEzNJldVme9fLTV1QUhsBK/4a9oXEzi5IS0RjjH
THqexE3ML6BlqavBIpTl4y0lKGEq3aKRhJ5XASe1B1rjvsE2YsURUBgGvRZympUAHgyMIXeTUanU
7RL8HFKVtmcGre8s46arq9yv8rPxpg/rkqzsFcoeZyCaC25ulD/bnsYW0c2CUtcyUpEmFFRom+rP
Qtu8Nz3i92ASVkYg3rE5XJqjBZy/e67U5mHEMaluu0rYfi4XpyDvJ4i7S5coRYT1gZzKoMRF1AwK
n5F4zix6cB5BLnL3FpiJhdYMF/xIdpRgq4PK4NjMSxcgAp6ew1+66Cy3Fwfq1w7EQ4MwdgKbRj09
qTlBR2pXh48U2R/8MJXwWyy7tksQ8PHY5nwrmLGX3ZVOwTlHYtcbHuNWX5s7XDzmPDBSUBAx4wJw
OT8z95ZaU3b5C+bdytoVAE08kz5jGbpt8vprOwfDVimABBA3tf5q4i4PRleoEylACKvgTyjhP6fL
8IRhQjy8/gIgmRj21H1Pg1nOsobpTc4YgDM7udKEQjGlD6WHSTai89F50zWS3uxOznC1GmKbKSdE
jdulSkdW0fkAwLl48+zLsHTiTqFW7NaJDsRB2S6AkMQcgZiGTCOnMCR6kcY/wP+UxhBiI5isHoKm
U2s7BufSS37ee60L8jMHwRaaYl/9/akardQ1JCJuWXilu/D7pum6REPvYR1VTKehf/gJuoObEC4O
xxrypWTqTE3U2ppSGT0pjYRkQaTHZlNtT0GtGYBHdUxWOcBiz8QyLteZSunkfk++XG3sUkqt7hf5
vjicSyMscQZ22u6OJC/+3naU2Qn2pPGcq0DEcJzwCT+tqOShY2mZ+Jn+3NBjy6t4qu/cK43SKTQF
KNuVQ2yUW5x4sdNtsArmE4Bc131Vxbpc/nLMdlJI9JyMDhfABCDxpYglKwo3MF30NQXQ4GrdjPlQ
6xEucYAxCCbHht44DoowYDC37reWyLfcOGR2t7fiFvfDsTeaWtPREcXLFI7UDM14Kcsla4rmlDFZ
SSUwSYe5alHYkoTonbl/42ayed96YSp6cqfVlJczTO6hoJchrzVw5JviVjlk0SRmZpUyr1e4w5yL
aHxXOjvolA1lb2Na1CtdAhicAI7WWgzMYE7nOG1nHYqDkPZCuYj4wGrMMVXoTUpsHA+3N7TMRiEE
obvw8jU6rIBJA+e+MRIxIyUU8Z1X9XUK710lyChkf5QxdLBi46qCWEuqrkcap5BZP3qYVPYuswYH
uLUwHHYS4QqRN3f4G/keJbelz1sUz4CrcOJly57InaJ22X4v8j66c1luatBKxbnRqKyX+ERD3UZI
3ae5lS85mRkumCvxhv5tceaDOwUbCPyc+PTYNwudplMggvETSixyNZqljctIs9b2wt6n0gRgeEzK
tSr0HdnGOa8NSVVf+OqxGxG4QirMAFuJtFgWZy70kxtz9pwujme3L2MZ0MbpJZcEIaADcI4PzGJI
6m90GN6Kp/5HrCC+U3lTnWe1q5Pjkq7LW0aSZIDW5iBA0hPQLy+VWDrpuvNDROkolF027GJNiM9R
/oZE/McA2kedQxZzR4iZODW4y0aKdhV3OgkuUhE3hU+wEn26PbDtVQO9cU8NAXjc9oLMwnzbLbnb
I1iG8GpE9Y3O+8HAWtRpFHq2QogNydOVWzStRHuJboS3J/htUaurhKGw70EEh843ybeo/RcdOtlg
LNgPgxdsbpaADfqNl+sGJzT+FC6vy0X0ENDspXxB6Ypbo47VU6UEm2QBWCSbzA7ezxaDNrC4egSv
mrjAjKnAVhP5dZn7IQD4Ydc2rYaN3kh3VIDCejMNCCwZY+TZC0bQERUYfjD26Zf9pyQkPNfBihCn
dq3P6gmtrhKHjme0PKvzRQyxebbvL7PuHh4n2Vy2iHejEgrCyTMxgdXQqbtgU245qi75FSf3jIGZ
ZKwtY2oIVKEqJRuuhU/RZT7AloQr6CBNd0GA5ZkLqTPAobyoQrIGimwO2/SvCRll3eJlrKS9bLzv
XDCOLw4r8xb3RBLXrwA1kS0jU3v6FKh8MhARDfHEEuxuYX2oBkADOwK0SZAY7vcbOnfuzwZ8BBGJ
TkiBjW684xYl6oPAj564ihJa1B4yzuie5xIX8DeOxa2SJfVmGplExFADiJ2L0v4cAH1l9ZUdeevP
1YdbnHsu8OugIw3lsvLe+L69n0dTQmXzabqGdhxK+8bB5dFs2sqGV3FgFnx23JL3Zvy1soXspaVF
8wqVgX7hFQh5bczT4WJraHoHosrsqZt8X2Vbf70tl7XEiDTH50IHyIb34wcnM+zdDTi91pT1CHWE
DZbHa2b07sIv8FoYwpwUWRy+HTr5aagdppzXUmKIDF2Vv3mhyEUH2faOQjYZgpifdRh/1Hu36h+0
iDpf5qCf6H4vlgbT41ASvyinmuWwZMo7bTxMdLc+vJ9pbi5sDiGr8ynIgLr3+igzIkmRiFnTE6mP
2TKLlbWFxzYmtEat6illLYUM4zh6bKk1Kk8TxTEF2fY5epLDv5w2uL4d4lFZJtO+7/i+twjlc4KR
BPU26fxt4O6Pqjs/yU9/VBM5Gf/QLPpdkSy4j1Lyrw7vl+ytRBEdCk0TpQ8FC9i7S5gTfDuEFR3Y
DSYZca/NM7RQorNA39/LFZyvvU0ite69H5ZoGnbQRPTTVzM+TaaYeWCQWbJYGRUyZxlV/sQRzgaD
N91w+CfgTM0nPmICXTYEpwGRofii3oF34j2Ewvu4srDqAFPImaElZWmc6oGh+fOVNMLmhRY2XvUc
FIeqD8V3Go44UveLjHV2JU1E3hBfWh3T+F0n5VJe9mhHovIaFYVlQ7okvaTeCXA84tzAV0AB+QIG
i9PKZVDJLJKRvNR7DLrYBf/h/5jG24XA+W+D1BdAnDcpV2XFp/Ly4mbJtO9meRfMnpu1u9ZHy2Oc
kQGDquqEdngfHJqZVkFx72DE0wlvXRLshJ2OcFZOOnZidBhUDKhTdvj9qsNB5NeQD7MlUOOWDtFj
VR0KQik11pMyrmo7Hko+/EpHjYPDJNupCFphpbWrAsv87nLqGThL1UYH2NzNmcnB2TYmbCYx0rp5
uIXdL2vUN+QprEwKZntl4anxVg/yqSfcHhwTllgkxX3JecA0+FDVxHh+myb5rCSgHmgYBhtutF0/
FRUkz5yCzl1eUrcyoa8bzJZPAcIYIH+j565Fgn8Qbmx9KMEsZRnuPpg5nAlNMEHGgaqP7nBHntJW
xLjRcUF0L/m+buv2381fNLajqCrXfZcPxs+esL1SN/Xb3afc+SDjOLs5QQAJeK78az0PT9Gwjl/h
b/EsnvrHF0WhTKtS0T6cHeNSi+bjmyOx/iVLYmQrkgVmYCseSp+eej74QIKCZIKJ3Gxa4oMSHsdK
UwiU2LUGGWTRQmyacZsviBbdi3/Z1f9R6Iq7iJl2wxJmk9VIRiVah7wZSZj4A1KApCUMdyej25Y/
UloBMoiRUk60nDhxBmp3pVBYKvfuaybkX7O+ZBFC6X/Bs6g2fxiXSevS7yc3zV0F/dfjH1ROtjqi
g0+9DOv0bOePUkC354wK9ReqPtm+flGLwFPqliowxBrQcENZee0r5O8EK9TB1XdxgTjvp8Ix+qrl
w24fY/TqOlZ3O4Y5UpFtd31gja3pa8pLfVJ6gZ0Nc+VjNbrcz/ogWhpBATa/lOcGJ7iCZbw9n/7A
q3jPsXGHPbVzomH/lHy7YrICW7sUsi4xntl5SRVAboUGSGuOGII30hthliNtnd08eUEVFTrAuycv
Zp0i+PIRwe1QfpTfbLiSyEcwnMkRlaYkzyuHnRQ1o6AiKE8pMAQTbQb8tdVMSILLT2Ift6rUTRuE
sWR2ti5qf8miTQe8jLqJiT4AEBprJIag66KmvtTdeW3NuV8Ly00CeExCGA1Szc+xr/oS04DtEK7Q
0dgqaLuNGdzqm+5OJpEMc2CaY5XdlJjYsd8f6lUtSLOcOuB9b/coWg/jWgPZkwH3ZVJOAfmYsEeA
Y0kfpapYLBWvNkE2Qaia340XNMuJ5so3QH85SwUrjDs1OWiKAI7eLlTx77u+hXP8HSOfmQIn98+l
7dQ3VPNmtLLV/sn8qE++O9hnvBbiZq0qjg0AiHYsOcwC4JJYRNEQ5nFqALOGYcktnaIFu0eyLBdt
BbKA2Lld5dh/5tUdwl4V+eg8/ZVsXiEN+K20hGsWBLyN74UXfXYF70a1hVXVYOcMaSqB6yyYqOkm
hAP6whFsxNuR3FrTZ5yLToKZCXti/dDhOUmCNwhBZrVHTUN4bCWl4Tb0i9d2M0GtcnBcHhF9BeYM
kqSRPPXMEh8P/pyb4SnxBLkvGxR7r4SADZ7Hp7xDxYoM3HDIv95Ah9+3w52wJAM5v44h/Rr/h57b
nJhT9EH1tf2BXjl85xwbOYVkNezg2VqoOCxaRueKNEOYn4C79WWSzqVzjs086EIHg7wyGuzIo2NY
qIadDGc1zvkZV5Vh+0UJURuNq9Ss7nmX+ka0F7siLmoSOa3UK8tCZNz0/TaPbII8ZGE6PvhGU3OZ
NnkQkQKEhXlJYGsBHq3lcb5dAeR18lqLVXpv/7uNeiEGYKSd8+1UY1dzFs/dPRFTS+tzUjc22vzU
/IBv0dG/8jJx1EiwT1RM6qiH3DrnOR8opomfT/qvMWk5HSBJH7IMwD5aBm+bYz8TlljzYmj6iJ/t
ClxJomwaoPys8jATHf5otkgQPL8aWuTeQIDbjVH0b09a0xPp5hYPA04wFJrJsNRvGsgoS0lzr4aq
XiJpZFKwudBXnwoRHzewym0mwDNsuPOBXEZ/8L0kuc3tPgEgF51o8cTOL3FMdQVURFfIPBQfgmW1
qxtSP+IBCUpck0ynDSVhRrTWAbbQNXHSxjQtJE5TElilwpx9viCk5M6tn1ln9HuOujvXNU/niD0+
t+wLM/cNKym6AfMRpbgMpZD2jcLUqSdXU9xNGDKoetslWyj3/WWtLzNdPDbom8MdS0sORv3HOTRH
Z0pm+NQ9mRehH628C99c4ctMpF/Eet7+tmeujdImjfOjLli9U7rUVm70V6/p4fJNB/O+PI5yh6KJ
XU9yrcIMT/hHes0O+TmHbzD+vOVAn4UAPRwxh1IFCwMH/bn3g6wnUW0p4PyOeU7901V407+skrd+
XnUdzo7f8UoKRI83eQ8PRd/ib8hn26PrGafYdaXU1T2cvHAOH4AlVYtDxNMbuanKhAgs9AuHOKcr
9t8FTJ/vHK3TwmEtNsQZKJXGbRQ4cp9VTD03X+Ffnb2KEKPQ/lJge89V5EjJiVn+mniFkcWhowdX
3955bl5deeZW3zmQMO25jBU1b48IRPchDllGQjcPJLIuSzOGPMi4Lz1nsH/0EkgG6FaQGNMElMix
hlO42Wtsxtm7DE7SeFX8q/aRGP50Gbnu9sZI9ZZysprg3VUAVxJIIJ9OGGKSe6aPx3KPblsWu7CD
hhXchvNTBM9QBTDdgtb5kKinGYHA5w35nt8arnr0AJoFS5VKKUGgJocr1AgFE5CLvRY49jaV3DgN
OAhjnhVNEUPXKiS6pZrgQpPfTho+Gq0+TqzNQD8PUU5BtROL9XUbDOxl9KfABxdKJVmmNyDE3Hkt
obGgyB45xyc5H7uhonMNAtwnb8qwcdzZLXEpdeDzdj9qz1q8toIkW+7it1CaIRnsIj0Nd6bGkh74
ZGU3zntO6rt6+xf5VgweH/xyzXZKD4ITykC7Ah9h5QnL6HBY5pB+vMWS8a9IxgC3DRSSMGUZVJc3
3rO+guae0zHSqXwQv0XCd0aOM8OW5wJricmRd9wQtdNphSXYwy9jIl6F65AE/1aPLh92My6clMX3
8N7KvdvkApL2RszPTlemMbBJK3qNnd/TpfP5+2hsGKLuybJMZjsNrLEuh/bzKA56peB3TppXJ8j+
v5Vm1TyPuvsQMEnlFmdITRg50hJfe+xXVKwKqpEDJjI9cD80riqgYc7L2lDVZjxdZRO8V4PcYNOe
I0TBYdJ0YpmhAbNJq96Q5KyRveGxWx4LBFrzp1Db6w/UdqruviewaE7AxfuF9byP4S35cyU9AhyD
81C9UklSPMlKsw4sdShRinXvj9WuyZA/vLFGiCEpv+3bj8cT+3/J5P55hWXIwXmkSt7bUUbStbPn
ioubr9ZNWzkuVB31bz8mWUzM3iMpmZ1Svn/3gUL5Dnyxf+3WqRek6L2n43RMEkZVT8XeatazhOAu
VUIwGdZPG0qbxPsnVQItMbujoVPiWvY48NXRHcTmzsjW3UM5xlzOxsul8aXjqtyYj/7bFvbkRJI0
flVDFmpPQ0WEfZXfHX8yJSpL67um7Bxp/29T7nXlvkJcaERUKXhfc3NVcXELNMJFCZu4mpys1VLR
Kh/qE8Hbdqtv6D5wmZV/VakvVw9AhicSMlJTMo9aLgnc3U0IveO8Jk8EdUSAGkXQbdypviJD3jFm
LuOoWqD3FFwVfwuy4BAVmFP1ipEr9xTQAwuiWPWfNmoiB1QrvgI91WZh/s7+Jq21b+XmWROyYfo8
XaBTJ4sUmgCoXrK00pYL1AIs4YkBjqWj4ypzLvL9kYfuIVCVu87R72v+7Zl1uHTKQ7nY8odNG6sL
TE35hkeddRfN/iMo+nEg6mjPAFhU6fKojGivy7WnoF8stvNqViSCMLpaf2xu1guD/8gEBQJybxv2
jtYdP1A3ASy9ewINwtNAgFRSDT6mCVxaMIXzNsZx2bEoa/j5j3Vh+WZAdPHRCqf6ko6afqhxqGdd
eLLsMH3h1JMaTWW02/MB6QR9wCrfzNz13ZvtP3NF0lVyHxCaruRRbQymqajQQ4AYXLVaDjzHY8Li
KK5EkPqNNy5gQcY97O62FPAMQPpI++U8JtlojwK5qyMPbzb6RdLAacn5rBiIMlYNKT3QikDmKWJc
dEYFH6A/lGkPvW3octp4V6gg2WyIpyqGUKiVuSfOeXVXvWmjaeBQ0YEtl7GtGf3SfnDt9iN3VA0E
/CPUEYvRL6zFRWiPza/UO0YnUxkPwhyfHQ1WKFN5Jwl05Gfmdvy8EgfoQ/KCG1CZi8HNxc7A+Y3q
sejdobYRBec35m1YuWyS2cEqjKafYcJiEzlIIc4dCmQyVIxSUpZAaRO6fmWnko/yXeJJkFIK+8f7
nrkkccPzT0Cg5H8DrTcNKhZHSErRDYTBBATf4DxiEACNkvmNnJ9pHrHG4xKtsmtWk1V1WEFIeetb
ahOAbuO4/dSw0PHkMoqshHwJbIK1ZQ4kq9SzzHFgBF8sp4IWiaBumyhDjzNwzLCcrs5dknoVx/ty
m3VOmLPa2HjcZqGMO6VEPWbQuAXtyq/pZhcFTMng+fQ/m7yZbQF8wcp1SXPm3UviGoU8SYsSdP5t
aSXfnotAhbQ4Xexz8eNPTAktfQWXKHla9oIgdhZMkxpkv1PamHjmchGlSNiVnYuEdz9Xzbe2A3q5
0oLtodmjLIbdsyb2xQw8TQpc73dqwQdIDHDqKlfuTLaGmm+wJ+7/YHi8ZeDAPEm5AbIv44ElVMKo
Qx/Ll22T8LoPSBfKwTmkj9arFl8u9qvhl8NzqrVW4KOa9ze9+ZNRwn9OTQCGCIAKpa6W8ONjIDLE
y+dW2n7UZI5HOE0fRzn5MtvFA+dxb+ClLvoIsttRe/DkH3ZACL4n8ziKbnxFbDqOHqsIpfBf1gIY
b8EBErgXpmdYD+hwR/6rpmCEwVwenk6OxCf9Ct/hmYOWsMZ/uEC5ZERKdwsiTO/ehJXvdAAFOf67
7wCTg8iXii751Go7XaQz6enkizxuVxUM/oTpP71PmpJKgApALYcvmue/DLJO6NUEaKZrql2/uV5Q
WCrvAXK1g6HnxVKXPKBpyA5LCxDEqVBa3SDENoeKguId5luBU9hLw8kV0OdhNSVoM0bTOxCNaFko
6vNCbc1x1klaKIpCd//hRhS7qLFLj6cIjirJvWxabdhcZR0XXUuRC2ibIyPPHNsGCKuVI0KEByOr
vzUylcLH8VtsXZqlo5xRFYhUYLS5V7Eiii8Pcd5TWBunv8XDelIfiLqCz8KyknZ/0eDC5RtET2Io
BNF6QaKnlMekwAWQ29BsBDcF83k25/ADiHMhaGIWX+9s2KdwVO6+gJEWb11+O7bIBzoMpjXCVZ5L
dyZco50FVMBf71jAkRZ+TqSfAPropNdPQ1bW0V9J5rerT845tV95f6DY9pBkVWXlq42pVvxIpXte
ZJP4uwifmsKI4G6HVIHbeZKDAJY+X2JIHgBAhQufQH7Un56ZurMIq5um7ME2V8JPRNRCtI1URuhz
g5f9iU6cYtjar7dr5erxONkVUMCnS/9/lFQGnkMmVm0etK3ndZ0+qhwn4E+1jMKS0A2CPdl2g/2g
h5U31C0VTn6MLPMunoNjXMMOspE+I3huv8/1ki8V9+G+BU58fDkryW3Pjckz59kuLyf6kdwi8o5f
zPMvzFutw0ofbng04IDZ9ueP91SokCMl4u88d+5PTeXvT/mSudfvmPsRn4+ujqn0iK+P2Z8AEuHe
HH2etO/1ysZl9JB/4EVSZV5cKZso6Anz9WUj+OMhNAhBFqkj5ieulhuV9RVw2PeV4whU8/Y78CSz
wIMcyzp+AOUAHV6QnCEg8nDz18zkp1BdQMCcmKrx7tlgl09S0O8b8a+UTrAhz79n8F60ooukq9At
lbcr939ypslF4AZQf7pbLOjEV9/pv+fO2XBueAg+/fFS8UwVzZlsAnP7ECm49dpe4VkRkNUYgaT+
oaRuDW2sbiSOZMrZm8gd3N8pna2ZrXgsqqpbtJQsr0FO4w8PBik8jaU/qkb0MKPFANl4BvEQehqU
YQvRMMgFa1Dmqfy1xSyOKi/j7cR+QJihVTtiBlxpMSm0/hcNtWbP7oykyJ9iAsmv/qu/MJ5D5fqM
Zxui1jYrPLGAL6xV+dcPC+gB8XjS8xkpm6ZMmL2e1GgiTWJkiAwFO7/dH3lkVoWKWsHIbpq9fAlk
MgylaBEgqMqCZoQYoK2ZTGhlel5MVRwQFkSR9AWC8mDs8lFqQgk/vmJX2ep3EHdApmj6YEyXcR8V
RxSxfOU7eCGhNjMUKJuwnivJVh3wfdYfnlLstzRn4o/sne5vYHyJdzKAjlQqwsRjiqjUMP40wuC8
bonLTlGOluOgNDso4zytfGDG728P3GrqahvYXyZeG/8UKYTLA2e7Hw8XXuEA5BzUDlAFqOlfgw2G
vI5C7u4ANbQQiwHMQnqBLVS6A5Aeze/xqKT20uzpocyGEEOKy2Af/uW21mCLdudk4tNcZpF5lkWX
hHpF4rPDyngVt1kr5p+ZTaHrK1epV/mCiigcYuwd130EF/usUHqG3oMbLOMGnJCMOigr/LwuRikM
NGMASXj9b8noACZIDwN5uNfrd88NbPiNJNFSOKvANG/UymAQPVLAA4xc4JR+FMOO4IARePTSYilf
E11QTogdMQkaKYmECFY9wQHg+mSv0bzb5dKp0Dc5pd15Vcw9OFLpXSO3ywc2JrqiKjy3xHngsrT0
OaiMQz9NgbbdV+uuPrQ2XBmj8adJi1Gfqz2l1yFHR/wRtJINnegBUax/CNCm7isZqDGGVZHxndwR
doL+VVfcX2VTFOgOBm7NMIacg57IAwbkYBktwdFva/JB3t2yO1IccfWiPTujxkLDKIarzE++sghw
C63w5PKRYtLiQBoZrBI1F7xJH2qBuoRc/dyIyvdHOcgd84YWNEfi0PKZ2rO4Awzd1+MjPTbXRA2X
qrZAKOnys7140uVTjwS3YNe+h/187RmV8+Z1tlrni3Bf34fly/jlEOC8Z0Khyyvzm01WC6FK4/Oo
85Ws3VzMKF2BNMnRN/uUWHo4WkqkgGYRcXhFsb20EZkWaxa8fzMznQvT3JJzO0YE6zG5JGJ83dvd
hQ3SEVmouzflYKGAtQt1fsl/LCw0NgoF1UVd8RwywP7EewfTYsOSqCvCPoN7y0+FNqRAyQN4dpuE
URu90nCUJE62oj7g4E3C77kVkSJTiattqpcnofkdWMThmLFaPIXLFPvXZghYWR4WORvCrevbUvxz
i3U+UMQOkQhoTy2JZgRXh0zCRZ75SCVMACDEOjrdCjojVpv+AeQ3NK0ZzP+2mP869p/TJLbNejRr
wSG3HJJtuBlm4+NCAucJkTSuDvjddur+QgwbqxN4vtbjLC7aOU2oQqFgz6HGpmPDyAAwetS1bJz1
hyr1+w1zFENo1FpPjLUma/uW9FGK89tn0DWjSWh4codcRUY/8ZXjEnHT5jHsQy0NHps+o0u1n1NW
eSMP+L9X3qHSsiqGtuHuZl8bPbWj1h/Nr8YzNdHvmvi0msSTioDSvku3AC0uCLWn14hW/12UyaOx
CoXgN8ck61Y9JLCyD2lSOulVDGTC2aG7YW38g8DqOGtEEYmLOYorO4im2Ck9p2UuGFeYmNxJXEa2
tSHL+HGYklxb+bg9FC1HzBDgZwydLoB1N5TxkICLfOyep/N9Fah8FivDHeccQPmqPZS4h4u9NWbT
remJ2fMkPjuorhg9btwGJ60PEkvzEJ/YtYu0hUNFB9+ci1zhNTvB7aBWD5cwyGrCq3PKL2OUrP0e
ECNppSrBimWP1jzZSaYraClzh7j4MIuR3Mi1CLbrfTOMvyNyTMnbAktIwNuUY45UWBFPF+jtGsUR
8Pe8TMwG+gBWPzD7omSBb+uwbr7KCsePWZSWz1Re9s/jbOqbOa6chytbXa+F38eec43/ebk3LtCr
9xB2WgxHT1CTvyEYhMu2jyk4YEN+uztlL5nSSO1ZB+xyRcg2l4ggaphVvG9NtQsgygdu6srK6qxc
kmEiKobWvDVOj9awyu3aYpdq5Mzw0P0qG1+3YeZNbYXBykjj+HM30z9GbCWrGa0ZnjTXgkghPBPz
PqUHUoMX9d7f9Hq60faaQsLt2NErGQR/zgOprhBEVXvfgqRGITOnRPI8M20Yjw9qzrusojM0PR4X
0r7NjD0fM5UmQrzbISFI62Dr4jwQwX/uF3+F5/ZRqjlnhIxSGAh+NqN/Wvc9NVg5GxQ7PIdJKC1p
6NxkxXeNc7hy7GFxYxouiusLM6ZD0ykhV/sTH1vOptrc7vophu5VUd9TEW9EAawURp54dyzGebfP
NHuIxlb7327Ly3Oti+eptZEyEdRMiMwQo7izivH4qqxXUMVOkL0/I6N3KRiPlbBaFOZ2E7+uXflZ
lV7fUiHeCkXsCTrAYRBDksDuB+Rc6S5JphH5tQ57oltzskiCntn+9ciUZm1xzpsfDub2G4faJoV6
3fpCeFQzCZgdJ7yELCoOsIcDcAl6AYhfWIATWbHb6bd7jT09yae8gLvaz0KUPO+6TrvuQ19RYtyg
3XyP3I1hohVADn6FsL+szGk/+32c1N5PJk5EkxVgwOTbLs/jKskVoUNSEaTRpe9AFhh1UZaUb/Le
EyOpOowd93jEufUdWvn7MQpkxPzjEbghRqgUdj+KpNw2dMzbfZ4jMfAgsy6qNkO/+Jn6Vm7G8SoF
Dz0wd0VjJoH7lvk8PvZM4zUTl1kIElrP03MoZV2+py3Ac/apZ8XXKSxvY4uO5eztyhp0HgPPZ+fv
v4BW4rn5rjcAwoPbkk7iwe3byq6kCXAYPZ5tkIX+C4ag5WrlmKPOtVeMURLGG0tIJrn/I1+CCAcj
57uwHLQTeO4oad3k5OzvLyAbPfzjPyexcsahrG7coUJPD+8jTyiQ6T7/WD7qnHtRP1UHvcgy95oc
+wWE92JeLJrrWReqb24BgUd0iRWBAwYBd1TLBuu0U/MZx04lZXiutVYX1XG5axfkC5+Bbr8Zp5Gv
2ncl+TxZ3bYQaacnQ9bte6c78UfODoiSJmIteRZtdw0hAAEru7dq5kl3xUWYlqhDDa0/TyDstbQK
MQkzaqEaXuwgb2dm1axVJU2/c/JuPgFSvTZKigmQIZ7cJkF+CjKPTIDdbOg4kIAUyUtNR+fn/XtG
2U2m0g5177tEa36DokYsZ2Tim+BpdJyj7EzAIl2lj8NyMq96eH51hlCK+hyQxPbk35zPtD3MzAlH
fhwpwVxCwbTbS24N6u0/JA6oXoCdZHUG9UOQ5b6mSQ04oo2A0KNPCXx7pFGAfsRCXFx9gP0EkleO
ooeC4NT4pwe3jQfM9rw0Cj/fO02iapir5tdSfZ40V3UkuDail/9TDBsGflR6zeutwMZlScpUScKZ
8IjZf/FTkex8NKzqLEQpvNletgORSD3VT+/dQ1IXdsmEACwdF1V0hWwgcj8yV29Raf9qLY0q7XDN
dK42lrSVrnN8MBmyEH6i/yD/El0iBfsMDD9fVjFRTb1LetbYIUHxT7BMMlaW8mpM4eR3hZWFlBpu
XhSh8cYdvlQb1VLAYeVyPOZtilg119yQZHXhTtpsgL78SAPdwbGOu8gj7iloF2S0fIzfVHRwRfUL
KsQR0fFzyfEx47T1Hi/XJ26AVeQJyJ9sHkg6DT9LsL4h83vxtHJwEvbN+YsGyAD77AF4uh6tNSyP
egJViNyc3VbdT0m/CBCXynKU3NxvOksu7YdEkFcq07pk3vILvsAr/QdyCh/R7MZ/7Qa2CCQ02ZnI
yrbIV4tXt5Iyp+pwxA2EarQ2f2urvkoi7awOEDhK9fhjEsxh766Tvc8N6M0T9X5UArBHWUPEASGe
rO/Oyo6U3rSo2PlX3neIDV7HWP2XeS/1ZG3remNDilCHkrq8gcIZjZUSas3bpnylVNDxMF5OO1Cn
6WIj9zS3VQOkM4Hac76cCc89DlV/24pP/GzIzFR9Es61we5+NFNHVUgA+v4PI82PCSErFZABj2sI
J+03vBVjAGaopmdadE4J1NjB8oKVdy2bbo8ulLRweRfxMUtPdJQ9xzGwg6gQnoMr/g62VgBoynLr
Cegd/PrMTghY7jFlriwCcU8I2jMCKOzkA8ZoP517+LFrbc44YLTjBHKWLbXvDWIcm3zWg4IyShCu
ce0503UuorCWwiIimMgTyVNBJC+86O85VZoFfRi1C/geN/Ei0qRm53fGDlm+Xjrnx42zVjK9x12M
xJg+Ar3adZcX8Yovv86L3s9wEcv3Ampdi+08zlvuQFN8OJH4T3h6K2q0bA+ZmWeQw5HzX4NSXzZp
wprC0nnAJ7AiS/b2dlR78TvUxl7Th71+wipGAPHA1fnOfoezCZjjm2mqt8NqkC7eTzIryr+bvZNc
4YfG5yRmjwhG+2Olvm1XIgISlL9TZEuZmkjnZKxy7UzvkfKocXoqkJKINZsG7d8yBg/OBIYGNVGS
16Aeq/MeCO0GKHEK3SHOQWZbVJXjXH7Wexui3SiiArmcEovLXV1hzYIb3Ng5XdlANzCm6xJPY30/
oAqVoxfOL6razWEd05GOfsx/9WcRMu3/crCUGP+52dlGqcCVfMKvnni6g6q7a0rZJmLAI2nksvss
B7dpWEcZkK2Q6t4U1vlINMVEq0b9Zny/QquhDbyvfCWFK48tox3TbExRHkn4r81ieB+RbJTcsZXe
d9pgx73RLd4N4q+lt7Yl8s5I7JllosgIVn104vvUs0MA2QD0wvYTJTpdmImdvmxEKqlOpSD6gzX+
ME8jLMN605MsZctR/dfY5kT5slTWjPM9wJnRq4+Cx3VXSBBWXUMzMy9Mgur3xN5phEuANYu4ayXk
ujgNEzdmZgPf7siH1FBHNoJwPg7b3xWp45PgMx1yZZY1blmIHmJDhwEpuSdhhru4dKqk97i58NuD
RQoyN10uUTfQPtFLSoXHwA8cbOshBOG5TvCSkS5Q26YkNPkmX4DKH0exYYXLMvSQfeB7I0979+gy
rDZgYCajuOj3Sx3HCx2zi1kvbkmp15WWVbEWGvsRunK9a6SOHGz2fzGoKkeYCZc7CDNxCvu8uuyd
/Q6D9s06GoHJT3Po8saNWMnMu5Y3Xn/9Q9VX1MUx+V2kLj9/QrCi7Dg1U+lNpJpnbJfMFJ/Svn1c
AXJ7yDwikzrZ9oVm4m6LJy3+vJ+WVliVfvhbEzFg2XiwEmi8ibtBGAzZaK8g/M1WTWamPAA07OdG
NygpYVocjjBGTAtJ5BAC+6ov8cu9jH6lpvqoh5OGh1guWpOrg41Od8fLEjdHBd8cAScFqmk+1EKD
jxrt8Yr+zP2eK+0VSIgi891EYH/Y3pEEK1gY2tidfH+NF51ONqyO2K9gm8ukVA69oWNbG8wIlGAI
hHpmh6tgVrr1Vx/ZSmp6ohZJvKjcsHFsmfOkjajxVllsUYfo5BkIeXudaQgDrAtmlEVX93QVB8iB
lakFhtswoYKCyM0wzeujNUp/OkTSr6euhpd+o9ImEjuFD+dHfbTaQlnZjksZSuK+NFTQmDxK+Glf
C9saMrm+lak/6Kl6UAK8amrBLnAdGD55g+Vbf9frUSnxnZ598Nx7DW9RGbEgMo9wfJhCSpQaFMcZ
XfNRu50092CP1kul4UEh23KCPdIz2WGsvYle67RhRWefK53nFRmREFJDj21QL4lIunpPT7AmycEV
pYKvlWZeHCzGF/kHeH3a/xE6OL9HpOiVWTX5YsYb1uQVqHAiPiXI8aOgpPqokVKI3CP20DWtsRLK
NdT7ew0tAxcF5GJFJ4xWowMnzFWbhKOSeNh+JbUKgf0j+tIuCcb3UqZgU/QgTgGVJzaFY+v+CRu5
FatJfoepbo4vvOdMWN0NUoGALOz+9p1yGZRGwHxsI4abRem8VvyTT7ypeMMxTtDljzmDV+XI8jWp
0f6EX1lco2bJstHNSGtv5IpPR5gsZQkzydh+5c+zA0vDoXwyryG+k/C2fRfIRIVDnz2ZJfrAxfNJ
luGBdy0qmaiad6P5Vu8H/frf70AKuTaFXODnMAGtnQ/+1yP92PdxPHU9EoVcWbchBxati/LlFpng
z1/yBghEm8GOiPmMYudnewNRi/E37pyhLAt8eHy69LX3cQDjLRuL8Qg5ebIoTAcHiCIGWpY13w1m
A63Dm9oHusqvUWQ3QkgiFy1ge8tYPVqbLgLkkKjYPGMLqHNGJeYEr9U9SMeJELPKuDjYfAsXBZxf
KQsd9jvPoPlbG5L5o2VwEofMY9Bt9gnWsmbx0DShz3u6PbuV13xwkq9L74cfApAxMWpVq7Ske6D4
bNW4k+Qf6PB5f/wmTXPR0qMYPs32rmtAsYnhPtxyUa8F2kWXA1tALJKWf+M4iZJLWxBZLW29GL8M
HxrLUdKL0JxesBEJ3ijI8Ds8Cq9nSZNb1aQs9azih8+PwvueHLJHXpQbFXO3UKKsy7R1nQSWVxn0
absb+xzBk8hZmaLRrNFmHY9j7byAZwd4jDnYhzhzX4VlIqBw05PEdLAWPFm4RT/gekaAptVWJn9Y
vE7SFPd3VQ6fwoJBMATqwE2yHZ8aFxZMthfjlSc3KKFS+AYhqtB7wZvUtjBfcUVOSw//w4hucKOg
fGKrY3HRWYCcSBloEfLoiQgcvY3ww3JxHcsIKLjyi6vg02UqlLQZ6MOmDNW85oZ63YK9xrIkcsyO
m5DrDxwhoC7R54kLtwspuiUZ+XX3cG4CC0U7N6bEXBIAXq2PfBEPWX7g7dIH9KshKXG2QmWeOu53
wyUOPhFBWLjQHOanoWUnEXz4HbzHN7QkLWbjqikv6A+QvjPm5KW/kSvdWPY01vc8HX3XnEhsGmNV
GyaaVv5nopBuTwWh0vy5wWo7XMNN3vUWMj8OXhU4nIBSM8d1ZWIzALuftOh9hTYB8XRZHjWIczii
0f6YK1cCur4c6xnG/zvar8G/zvoK2+TsuifHZSRRq8jaE4TRsFtos3GpB/cPYTta8RukLFtuieRU
Vu7FAGLPk/U6ZUapsNXzTgcc/+BL6olmXd0vhAA2vPEMMy3qE6ETN12tQoz7W56mCU5iiiN/WB3F
/agwNt+Q09iMiHwSEXutHHSya1Tsfh/VZ1df4Bxul7Wn4pjlwH6EJ/qvGmNi5aoSxBhKNMTl/AqE
BxeUIvcYGWHPDkgPw6LOV+96253rWA1OV1MZ75AWfTOxC2PkQWRMXF2JyRzwGbp+3ePFer41/B4h
4rRfbyBfsDNILUSD3BDqkHMh6Eg56Hg5XaOyRnZXJvEmTrIjeSxBV8zyNuJromeNLp3pd9Ao/7ur
u23RnX++EFe/AR4l5AN/udDBUJH2PdsSxMadWubfY7P6oMwy6QZmw4KpLDdkRPX+TMeiTAnnnVaP
18DFGjMWH5chN0UcTT7IPg0wB84i6dwcUA3OSACSXeMDZth4+RufhSPLY47vTxPZyxrkLR8Vx0t8
gEpqATIo5omzP5PCdMp1CU9xE47SQSuB1fRRubJXfO13vhyoMGXUl4Ody6caH9warlLBR/N0RqMH
jfQJtllUm5r1Mkx3vOZM/bgCU4VKJvT8OxavAC89UbxOpWy7jJP5jOoV6xMbu5a2PmVywTVWVo6a
nMz7rtJ0KbRiuUq1a8yRNMnpFfgDaEy/Y6F0djwRxb6UKmQCklniIKsxI1M9abrxuVKKZktDcNY6
BFJrvz8Qu6bwyirSTEaoxq3TLc9NlCjwDx+B+CTwIGvqqq88PP8clmm4DOeGLZNTqbQih+uahJla
5LFHHN5fw6bqwPk7kJAvwH89LesuI7Uth7owQexWByDf4ou3yulv8byUnr3ST/mnUgEiySpXizR9
wjbbBcan4fuwMl4Wf+Qrp2fKxazLEKtXnJI681ocB5p7WF8sYZpnT04ahXfZi1cYjFQS9rJ0WJD5
ztklgiWMyDV3iQtSZ/z4qzvqr5Nrh4nC7AY7cODkASaUTb+2dzCBXuFMaWaUi1G9Ba+FZZAKkZJY
9v8fSiJBG+U3mguTZfsBi59js78M6kK+WNk7c84amRSQ5v1DWy04ZLGlcoASdF1hIdAccqXbweDQ
xeN1Xxwq+BIwhPHNcAaN3pXisYsKn4n2z8XUAcA/ntT0nXt97qzmvLQlzn5ceLnX0drUzvH5NNpr
Dna4dCmCLKbuDS5WMkwR5uowsFsS6q0OEz/DmRHkk9iK3dERxtiRKWSyhMGwvOq0YqTqMgTNZoCx
hdqbfmtZGC4OsPC8M07We8fqCCfHqAm/kNdeyI5fNypV6Sw4OVfcueRH2H8xHcxGfGdSHY6lsuLe
AT4owGp2YZGTp5EXvXsyjxS847YuIn8mFH5Kf6hcyitTQWRRwsoQGRCxvL7SiRm6enq89ZnsEDrF
Bi34Vsn+d5N1/O9HsjnNBXZv94qRw9TfnBa/TrXTgx4tlCccO7y6vfTaB311aLXo2h3ARlazEIl1
6KkScmvvDJfrQZet3QU+a/8CABxAmDbaHyP+Er8kIHYjOkc/iNwMdKuIlEq0TwNCGZEV/aaOxEfA
k1scK7KN2uRYEt4mRtzQXNg6GP5ptkwutZ272XJVXeh79CuviwlyTsFYxQVssd4I0jqFQRKRH42P
fEiDt6H0wMMvupofRZSFJGX4qbZo2fpzf+JyqK0zpLFYvsNj6o6IeEaAW3D1Ugurs8Ew2W1yfVDf
VgEjhGQBOJJHyHP+Jwyedf46eIPs2q0VpkR/jWYeNgDgE5x+Dx7c1tYltN+vzaGG0ZvbT++L+Ceg
zbB5UdRb0X8uOOT3fUBar6tsve23hRiNkZFiGyCXQx6nwAuj3JEOn9vbgAzT0i5+OM/6zpnWnezx
9CdT6nn77rVCbK7OQt6DA18jyS9MH5RfpWY/WQDz/+AGX3vNABeWZQhUxH002iEUacZ1aDXIXpST
oc4xbkX1MHmksHTi1z8NbKe5N8i3kob7igwk+s5DiEvs0kUwHtemwyzW5SgOOkkPd178p3Vx/lGx
UlP6sed0hMCYUoXoMW10mXvPG+HCs2ortccYAVz2gbRlFZyldf3+37vv2zZq5XrUP5nopsaqdXwd
b12FofGzzeRMFc1i8MzRMWfmVACileCZIYvZ6s4+Mr4vts2RLNlcjkPyj88v/0OrXB+QIygAhk6H
dwmtVoOYQUV6SJCESWAGrXr5fCSPRbKnQa8G9wugPyVxIiy8SjSGPgTwn3dP2tojpl8cz/gUq9ED
JzdlRvJy3q+Zpu5L1R7zdWxrKLr1pNqnfiJFqIGbZWx2eN/9JD/XsLQdeprSjhLhNdZyGiI3GwCU
HUwG03MxwU9uSFrPzvH8bSgQgSQ56SV5XSBrTbe/5BSMoIU+Ce7gRv/2suR/zWrX574UO6ALZNbJ
w9my1XialTKsftG0BJw6PFenUosnVUmRQwANfihKwOO1HBukkRtC4+B6gEIeZl9sz8eVqvILgVq4
ytx3egtWH76BcjibRX4KoR4dCeRsfQKVGh49hwFDVmOFFLRSWKAOF+AZ4M6nykgbFWpuwUyalTc1
Q80wfDiU5BpFTjS5rldSAepv8xH7MHFQC5YJBIi6Yz5m9Lcpr/k01WiKNXmX5cxE6gOs6J4PoSk3
bLKbqEXXLoTRYFvJtvQlxQc89hvRvXyHiXST2oMGmxqMwH6F8RKEI+mR0yOEUV8/WgsjzK/c2HTL
VxWJQp/Af6PllN//rN7PalPdqUlFFemzxIP9Y67SCZI1m/EgmWZSjgHZoELp9Awdrmt2EhZguoTT
1Jwq0/9hu8SXev5gESbVhOEsdxM3SsT5uYB3qygZJYSjQpFsYk70oitx6ty7wQg4rttNO06qcJo5
DGFZLZjQ5n0twKvn4lBnbA0Bls5BHTiRAg9g7PAvQZXLo1I+ldaFHNHw2XMNyZXQzgikhUU5seGA
BDW+TJLOT+uq0jRdDkNccXYW0SUTWRogWk0D3SJg4+7WRv4eGdoFVMrgFv0tsM62HzTtyWce8BOL
qMwZmyxJFjkJERwL+aBA/i1gpzaDXFVIaWoUv797gr+/BVnrxmBI6mjROxVf2ibtgQk2RXHJjvz1
uXP5tAVNrCD0RsynK6lOjvc/W8QCOEZwIcGXxlCCepjWvtVSrcpSPK62raqMdk3JKnM1LtZhkxAl
OPCDzCiSYaTwnhrZmLlghaOHaHhNW0tD54rIRCb6ZlyupzATWFYlVhL5P/ibQJLnLMVpcNCXyYI/
exAijO/t4ZhnRih67YJaDiW/ESMFm6zhJdZIIcIc00uYkAG8P5Ay9KtcbP7xMWTZRmJ/uABaH2NH
Xb9reb6kGp/A/34HfPaBhCJamGgYX4uFxrxbbVNtCuqpMCRSjTsrRezLr9FNTUvLt7G70069vuK9
gNqtYkPaVZNF6sEVOQIplhPD8251uf2hC8ItjiQuTsSEJJlgrgPpZ7oKoKq8Kr6eue/g2kNk4Xls
jrD+wmKB20C8D5W1zEHoi2FjqhBYhztQoTyXc/699IqbLfjGT1zSyMXkvs6/IMIslnVtwwMsuIjO
2SZgDWoQA+svCMKLKcVYTPEHs2pALueRAswEWX7CUTC2Y5XrLONyyrO06BSSTVSqpZTBsugMgA1e
zAHMdxT6TEUjN9W2iuDldMyMsXRX7JOvaWbdqWxKCkljbEkovKnuNdPGvVWbKyi7PENqzxW8Rflc
KJePfmjsi5e/3jtjA4rHOaM8YWcdHPwfm0AqaCAUgxrtbV2mYNF8M184CwAm41/Z8+hwDxjb5xXB
xXWUjo4RofF/A2s5BDFRh1oAzr2/CB5TTKbQp1ObyWxdrvENCsGunK9k6yfuSCGfu11abcdbrBQ0
xIAxH9MwDSSADcQHYWqGXExIvXrqlzbLUFfE8Qgpxc4OMhRbPxPTFRYwOAg5TGvtdrRB40whxfFQ
vLLkCAJFgM3JXZWZMBX4+oaFmfoyP+/Q+eGuPMn7WJUydhXmMGxzX9bSqNrEnS67zz5L11UsIKoU
ySlGz+cIYgNMIPTRRRsNRrly4Nco5Z0lrpVUaUm540I/rYMSti7oH9GR34Hy+I0z9ZzEd5Tu/Bpc
qw3u6qHSe+mH8IBXQcqJZXnjRxVqRggfkl2GWPGDrXkMADqpX/1a6wLPP8yKNE6nomdpDrjjVXrw
ddkXS/tzqVoQa47PJIq9ZimLe54n6I3WNn5IxllTCh/MZ5zFFOwiV5cy4j9HSZJZDQnm85r6B7P1
+7zKRAjST55mgr3YedlbR02SdFnnUVBwOOKbpro8gHsrB0I3JIwGtSaR2kGJIp+pIU03rdTBZBVj
ZHDFJtoXmBbQYHbjsKImcfoFcf6AI3Hg20j4PYZehyXbIf1HywH4ZPRCrdTW6qPKzC9GGOONpi32
J7uGjCHFB+qBaCIaUhGsOc3/DZw+zZJdoMufBD8rbLyzQFLeWfi6frtPRKokEEE33ySHS2d6d3V/
cLQoWaCQefkBIlEdmABMye/2JXPgTxSLEmyq6b8kh6e9Dw0XEt6gfBgR3f1PP981V1WomF8GOByP
Mj/g1IL/cOUi9Aj310JAjz5E8Bu96AXJn1l+yabsGUfD5E3oEoWHt+mF2z/H3085FHw/9+Mhgr6z
1EADFeHYp738X9wXYCquEtaao6ZRlpHDFt8oKbvg+KA8XqOGfNr4yQG1sJUCULcZB17vyXMdHv5V
IqAXv4aVXOD72hfPp6PPSiihAnrhNJOIsPR1l9E//C/XdVS/NTT1Y+x/hFB8QouJLI/QmSyH/0M0
yTZqdpeb76dCyzw/bUpRUCj0Znb2zaxpPrxvTHvjq3fITxyYJkDO1Lmccmm6OvmqiK63c37kb+fH
2wYzwiOEGu2KxsZhZsC4vhU2uX72xViKvt7BqIfaSaKQwxfvK+tTcq2NnAQdYberio+NIuBN/C1v
8eoWCc2SxFN3dpyTalT+t4K4A1SMiJW2t+iVPee+uoykKYcl/JhvycHA20BXLOLenxtBNaonji6d
zKb7WThzsVx/nyCF3vvCzYPg3HofH5StW0i+nWGjUerru0fefCw5aVAXDFhkxJ4hrt6Dyn+rvQ/1
SSdWbPLjwsXDw83pfRz4aPX7mg3T5NxolJaDetdcUNNcsEiUn16VTlHM3vWPc/vzsRTo1PSSBHjs
LPxo2eUcmxlxngKkL+TrdMv3hDRGT7Fai1/nYOBSNRRaXEA3yJW99aefgo5U8X1Fw6K2SAXQWQCc
sNv1FgAdKpS8Uh10v/RVY+cPR5tkCuBvOKaYMCwVDZjmYj/Q790Vn4XNUo4wBMB0efUvOsNkGUFC
Ih8TaWKCBmL9nrZLYz53uEDrGvyah+7isnGs5y2W3IqRaHXlhQks0LK+d0jQkUbswfr3fL0C0wlJ
u2Stg9VnjFekwwJlKb+kKluDadyprl70qBtrLW17bya/FXESy4nfPIlKn2yabk4tvn2mv3U4vxAc
GtX2AyvPRCh9adfWWyiOwIpTIQZMBpIhh4oKk4oeUeW42tpU+z7RmOrVkGjhvArtpbY/kTf7j4kq
pevvA4D+wwYoQHWERQ14kleBKsekhHAHgpfSzmXP7AkxeS1VXqjOsGBJFS4iG07anRddrvVAflte
V9YHD+lf7L4sVvoP5Nzep0rVyUjSAk/SKRmZpZXhxNp1FUBYTWyVDcNg2ukizdJGieOsGFYJ6KxX
TxH3RKYw4eZ4iEA1IFCEHIK2hfRKnz8awLA4g5CcvfQgjBlVucNJpGspk/+Y/WXisVOtjkargd+v
oUMGLcbgZqviDBOOPmDUC/nhcHlXTGGOHYL1nCN1kfcHfnNakqBGOorhPZfGb8tY6x4eg/7iZ+yr
2kNB/1PJgZvrarEYHgMl36amfJKJMuUAKTMQvHG2WAGKv4d3AJMlSgx+mvpwSHBt4AXyTu+qHukG
oX3iukwXn30Flf8qP5zDnS6GaIuLbciExvrZvU56/XaHhaO+/Y8TgWNsI8zG6RMv9cVvDEI9YcqV
ToLLefTlk5JZI/m8kreyH6J4B/d3gkT5kc6llB03OzVdt0kNe5svzZuVNuo2fjD3wnfVdX/+uot6
3i5DkqJduIOX9UOljuvyXqeodUY94rPbth1Y/ZuN1e93Lphx8/TUNnsvA+Q/zv+Sq3M6DIa3PRZu
c5zpGtzE1HSHJcyQkexuH6bV0+ilk62yONKH/SZjzAqBmexJp/C9iDR6sZfCqbfv+eEFZSDmw0Ed
Wvq0/N+LaHK8xd7w/oV+m1v23XKgvTNzFj8OiDy9vGwOkOu/vDCKVyDWzOE0J0nU7zdPMrn6fGaX
qd0h5Hgm4DjEOQ7G+PwJQ9rlkT644RsxwifEdaasmF8yz3T6Cgja8dCm/0oTVwTjHESJ46ebgbFO
RZ8CKeNL6oE4A+/nn+y4ly/fmBGPWX0+57mTzyIBzQ30YVO9MvlmRNVoDvzFbDeeviAltwMp9214
c3YCNk3cvmGyf1ltyntxt+p2zTkKCDJ1vTB006p40Yv/skulBvbLRD/fmMOkNaFGJhUYCS3x72GD
FxcRO5tCcZ83swt5TOicx49vOyhd7B3aqWW182edvMcDn2CaZ3ryMM2siwGMD5YnIa/ao9OyoNZO
om4bIHn/ew09NYjD5SpRVnlzYdvItd+ssiq3UsjpZOBi7PrsZ/OLUEqznBRWxz4JTRvMyobsvDYb
v0b6xURHhkhKRAaU2lWyiWXR+qVeAZ1PjO87MeM0sOi3DmIxKE2SxhuEAvSq7QSPb+a4D3OhHd5P
QuF2m/D7yrH7MDqNdPUUslKl6AlQ2bmqn9s1UBCQG6xJlMmTKjjwZ/sYh4tX7zz0z6ANXOm762J1
l+dh1bqYxrr4Qt5Jg/5A8tmu3ciOt97tiXObMsVCyOff37lgkYosABUsWTP1Ylfinsrraz7toRHJ
7ybWjfByNCnwmOx7VYKUmyD5QX1/nOqBgyGFRPu4ypv2qtTNtaY6KgdcKqElTkvaljDo6qQUzJn8
KWqi4McsAKHipl2RnQ6/+gAupIpojPq1XbG+CnX47Dyl3x22fhThdEjhwGW1tmVFYCE3csMaqfsR
oLQl3MPya+qFzpr/RqVjniS/N6BNiCbELOnqlboTErz2LGwpyDAtSm6nkcCYk70AHqcS9f79Cl/J
jEGgS4SAnYnXlNg/wE3ueiD+c5lKdvJTHMHvkzzDDxhERBwT2xignlh/aTgo1lUet11hunmYCLto
y5qxZFMf5bv1j9oFBtR0qHAoaqeJq1qwqQB3bNYmiuLAhWuTRgCniN4Y6CxgaVvCzSsUhlBEl5Z0
pOTU5gqWo2b1g4IkSDehqUii4LImb6HMr7c04z5Pf/fDfeTfiTfUlpi+dtkmuMKBhgZVy9p3eOoY
3sHD/pOQ+4sSVcPqF/67hQ558wsg3JaVTU6Zf+xxKB0QwvYdnciHq1eSY+hzJ7AWGKp1j+cmXOol
/nvyoJlnkpO/wBCMS4vN+ocQcObj9BIUsKIS4yYHreqk7LsFl5it1BL/soDor/voQmlCDFHJ8Bpt
9DCyCMARC2dnTv/Rm+qobQIhlzvH9OB9CiIupU4RFwstr/x8ulCgjUKTDfUxaooKl9Zbow9S4pKx
XX/qzYrdzBuyuAvnNorx94RF/Qn+h6wWTp0oxl6VRSTMfyAdsOZ8uZXkvQzrhWWIdHMHgkC1Cqfr
vtDXX9vDBLfAodqXuDSyvp8nuSC/ss3GnENdr4QavSBqEv+pFcC5VAB9l6OiXlnvkhXQNYwAe0Lb
Kcy/uBr5d6rMiwifU1tsB9G03/cl4q8WXderO4qUDv/GJTlXRRjejPouiLJgMPoepGfvIZEX9yVt
k50tSjcdjwYFN8IsTfA0MHX54oicPxZSNojG79/qk48ZlmRawN8RKQ9eNMRO1Ly6kjsZbwsA9xSW
tYJao2tSh9i+F6DwHPF1Hu2pWITcWVBdRTX4MIig+D2ln4+XOqehLqBCKLQG2LVI3NGXhVezIGcK
jFXfQcAHpT9djdZ+3dBNISqBJwnE/jQb35EL/ePfweSHl00xNMkazYootxDfGfQUUSgrUtp3zfg+
5D3qs7Naf8+wT4a5VJJrPForqeWzKX3HQOlfZWF1VKBmhlHSgjzq6bwsCQsLx16gV8T82C0yyuLp
E1hXmntJjCVIxbpkVL/Kq0jIHc3btgqPeBBcY3pCxVFxJ4i0EmoWCmjUU6nSANLMRVqK8Yd26W46
5KfFpVWShC83CyEzRxAQ2akfsH8aepsXdUtp8lSghga81cEXtdysHWo4CSOhnw/XOvIsHCn1aj72
U/X9MTDl3f6u7Pgra5fKhhSoads9vLmU0WemdFC7SJRYFhkoYxaCKTdQ8OzpiMjmufkM95gGH10Z
TCDOLyQ7/a6VUCe0aCQYrtrQEmd468UQSnqoTH1IXQ424Ff6QkDgosNGPs6Q9lipXnIshbMVYvuM
3Sf1SvRC5hHod2to/TrMJ0PU7F1aKPmyW7pwNJxava/Xg73Gr3dnWdzl9cOfPgMM5RlT70ezf+fZ
zcxdmoXUya5dUhFQNRkW5YpwU7lZwMADW8Ui2XxNf7nfe4hsdjg4RukwkRo1UlxnnQyvKedtFYrJ
3eK8t++XqkyKJ/iDZodXosCq/PF9DDKOIM4iRgwENx6llNYS/tiOMyjFYGEuCTDc/XplX9axfOto
/HcbGjfdMscmLL7SCWfv1VA6Jv7jXWCUwH4n6bN8KMIuRDrwnGftS8m9ViEzEGb49lNzZCbUNZb4
wjLnraXCgXOesqAUSrNRciB3423Lemrvcc9JSJONF3QlKKqtY8HPnjGGqO6v/aghi+S9uPq+vkTH
eWBMvmYmLkUJyaYBBQwKSZNoLDTYi/3x+ooiXGqbN3l5a+8Vm5BGty6uA87bAoVskXY5krJf7Piy
sLEgXK+CRLl0JC4od9phqyHIm+Pqp6CN/hcINeYlor6C8jdZPc/yZgDZwLn0PzOuc95hWeQlzucx
3T7SUTJxLRXg2N04zCFD4931kumqP40kWwZrYPkMxdENsZJE+MNeERe0tmjVZ9gpbU/AiMAWyJot
DhdO642Rwn//1xOAxEKkcgin1kSghd6jQPA0HGnYlIisCXV27A81n4cz/0S887WHTuxjPuFppSed
iHtcjKip7MeOxlkhB5cgqfnpiJsuu9csx4TTAK2E+0pRtWlG4ozfOtjvdl7ZHg+Ejjg2tJMrt+MT
Y7nCIdGjMzezctStVnRFRurGesXk/T4DBSZdAMy7DYgcz9aQ5DRZmzROZj/HuFQNvbF6RM/ZLbO5
J7bkG1nryTqZC9m6qn1gZh0RzPpAW/Bt9qvXWn7vB2MkMoraKUA5g29fnG8/NSefFIO84cu9ZCRV
QwOBy3lV3WgHFzlVU2ZqW0le+dbcYCbL7jFPpOFWghwQd1BmWjK6HzwwB1vn3lGHNyu2vLbSuxV2
jCCYgh3H8ZLyOWSX9ZBUOKi0YyqsbaCCyaLH/C4mppYPHtNDs2DsJ9MF+sZZ4+f1yvvN1Ca/WE1d
QRiXTnZsyl4bX8EcrvCfu8TcRMk/SOmlb8YYtZ6FtG7aX3LnnT7tkE4YL728ndl81riQAmUO/opI
lHU3FDSPou3CtJWVU61B2wdoe7/TWezBv9BgPTL978jPVV7qR3FDTGrf10iDHVpqQ8yy33yEfiU3
d/ZBYySkStGKi6HMl8NkwiApRvQZPEAvqW4h2lYgpQDB9H8LNWUvwUy0XJhbZ2r9t1zYmmfUx/KH
spxa6wc8NGLPdmRPo2q87vuLz9Vd6aEHP/xJbelB5iQ9eUCrZPLRGsNVIUKrtL6Kcp3uO6cIf0uz
KD39vSWg5HZ9N074BcjXRA230j0PDOwWEBxJS9+9ax1ljHv07QWUVMmKApEGC5Uc1hJ7Qaa2zHz3
fOzoT9z+u8Rx2sAKKEmRnPJzqI2DIn2OVzNpc42jonZhWBeJhKchY2Ba7AH9BSCV+p5d02VHbFyy
ednZIxBrBpMw+/Yox1spcw9GqsyUfULIdr2/dGqnmjE+VZbP6CW1lXjqRoGP9HPbzAUa1juGx0su
aCaszbPjHBKp8MPF3DTK40BUzAV720ix3adRL8K53q3MCr2pX6qAh4LxYylRkZsUUA3yoOKScNC9
mSH4MvhFl4gkiCFUCbYJNw28QnkEUesjdV2B7N4mbwMrVCeXT3KxZllhcJ71x76kj8bVITDxC4ej
saEgI3TEBqmyE6iPevoOyhGxFkH00hJQruxtA2bOVYVxAMv6gd1iYno+/z0V+5OrpHVJUcTh3qOw
/q+0t9hxSzUVU5m2ZPRX/z4zdQkzxRlwBaj/tPCy9QJb8ZYvjpw1NEX4GjevRkK5/5AYNFJ/7h6w
PSGheHbBotKzan30tTuH+4uhHR7CB2FhFTzN+kT/Z1ct/hCjaQ1BIbiw2UqySjh/GTQ0xcBpouPT
jS4CIdN+nGY+GWoJ1ajA8w93h5KPSQrWEqmoFi0BiExVujltt7Aooz8XVCVU8nbHAlAyF7/jw7go
o58UM/DQi1DKrwZlAJCLw0q6Rau4PbMR9wREiw0FYO+Y/Yq8gDilHUUnotUORzCeeGFFMEiG31rW
6lbtD+Ty31Bj+ETW+6KXJ7ysjzQbeNLYtlV/SXZkq1BXsjZ0lfZaUfb8CZIxQq8aySSrDu87ehr2
cU9mstGZG6KwRb7i1ewm0jJN7pOIZqsJzUJUycrhjMObXfRwUnYnsHUVkuL9a2eKk3ELEk3ZVy/N
//L1SFiwD4qBipTXO0yzmO/2aZu4VLtogOV+XvR5wXxyAJ9oT7aN5O93x31gCt81+8FOUv9MSXfy
rdfHBdGMsBUgVgCVBkLnQEeK30r1Tu+xaT/psE4Uo2wkolrD6aOmqJVZMvLZX5GBOjzRg7qyTkJr
tKJAItbepoRZ+htd5iOG3OYX6FsMGmWnCdBor7nDp/Q+qDiZ44QP2IROHRXti0Fo6fPdOQ556WPc
AkZFXtst4S56wMWX46ylcmCBrAa2v19D3JJldwjtrvt0LT9+ftCk2njSdDrEqdi1aIaISyL7pXGy
WKZQfJbaizCMTUeWI8FSP2qeDqQ/8Vu78baA2O2Kape5/ylwDHvzAP2BeAAW7cxewXO1jKqaSPyc
ontWyVT39L+iF2rriBqK5eXa431hmMMcyHRDKjs0cNPWdVnx3CXr77gkbpCw0DmAb7b9DtPi8/eA
2Q6bain7RTyqulmNSwjpQwPNrc8uAnKNYX98o0FNzIFemhVW8akvn4QVigsqFMfdELZ73vQI2tFo
5LgWMGubzzK6EgTmlEG3uc1yqyFHR8GiQzhChLtOehjkCvr3C4jfrEmKpqytUP8zidClNTERqJTP
CDobX4BkrEa4wk/+Z1MLtVsRnXNcLJlfYYJFYZo9xGcuqNwk1kvgAnW3DQKvW2O4stt+1HXJA2e/
YYeeq3pmeH7VHbWEyxJ7GdYtk+hb4gpsQCmcrlp5FuQOb+lAkZolmVFF9lt9qt2aGz+m5XEWJ/yw
bcKq0KY8SWs9Kz/WxwG9Kr86gIgTqHgq8XdbYYl7AXoEzq0lGus1aROjd628mAfI3bg12w2YTDcM
D40g+nLsjwvKOhPDo7UFL81+1ao9htYPEWS5DL/5N8nzbfCfmq8FkhL+AS46muKL32UaSaxTqk/i
DCFTRGzNofJDEvLq2z8iVknAlC5oV2OIHpj2Yp6knlJhzz5GzJGcImjLx4BG/KwxA0OeuaTgHmoq
zW9lD66fUby5Qp0yCMrl8LQM0MX7vDYEIn1MzN/uCbeU5zPleTj8g1TwhsMSwT6T05zNlYAQ8C/9
ahDU2I3er4wOYlMZhdhmtMgcEvse31lxN/PWV07ifiBLqJQu9yNKvwLj3yRYEJKX5ozpN+3p0Mnf
9jL6qV/lIVaccrONI69+EISMjU08/alCHXABpELzay3aRgNb4F88BEv4XwfC9ZZKaSSDgasVtUY+
uxmBuwvaunyFKe1v+PBB/CCaGItl9zL8XxZycyjX3UBLeHSa1SogdWavfBkLfzc2l81FV4FPCpom
WGT/wUWY9anKzdTT3MX0WHqeg+qqP8YZlB09NIuJ5nEK+ufqh9lWsDMWvXbB6j1Av9X2E9Y3tcSY
jMUQgFfdEc7vjLuYCCaefyNIXW2Bs63semv8b+sso69Wvfy2WNUSqaXn5oKfcJ7QD6NFiHT62dP0
h201ILSyXyta4xCyXcSOOpgmg2yIZH94Tvo8NoRS+pGeLj/a8RZiyxrF0ztx9Equ/tQqWVY8Sq+r
vN3BLcSsW3UnmSBLBwlJtf7wqtuCSnZsE+Rwb62c5xJcOBpM3/heUnBadqMGy5dokr44aOO49YUi
9ulUzKHgzBI6rmq6nQC7cEt2CMi/ToDBgJwIxgdk72jxC+/Wxm2sdXljBN0zBcsqYCYs7kySK5gH
iGIz6Im8g1a3K8Gl8aSixS6sUv4vxZ+cs1jE5IwvQykNl3Q5iCaZKkQw4WOVjQx2Vh39+9mP25rr
dRL9CCjZHgTBKofXQLEzZLWYnmR5EByOqHqUhdxqdwTtJftch8vzpojALmthhT2qPEj5kf/04DYT
xNCFZFq0BPeAARPDrKLrkPqu0JHlCOHka/vDHzsSh9gKC1V25Q1LMs9qXgONhwxPDb9yTW6MLyWw
tYuWA2od4W2xhWbtL7SxqzudPHLwY/SpH4s1fWnq/uEkB3UTcQE5wGYrYlsaLsLj5a4emJOPQW8Y
qKDpNK8K9PPM2QVXZxXD7qC7FFUsXb1e8phAqgftwRAS27HzIpE4+2YE1Fcj7hZY9ROHqPzw3nSu
QdfEWnPMX8ONjFs2/1qn0NlO58c7H3n5+4eLDJGsTnNw7n5/T6zVdj1VESfWIupTkK16YBmY51yM
zhXRM5RBFJIPr0+OYK7JiLwMf58Ptje3K1ABjW5hA6Ta0xRgB64z6FN01prBDNYWYh7jzHtf0VaM
5AmToPedjOo1fEXbGf7u2mnLrUsgitM5fIP5p0pulRB2pPG5A+6a35iD923YsrgCZpL6MvKkn7Cf
5nvwWFc57e4jSQ1odjtv/OK1W1CG3s3Dm4Mlxyp+8aJNW+6zFqk+d4/8cWVFZRWFc1iiFC/+mR/V
BlzzrHe2Oo0uhKdNaxZErX5Qv4As2SMDnECLbwN1WT0kmQrXcnmqXPoAd07eT5y0w+plVpkmmvmn
GoZdH1QqRNVizyT4/X1iKTtZzk3HaPOndWaN9gIF8eNavsEXBAwdZmKRlXhXrelp1AAx7hP8X2iV
bSZrMAX5QuCWgzZsO2l/8XS3U56PaEbtYUleg9HeScqGSrV+rrNadFsOeVCfLS2MK8ccLtHfPFq8
097KzyIyZ69KHr146CFeEaHyQFY6+4+KDOq1x0bJq9pP2QpN1W+7bugdqpE9XtuMwPa+tE9CcXtK
e3YqaWVa0Be20H9VOyOU86emVeuaU/Cv8+kqmsuN5w2ViWnVsSimlII0/RDFlGNUdf0CDjVZ04wj
B0qxnoVNQGtMwxF1UZVttfvb9NndAVpX9bAh2iMcUQh+4moO/HGkhmcJhtT2DyDmBiFCEC6kFJnP
tDhKnR/841xLeIHqYvPmGr/PtIApQjTUeYZJoosxlCVSW5ou21Q4JVUoPb+xq1tDxmjDarqs3dHm
0/krsyp8g1hscX8a2fb7lI4VrEEGd1IyKfCbkd30aADH+hf1Qbp6FXBQobsktjJCFIOtZC0nYJ80
xaxWUmXXrAV9U1fKp0pa1OxMGOGpHmSJtu3QIqc70Dqh/8OHdk44NBvCuAIGpJt2406RpIKDEmwg
oYNjThAVFEzprgH5OgcqKy9ymgbJpsdlHYTToFAq8aL049qT7w8gcmelkGlwxHIc24Rc2J6g8iEo
O1J3PM8Jc9r1KP2rKnhnKvmRHDvhx6F9bLqYv5QFBGh6aotwoj3WvT/lgfzE60SwjuJkNJABRlgH
UNTQgNM3S+eaCiwg4gp73v7Ky9yWPXypndvuTIfHYycqcpgavW7qMIiPDeI256vFV4w1uhkIdY4v
NSk+C6T3tKuidkApuTQ2jEUOKgqHqNpTXlGIGccDQqcdrvn/WMROKjuWUoYw2JDDMMl4sHoUb7zD
IiQPVxkSl7akRALtf8iLr4rTSf9TpGOZ/tfeaeyvn8mpMW1+mb1ywu12W5snvYGuRnkA24q40l3K
9Bn9+3Gl/WL2mcpATKRQvlrtK1kmNfHoHM6XHe31KF77xlopt3frSXbL7OUPVLq7gB6m0UbD+4va
fQKBx+TOP1Ou57LQ2e7M/2xd9168rqcjcVpXP4ZddAiu56i1lHl3XnA9aIlLApE9OHZyTqED2CCf
sEHLXjqpQ3BwtOd5ORkcdwQrGISVTWaqFZrSCpTrB9PWF2wZo4uD2o9HNV8UZe2XZcaKdzhWXJ2n
bMPfSvTX+P6Cul7yTuS7Icg9hNE2rXlffL3urWn+OFQUuGdEL6mVtCZZsEGSDO1pbVPdIrrDbmCI
H2qDc9VwwSSGo6hmltVg+/pczWPXXDj2PYmVXVGbsIy/2jjhJNAYS8o9zBxh04ci9pSvhR/fbpkF
LTNUyuWeR/N9SMKHr8DyDQFlXa1QwtRNUUjc/lZ40Su90PssAywR91uqOQly7o8PVDD08iM8cE03
xliGYlE2FBUBUAbd1KFvfMbGLJmbo7EWf0Yg01vidbT92biPVY+ll5uvCqSdvqqaiUYvawhPpvCS
L7x0MqhoAA4ZnY0EAgCfojUqW14vK7IVb55Bsa9MDzo5lQP9TlpZoCoE59mnSNKlrSWYe+O+S2Nh
/kBN1UvBxdVEghPc11ZOf6sEj0kt42WMJyTHIiSN64EHUYWgV4VEohrjju3ig/0GFJgFm5YeVQCp
+1OjDkmH3qUltIYqtATBv5Cb2Ii4z77PwTJZm5326R7i17T+AXNinv0h+dN6T5bDcpzb0q7hVdyP
jVafhvdnvtbbV3U5plq3hmjRnyHtfQg1z3eLLs04K3lOv8IQRk2tmyeYApJsBK7P7L9Uby4IVWKR
NHIsP3BJgwTqeQNywJDGg+kcYGrUZ/OXXSoyEKRZX6b+li+wllN5t+QfQhPA7ozXGRSarnhz27NH
0aFmARTVNNZFLe/bguilD2bIEH7Bk42OOqouRRNnrSBovLwFryXhnsZPy4ZgZoFTLy5sbq6Z7eOm
8QRqT2i1lvptToOk1NF+z9XRtpcF4jDN9RvlWXoBwmTmpRIeYoUId6qyfRuwXzE3cDtH4hQFIGbU
tePtqaOqBZkI3KuQQVMtHAJOfil5pQlxHzpryKuWmPLSXmf6iNrcvISDEHu2j1ceAuecR6MFv4dn
TqRQz8ImGHsu3Zj3haSF0gi9tVWWT9GaHTik+K7YP9wGE8VhhmSBOBWyugMShPaQyfaTm8FIs/e9
Cd4vZaSJTOlsVGkyfbR8jLz51KRQnLeDYI8r5y8014mDfj88sB9qbLTuCTWmdHTLLx92aMfRDpn8
zFj0SbLp1M+UCJjZ7f9+ar36WNk6gO5lCGWYJqMAQcJgsT1roLqjOBQHOqnsCvngbOxLNn3yl/+q
NvH50T0xz96B4Q6PEpw88ir4+i8RyjSefkORTRnN9AW1Mj7ofoY6unwGtx6cVcWVwt3JU4A1c+5x
LrSHNKBPDx+uev7UvtLqpoGdpHp5BlHFpphGpSoUHPMI3UowWFQPH8dYMO2/KJSm/4PR+fQIW9xC
zyIkS6FqaDgSxeJ1MUJUIObpZ0hYNe3o6lhhFq9Kk3mVp0eM/yJ0OZgcfVl6tNcijjxPWhfDSxL7
W+6tZDfEEqjIgt9Uti8D9xCMqmOLx7Q9rYYl//sJHx0xHUDPCiw0ersJCA2UKTQHo0Kp5cV5iyXr
s8x62ZKHgw0hHVuCRpXB0H07nmsB2EE0hCWEco2UIX0Z1r5eAcRDww+qs/vkLDnDw3pKDM9/+N33
2ubF9Ox6UIZIfmU0sljlY2Ek+m5cZH+rJb1pzPMUcLYGDxFlQF0qX+9zkXUJLWFVHmMhhGwxiXBd
8RX+P3D0WTbX5njq0toJDd0rVZgpZE3hy2Xeb4YQfhzaXUYZTwsesUYTDQuE9qZ0e5GQReWIwm/D
TOHx4jprdFryNjjVNJN6luMlgUwdW17pRv9vGjMoq4VrbW/HBBk0Xx1sXKmH0aXulb7u9qjfVtWG
6xLdi52HK/4cac6+mRVac26sjc/Zs2A4rgQcW9GPP0PPBufpl3lGBMF+HykzBIMKbgTilFiE4PX3
GOwDGI+sXoGzGq9BoUFQaMrC6TXGO9eF6ASB+WR2vggp3oD28KgaBRtrm/B/DFLGJP4MdQKir1da
Opb6znR/WN6QOTVzWa6sPw4m/nUHVdGOhI/Squn/urb0ioVREtuGWOmNQnCJETNRmbF9YHK6o/bH
/JIAORvcsusyDtIWVxQDFtYxylXITIg0z0kZblvhMz3U++uIlryXTwvs5fWs2RMc8PGeHzH8PYkk
QzbnW83AT3l52dEOxao833jNGurmzh2lMeJAckH+w2QUBDC+wynbGCFlXAaT1NiV5dgDXs7YQkAh
W/WpytcC4DLuE+Ujc4+udMjz3fr1cTVfYRxB6dtmYEz0LePcMokXVfwuEc/AXNHGnWeXufxN/rp+
/o7oUBTyHdJxKB0F8xBrv8cC0Xdpvur4VndzpC8jgyWxjyw6jpL7IBxPO99rP9l0gr1fNWj0P+2l
2dNypj37ezJ8BQ3TAmAf8hb0SNFxafBeZ/ozJNeGxPPpJIpF9tB+6Ac/X4zz+x4xi0+UgAWoYn+7
jDMTJ1vvR2n9jYcLLP1SrIpvPcXL4i7FXmobKY3GUrBSyfsaO9iLIHBGEc8esag4KBVvP7ZbzNL7
kpUqdzbWfblp9roMQG3K5sQsv2baL24DCRa+fSxfkdfCl5/mHstZjoTCF2J2Cdb5n/uzcXKkPCP1
au7QhVN3Bn0NBGfKJ7wuy0TejXdTqJPAmORBR1Hox4hR6vmTl3QVmUv+QVTv0upO7kme9IYJ6fyi
I8OqVUjtF7GVVZy75+XQcixOBiHEhRPyP1duG5GhMIqS8UGFVfly1NA4AUyuxvgxSrHe3Vw5/clw
mlbNJ72ph2a+eEdvEqHawwruxyUa2FJk2DtzxVBKLy86hWcF4VRNQxSJEgN0rF2vlv4/FFpZ9di4
MXd5KM0DuxBswiSnMfDkohimW3+cSV2jscK6YagbVsyvt9m0RDNQfz5PB/fPNpOGW6NpEUNHhQ+i
KSSoDgFagW7wgdCkX3cpU4E9R696eYLTQRKkX/Ae14isZ43WJq4HUP5tnWDiajcaAkexhKyJZyKT
YHFN6IzmpWx3Lbpj8cxT9kCbqUQHXTKvoBTVlx8OzYhrOki9kQPxf2kw6ePqX+ReRFJFdqlW2SAL
rqyVY3p/9QAVUvlxyf9CZAncN62TWwdpKRn//MR8Y/K2/qpomcCLpAXLfREIM2KVlXSPs2dP+413
nz753brt21SE2IGJEMPfKaM4koBLTZWP7o7xd2k9VTW5susg/tvMCk0TUQcFej1rfk27Oc8oxPIX
16o1MX3n9fRBwQU6HLLXeqlY1qHXzRklnMNqyTPGYqZXgIfDm2yGviuZoVs+i8m301jN7IH9Jvaj
qQnxiBnKw1klhbNk0cxlYtghmcIUNLmq7wytZDN14i//ILxrqLxzRsc29mAXnzt3wxii38Y4ek0y
5D4ZRJJOKrC6HLDJPh4XM59MjVX5TL7gLn0ypbLsMAOwAABJCQMb9zah45R+BG7FJ3yQyZc/URLH
syadvCsj+xe7q53JQva5wKvrVUOepnWupjshutOa9+8bHN5FyTbHAlVwk0kuyKjSPuDUlnPIVcDb
byslEmZZtTLJnjWlGQeb1Z4fkvWM39UpHMnCWhQdZ0DjezsSRQ86k2R1GgApFJnowmW1djVeBJXn
NINgjWDbX1UbYOlcs9faJ7H/KyuIZhiWp3LaCdzvSCVOaD0XHM7dFpD+cmxGlFAIADoTBSFUo+Ik
tnF71hcbzhPL8+Sy2hauxnQK3for146iCJ5aoEG06a/JM5AF3c5IRwT+Jld92Gj22crWah0Rib4D
4FrdHHGnFQtwJwcGA3J2gql9n0p8dELLXz1MTGP2mQKUc+qtM4eg5nu1bySH+SkQv9R496R1XCVE
3FRPK9vS14rNAqnVlk91nWySYHbLuTYkdsyVsjRPAjVJ0URVkgDwHm21G4qMXh0vt7XfwhfkAacW
OKMCM9jn+FfTnKBXVhE8jA/9xV9P4/dNoiKlina9YeDI9zFpV1WHpPl48sAcn3keI9FsbVss8Pbx
TRGCNDY4y9m9wwQz9Cc1HAJVzDXuI3agkZIyrE6vqYmUbsN/6nC7uy9MhRStKs9WhyMfh/4s8Uql
7cqCVqmaQTh0pg8xBaWMBetOaE2ZUaF/LTni/p1oNhANWNqkX2raWpoh1vyEWD2xWaFrVnQehewa
GsBQBXNtd+YjRQZ+JClFCAetPYe+LMHfBKLxP7ZToBufJK5ZBeMOciW7JFpyxqYNbQhc60MTSDK5
6KDYdTq0Nv9agELdi+dsoo0/+o5JXivls8jyPbz3SiUFhW/PVaJfi02nV11GQgS5OFikw+tmJwUB
AAcWljhd9jcO7Vb+CO/Xx+V4G0Wgm0lPwLM4vQdXBzMbx0agKdw+g9PmoYmMgelkrGaGAwk53RQQ
FLKTOxvaT8OrlXaauJphwNf46zu1gShac9QgNYLytnSsZYUzPMZxBNgWPptZ5gJRtiUi9yxBGJzS
nERqN1my8lVvBbO9bv0BdGGpqmR8Cc4+uNGDydbcrUuBqZlgLqX7zMtqV7B7YQemoMeHi16TafFj
Q0fU5LoEnaEAFU673cxnLw4FVTSBnYYHM6WhvqFw/81Oujxh/BT5SGyzOn1UrO/5Eys4g8MLAGmc
3RK1NxAEJywqBoX3Al70CiOsfyYcEkU8Kt4VYL+rzp8nAX9VA+So4w47X8DcGnZAQTXLQl361jfC
aoiTsGkAuh10x4Ogqu0sM+7aYsnFpZt6JK/wpwqlE0tuZQh9pvy9jc+HLoqvf5DWZAyyTosg6xfZ
CrEB8clGycNrXY4tZLpTQ8BR3L+tBp9MaJ9qwiBhK46NZCEYD221V4o4obZLuGGjSYQp3Ck29/uC
zCjncaIH6+9D/zBHD71TIkJWWuuuLQfY10PQsoKcebl8f2H+2m7o90m0FGVQvl66nkmL0grDFtRz
rcL7ealGplDsz3Qkc43doSxUv7UW721Z3tsBvK1RlPFa0fsvgspYtkm3nChGcpXvqOkxBjbH/MXw
YQA8w4YBqRBVFMPkIbsbD8TbeXzJryNBPpjNv3v8ZNK0dRRA637sfwmSYKcLrXzdTmK2nQEqqsWK
6AwYNpxR6P45nG1OTfTnPKSYQ8/fztaekRdubtRSucUu/2Owb74vlAxqK5Y6kR4Q2mLfhi0Evq5F
YQQPAabu5TtNlAp7ZSEG2kF0OVJ7C9mECw6FVPpFPOWU1geLuURDkFucOVBmA/WgeNwSAjR08oZp
S8VnSlmEtlcaNmzgYkFlC1VF/YuCvqi33ljWoWMAwolLjCZLH2ratltAjyLakKhR7+74/6PE5Tjb
wtaGsnUWBx7XEgncdVMcp9WoPV9SGnNFFnsdhJLpOzB55ueXrWJ2G7NTC0A17imo49pYKYSExY1g
sPJPgnt6tBWO3YBwdJoSf9sozf6H93YuqEGp4wqdfzQ5aUBgDf2ddxavYQtiJlC9NrTb531CJZ7e
Ov81KnFTD/CzD+lAag8TMWkRGwm8zf6EQArIKPxyc7bWKE+YCGb2edzTDMIbKybhcPuIy+JHU35H
/6dRhevLfISI8R3Oks6y9MrxvIHL6sable1QRa1cYBW4oHLoCsBDBStT7vVj7fHXiqWpZeYm2Wfx
LFCFC/yHPqHAa+K/B0YxXtJsDqpOzoKSESwOocVJ9wBGP2SHuxrS00qn6HWoYcuVZxE9Xf+o07Pf
ZVZRgXnbf2W6Gan/4AYqBkhR6xGtTlBoODgTMnhoHvxYu1LrbwLBARz+/YFLMCy4HUJagOzHIdkf
gYZWBDuFKlv5IzloHhJM6/RJgsIhp8jpHTdo34GiRMo8k6HTpck0eoo/fWWJZ5pByU8jahIJwp4s
EWDO1XMgScSg3vZ1EVidh+yuoCNnP9NXwXTNapB/IADMq7ewHLHku9eSsYQF5Mf3JRKhqHIbAWAa
UPpD+wv7ZVFDcEnIDtAW6suwoSL1UqAw7MCZkyYnbt+oDFJvhTcylbVgUFC/eWjHBZMehOLUuCE8
nxizhb9aRXeqidb6KTf3A3RfEq7HqDVhCyRA960hZbE/YM7AcSBnKeSyE5hu4+cyubUEiLdfKeyK
a7jwsxNdQKA5mwLhf26zeNq30wCN4xfxdkR2UY5tJApjQsPv/k7F6aItmJcLAiPofp3ROaxf2QNW
zOTjIK7ihXuqJdWiBlLQGO8PZYt7+FqXawMYD6cDKqx9NR1tP46iT8GxvF7Ek1Neq4CvZWq0ORRp
VYY3HU3qAHTrSEqnPsAPNHvAgF5bbAWBcaAmTCPvojTZw8VCLFzkRRT++6icT3hLNRIdB/Jk781e
p61hk/dcXm0J4fVj3aHlP12T0w8DGTaXxZ6lV19B9NSjbsAxvFSi2WBUUMAOvSjcKR2DStXWtCC/
5lJhCdUpY3v8YZQcXfkWxt1BQJggPx+SYOSHxpR4NZPD8YDvN8uunnYMCJqzjbmchutwRwlvNy4/
SB0mY/hnhQuNm1z/HcULwfr/SLGFLOlQ4t6Gy3YxpkRWIsa82fVMRZmS7nFiycmjIUk18gQdGrNU
OB8ieEQTHFBLiQjAFlbrAzSl6G8OPN7W3x1iSo1LaLkZ90XchqlH+tLsh/mRF5RaQd0rzigNh8tC
7g4JJu3IeOs0xlUHKlz7PV8Fzh0Xn1RRTrK2DaZkCBEzBS2YSisxR5hl/YXzBeFR1WR7+Krd7aGC
ot+9zYerJKGoQu4KWbBVQMfgc05CYLloxhEhY0sTmPsqMP09Ix8CnWFh76CH9SLBr2hZzoyEd/sb
2Nc1l/WJ8MgiSWorrIi4fl0qRaH2WFpaHpCw8ydo9v45gTIHEo+PdWjy37wMI7n0CL7k7MpHZeHp
IJY0bMAqyimWaD0o4DkVTpkFXUn/tUWq+9RvhQw5u5IS+B1zEI5tEqm3X9GydHbCoFT4Y5pcKKVu
2t2KdMAC7hLGp1pplRWFemwRx+80E+G/Mp+MOxQqDnpEdIfTZuNwE+n80Ur5YlS9pZtELbkF40so
lPGIvltmshk9dBNmW//Jx93josvZ6Fti1+ODyGF0FN+pdDwwzzye9N/Kht96vVL5OU2mgH5tvHWx
JwsByEQXePd3WTbEYqH9JxiX9YN5LcYwHFA9pVA6c/AL0WL/o26rA3BjVo59XQcVJqQUke8MdoFs
p1AEewSY22kTodqnWNjWd5CUk3wQC3gZDflpi8fQIfgEb8JTN7yB6gD5SLXS4ywV7AkC+nMwogBq
Y4vlFQ0xY0sQbPGexWFCLiiRuvywOLmQEd/No3jW7KQ6c93Ph3xkChA6TM9MuP+qG5mhBdkUttZw
knmcA/CZZUkw4KlQuAY2Qy40fdSQgg8H/RQTaUjT4iFBfsbONbdjO5T+h8I9MdN4yT5gcTLbQGob
vxVJXICenWK7o9OvGX9YkedzYo2o5tVqogldHfy69Bt4nMaONK7LyVcB4RL148fdwR28o+hZD78H
ioYEB+9937pzmhpZsf2rJdg0JkAhJyetS8URr06n7ddo/SioPtlJpRl4j0HQy8CVsDUHTVQxfbMC
lGujKeKThQqDQ9cLSGruktjfVq/SNxno6Op2GfrB3QyL//ltWiIuZXtliP3zQLgcQA86u6bQjzHz
K0l0ZSpEPqI/ZTxnFSouGgbE8XfglaIKY6/BBW0XfrzS7+q93bfsYiqQFYcru1JeB3Orh18aVgCd
Gwa3UMfBbce1BHbrqnBzHwh+bqK7QhAg4AiyYroTBT0c9ok2NeKxYUB/3u7BVxwjCqxyjsYjwrmN
wgyYVIPJjXaBQt9Mc5qH4dHEA/eTZ7QJ7+fFL9rgLvEBA2V9WJd7hOg3tWYCBrritrfODe8eNXsM
Vyv83bjhfqumwaAqPpzoDJkzGZpUkzx/hkUPsXoqDkPuWU1Wr+yIFOpVc97IxEpG2MUXGIO2lPxU
5nemtsPJQOqw2G/dL7f9P5M/MGjk/NaAKlJ34DV/XfkVliN0PNZUwrBgN1ZDw1j9Ogq+jXk+6mYL
4FCqWChMn1qs9e/c8l7pxCqMXh0H2d/qBtyYND52pbJGGc2cjDrUJrOhcsUzUZ8HYFGuwdnv48mI
yG1TPOIgid+t6ahZY+kqrXVr7icyVpwvvC35WnUYV6c0ssLC3va2CZm1f5Qj4g3l6Tpm5lnGqO0+
mW8ilfY5bfymj+nmOdDd3psSu65ZnjM47zn7JwaU0kB83NN2Iz0+Wf94Lb0CB49M0Q1QUw6I24XU
7R322kh11Lp8ZH+afxKQgPuwX/rVlsL+qU8TQlFfwSby9unCvD+pGdhNf6Gdmj+SscP8qZGASP1Y
2JnhFcN7V675WT/WPyJZc4mYmc/flu7SX+Xfzvx0gILw8J4Ymeb9eJzsQgOaU4ZkUIMr1fTfwrMi
hTEamzF21B2n8p1CK1veo4y7vQAWzQ0oizpr4EHFdrueBVp0pApCAQZatCOMLW/DNv7nNNzpJuM2
kbWX6mCrYiS9T/A5wrDzTDQibSI/LGig+iwAPTtB/mmmwpd35GkfsqOyLOCkIfMuyieHj4k3vhd1
ZhB9Yn+tTuKPkDyyHednS4U6V2ATR76JtqNxcjSV3b3ssiqVNU4aFYKH3SDp0cShj51IU6H/172k
kgvLU/PfZ8FudyeC9rrTtB1RArW9miQXnt83hJTKKgpeTo3ua3ciPWaPrum0uUypQfT3BkmwPREa
lrG+wKb0rseQoNvy7wm5EMBwZyWTuNbbWU76Z2L3HK0l+A12f5fztvHvj/4LJTWGYyuAQwuouO18
2T5CfN23cD/5xbnJKo167voLFU0Z1vcSlLP7sj0rc9kSVb+tj9GRTi7qaxOXRSwAF2hN62s8Rxww
WisjnTBE6OpgtEEGO8WvkR48/auWhDI4jtK0GITnisRCNY1TtFDevqyhS6jISMp0PFdmdAlRdYHq
GkfgdJcSickvX8XmkHsooUzU/dlML565TmR7WRSAF7YIw4ngpp83liX6PA+OZu5gkDe85hOW2Jft
HZyJ3jZYPaZ+tx29jzn3gPf9qslR/PXX1ZV7dTw0322B3tPE39UjSrZwVX3zfcuBV8jdSsIvLSGL
4iOzL/zizzS0hP/0KYNQhjkiY1F9vGBYK/RVCBiHyTxrPTQsg3JERgcVvOqPhYL4pbzPOXMVLKgu
wpzosQfpUOGV7fsVvqR+VZ6huV8LQgHRGJQc9L3g6KyacEUCybL8qy+p1EPAbnIbfuMQiSbwDf4w
DqPrjS5t5tpYCeNjUMJrPG6D0Qld36dK9XeWpxXZr2HY+GkZAQQSKCIMbWVErLsDPrDDV1LYZi6T
ML7WpvuQBgJxIj89jtS725vZ3wKiS0mbu17GJ9P3Lf9H9KAPdI98DLXGOM6CoZA3WjnDSgKM/4ws
c92HnCElMuhAAW0xqecd1V4CYLKI1elae6Tz/j3kcfWEP//zKNv1u02Tfvb235gex9INyW5PFF44
3BOwZryO0zP+k/4uo6wgq8dKeAMKSZ0lSw6HPr3MJ4F5oFl5SuE5wI1pM2aK9lgOSyqNk8bYcm1y
0RY2MSqFozWdP6kpccl67d/0tRzhA4r7Nbzfmilm6JIdCKp6AUsq2slkkcOeAhdNVU27v5+Pcqzt
tVlYfMtGq1eOLEodV9oBxLLHnj8WnmTyuPfhoG9B8bJgIe+q4VZ06M4YcL6mCjW+IrcMGIsASWxq
GHRfDnmU1o/2k8j6h3rF3xBgFPJT4cKyxsqVWxQ3OZzbDCeQdN0tYgt7QFmFDBV65kpkp1LQOgVT
oUexKiq/YA2B87pzOEHDZ7AvScLKTEi2yoyn2Koau51L7giME7C2lmsjEuPnkx2Nx+E2+3TriWg+
Xfh7SKaiPsf9+rGfRJUvKBItROAwlEpCso/pkJ7rku86yh0d5wxX/YHnE2r+7TP14vqiXa6uSoUS
qSJk6EkRq6QTTNZ7T8OnDs3LpPOLc0iymADrOEEi7QVgBj5opL4/skn8za49GjuDgXcdaZ3FHhPS
XqYxF27uZk29WoZ7YEFlP/aqOvspzyDdES+KT1uRvwm69QCHmZuWq+0Jov6KWHA4OQFUOaMzseR/
6D/oyWXafCN4S9enbCExz0SSCUqJRxk2XeJm5EjLYLboW/O1Vx4+2S+HQDRUq1INxVeQdvLKiaSi
ur7KIs1kBRa/wG4Z5r+GsWX+nNgXz3NnBr5V89Z7knh8KYC5yRZMBMRYq4AI1AyjZo90D7dXywQg
1odlTj9mZ+yR9srxlTxZ7QHbyyuBRa4X5/VFDganDBkUmkG/uEZhkZW6M6Z0Pn4UFM9A22WO1GHh
RCoK4Y/SHENRl11DrXCyGzlIHR1wbywy2Sw3FUdWvY9L/oygwm9Hh3yZsPxzo0x7qvZJlxyYzf19
rU5fkGFUQ3Qk1JAhEoYKw+/QStSARwkLxjdJ4yy9GCeDmvc0IQqCivq4MP9ma1EL7ZxMJgS0z6cr
ucTTOOyoUh9nP30J5Rfg4VuzzIFgiLA5PDatGd+i0ezTz8Y5cYUtSSzxcfoqdGaGovdXxIomsUkr
8ZIdX94KA+kafZnV6reIf0UpHeY8CuA8VWtnMDtuxzD6Sv5BVTkp9z7WSjLOI6D80anpaZAEbhUK
CQT8BYPpgArxogOu/aPzz0qdizCktC+Q96lxsD0eVHOGWXVfDOhxCVScyvoaOIbTMFU1u3XJ9Cj5
SBjQmbQsXyiG1YQ0rV3Q62JStuNpeqcg+ntnjIvHsavVmWW3JvnM7UQiTyIq/xLrOqxkEj13TlHb
f2Ub4/T+YJ+uU24jRZ/nyQE+n6JZkyD5hy+TwL1SAvK1qbA1Tyguuv0MxDwcukrZv9FbKxxD7MXW
Bu5a8Xh41cj/XwH7jE4cTuD99DihzM85JL/aEkl4vLjL7kI/uHW2GwCH+PBPk4gcMvte9uPOFGwg
ye+UtQNIPflT/mzAI3BvNJ6ddgcdj1aBCMsuZvmbzNtPY7IhQAXf5VckCbM3erirKpSeiKXeMGYr
6r4X+1fm7e/fguXHDpVCRQjhTigf3vKHBtY58oI+xH5UUQ0ay5jxPY7n6yMmP0Hl/ityTvH9snQ/
l7q6oSyHriKFNP/L1x/pgJohPFIZzXxy+H254+tsJxx5HUjPD2uZJliFRao59igrQvSmsMgiPBER
g+Ygr2UVpUEOTum9YLIIOY30Q6kSJHrY3EpBW2ae/QH2AQotoTpFKlJ+9Q/VwfUyYjBMOx1PA2Vj
TFo1pCpgewH5e5QZ/VYF9efpq+IiGJ9ZVKLZMfx/PVtmEKHUkNl4LS7HpLLFnxFU9kEG93Qc4aRw
ZrCyj53RZ7VKuIoJ2KnicK71KVjUKYUhn1ICd32iPqjCSAaas9aCSnVfYS9tBFhTgXohRWWo9y4T
BJNKdieNVnrmwLYRT87w938kneuHkBWLlB8IvKc+nRsJKHd/tvdVanMLZ/A/hA20oy3sXcAOD6Bk
0VhrCGak0X3oRaImsD2vdVoFmL9l8ZL0QRgC3OmPRoHi/iri/2ZKKF7iMCA6iUVgPnggobzcSbBb
SfzHML0f0kUN4gYlLzTpGg8MFMpWkwH6nstFF+YUQr5csHjqkpbsbI/U1SYdZyTUaxMClgknGv7u
dlx0KO9Pvw1lR1lqJt0IgnP3pS67OR2lb4xsYFnjQxcZnX09+zNHpI1Qo1wCkcrM4JWV1YWtCQyq
vSVjqNubr9121WA+8PFjZJr5l856ZGJFXZULfAKJkwecF0Q6b+AS4cgexTDTk/IuaV0iYWtWt5Or
owdq/bUhqR5xdqfQfIvACsVYUjr6TryAuMvX7DONP/ZQ9q7on7w63N+FQKLoxX0UgfNiV8hQRKoH
QCXzxdT4DkVvBt5zSVnN6xWMvAUaJyyUXcyEXxjsx41TPUu9ycAtXt1bwfaz5rb8a6XFik72+aEU
5SwjKNc9feFA81M0VdNiqWJG5hhU+xge8w+eMRDbkMvzK7cPFhT4vaPPGUG4A6nGmdawb9/iwaUT
V6pMXNxHp/Vx5S0S2GTKtl9aJ8nByHsi7u2jdsQwJr1Ah6jQKDlvpfh45SgQoOU2pEttNFj0QMVy
WGHwi1b3FzWFNLQjV0E3VNTslJgFoObSerKe5OuZyiSbTIVsxh4LsFgu8i1P4UlBKp+vS5Uon+HB
kdY1NjKR84NLPGz/MF+vD0s4Wyhtl8+dOOCjmKvHUY67mOLJGY3pv26sLYXG4FUpltYj1ufCLjJ2
TUH0G91OshY1bqcnwxRzpsNElq/QgwAhfd6028TnO/S+jE2HE4qbuYQeStWYJt9ZF3cFzdERDXD1
PImsUR1XSiRj02AQJ3KbPbTZLDo1+rxPlEKuFkSltVFMQeJ7VxuXc2s+mcKKRS+vmocMGyvm/2oa
Vxy3Sde8F6s5f/zOGv4A/ngOLiB0GFxEf7e3ZErt96DvmePbx0aSNMRaLP6kkUXzG5/6Q1GSzGc9
X9ViB7BI1J6jbPiONk42IBe8MOLaLxBWV6FoBNW5xYfv1ojlEppYtm4To//QcUstbTf4FCrWue+q
eG6yL0n2saJ8MPryW1MXkkVdcPphrlbiS6eOl15PczBNQX0OsAXju8tl7DEj12iqADqkxO4FCLof
JS03JLfQwTSR/OL0MGKMI5cpNs+LiJe1ZeIG3LHdQZtqCpIhOhh0KTMuRDO1aFmDBLzMP2y4PeWY
VKLbL9RID+GPb4E1t9KRNjKf3hZ+xF6/bhI6Vanh87vzAU95G0uJpC70k1HR1bVLrOOB9/sIVh7v
NozkQ36mUT47Bp+ADOAFZgv+6cE1TfblCS5Hm3kNbLvCBq4KFHGEzTxnPBHuyVmQjKEb4JVM/uKg
mdweMi8PQAJeT5BFxwF54N4LAf7pWQgvg/9YMds2PCnNI8rn61Jqu4Q8y0rORCBeirpZRncdvUQM
BT7WE6hdGkTBQoeo7PPURlF3UtbBq9uTq6X25dq50FWfCE1YmbH8QaUs7/QqCw6ErP7ICoF+9VxD
5s3S9S9x5HYKjWVnEiy562fk95t6oVbhb24yP5evvP+n5q5uYmwTFk+TEswY4uvzM2dFuchuEr+2
pC+/rfbPYRVc4+ndPQDV7Jn7z+aXHDwW3XD0XY1Ymf/2U3KxI1x0VLMYAwsVEtds/FCltlJJ5xAh
Fg0QXXeiYIsbrSZ1OpJ/SxWBDI4hFHJsQUY9OPUJZft/VVQPaHTnTr550R7uyjuy330ZQzJt/LUZ
RS78fPytcSLCc5s3dICdmgVIiXy/S8apbR3uYXrcB+Q9CLjV5PmYz+epXnuAYVsSNJafSTVFxGFa
h7rbaqhwJw/sHRhdytulhuFiXK5l0E3kQlRzJu23tMi2ZwSbyPmw0T0hmEDB/7iHBmvlNrBKu6nk
2zBfRR6Vfzk/YkT6ch0EYPKLkw0AtCegMg3VBDfTzplBSATdaDMA42fUzWBbLCjV51kwGQy5ygrK
p0mSUcmrJDTEqJXu3W/snM9FxrpGEpi7Y7Rwj3lniHL4pcx7T5K8QL0p2rpuwZ4HQIdmUdYKR2dI
o2n8OOQl/zBx0OEyCFdgENjLX3dfQYeNJWGw8X3SZxrgeuRM34B9Ssi+CLhfZZLCSlgWAZOd2yVh
NwHqxHJ+rwgdwagEKeodYkQ+LSB8jkQWBsd7wkvRp9/iXfhEWrp2x4hiL+YHyNn09e+4T052goSd
r5yZ+uiO9zL6tMxXCrgJ881QPP/JOMR5fhKaygt2MdJtFSfFiu44ZdNiG+zAGGpY7uIPiiHydF7A
zYR8SpRq991B4fzgAGi2RoI9cD5rH+bz8Nb1ryt5s314jjmLwVGjdb+9ZQpJh6XjpQOoiC6YOW1p
nKwbkKhBE/vlATOsqnHx+FjUMQbMWX/5+fdo+3d5DklVer0Zu0D0WqLHwNOh1AVFqx2SkN9SGAKg
Jn4gpXS+pfnZMBI46CFY69EU/5AlvIUSlgzS17ls3/SrPmMbsz9pAepVSwHE3LEJVzSV7sfltgZA
6RnO/hEivO63gOxatuAQFyOv/lM7GI8bzWC6YwtHEn/N64pejwx5lcbUx26RKhxIKo5nIdhdLzzM
8tYcg/RWMW/y2JPxvVAaNArNUv5vlXrfTIrikdw9G843t6THgm/zVq4EjW4Gw7aCd1T/pVww74VD
vfZI7TjonYTKN4/CCe7q87Lqf0Adm3+4iPAeg7hM4l0WeaBDrQyh6yeg2p6iDI7yThdZLe9gsP8p
ANtt9boKqaCcqoIZwX8o+cPdHUrDFVtU5ClXHfHFbfgljP5AqlP8y9mauAUQwSIz7T631CT/XEEY
rGwigRcU7YvRA4xTlXXjxldZE6gzaAA6CAW4z8Iq1V0hp/aPy3FsAtl1nhdNdeS+vdRF4ytPDg4y
i+wWLcL8gHm6wKW8cIiEoUVhrN0AXxVxPJ9rImQIEoGo9eR1JMFij7QNS8cZm98VCFAgNIVPbFiR
MwSI8Kar37rpIAf5BwPVpeV1XXxHMGPgQjfKrmIAQ6s6lvta4xPuLw1LIVapK6afcQONSjwk91V7
RGakH17nDMzC5Dea8NHZWkZQ+yp93//CR918b3pkCAEkAHb+6fWE/IM9ivgN3RXVJYSAM05cbEm+
5P+81FIoSJyjk1uK6+Me3kzVoZJYe8YGHKLwwcpuQFXCJ7kb9qLVC4yJdz2sv5v8/cuIIg+FGuWO
toRp9RWJy8UDnS2p+IEwAq2AxqpiDf2MYIz3oQ8IRxSRotTAq1Sv8GZSoCLPEA3nekJHoJLOJT5u
JLGvuM5H5dx4u0zbSejIjsDQeLRXkVR0RZ03mF8bXP2+bUlX+rej1AymLZf7pKzcycS43v/HU2Or
eNuRmfXH4myc1WdcSLvy+Q75KTqWjsePTCQzyEzbeq8fulkwVCbT+9doHpuvZZEQbXhOhDwAJbf1
aTuCu0NhZSvTvK0qmuIKaOsYbxrOGDG6UiTxmtGQn3tcTuYJT/JaV/QjQyvOF0AFFz+dk4kPM61u
o8trECWY3161XKfLKqGh2BpnDPPntJ1yN76BDw2SIVHYIogqZwcsdqziX/PyMVbikxFcZE5nnxr9
Y9wUBDt1cSjjjBGVtZtB0XoGEiMojj0l6rdbDfjg6HmHO4z/OVEQ7og1Q5EQ5CRku6V7pjwVFBJ6
jHKo3mUkpTleA5cRMcQZYiuvI0NRdxKDl6RPabcGnS0cPOemWPjUivuPVs5UHCpnDdnWaeuc6Rjl
kTztyR3v7LZWgp9ioFwuVALmyq70866asUWDL3yBzsztojq8l9Q4JPRI0UZNHLFyQYgblU3Y3Mgh
bilCpbpIZxtDhFMdUe8uosnODgDUSxXXmdJj2hyPJiJqee3Pl6EzqqtK6Ywrypdf466GFt7TGNoo
7mPY5vEVsK8LSB4Ouj4SXhSrNbRT/oqboO3ovJ0itbhnNi5l3aO3e1hKXLzn8fw+SDbudDSdd4Ms
Ge1A7E6n7I1LxMaOAoZX/atlU3QkfWb0VwHo6s3+GaZLKR2FfmBRGwU32Qx5fPMuPE+rS/2dL5+f
bINqaa0XaRGGmlTToz6scUqe6rTtjWOTsc2cTPMNlXodBOoOaYZ4DCS6zhms78/Fy0UrL5ApSDiK
wh63e3rnbJDDSnXH8eQmBWMy6oi86FpJY92w14/dDRbWCBXPEPGHP+EuJV5+YRykOAGiO3gHb4oq
ZluDWPVv8hFiQ3vBIoxR1Uay+j7f/YNz6bUWyFziWMnga7Lk+qxSFHdaGE2PnTQlS2Tk/VubjjT9
gCcIbg6xsO2wacvepC50x9NjXRE7CFyoqbSEWMvSncV297rucFba0qhLWHngKTyQvlKfgD4OawJo
+5IqFa1gz+b1phlFzQqmuoXda5usJpWWIbEdh/b2hWJwZXBFJM22LI5lER+0E6YU580vkhaY/rPO
CUSm9jtWqt1wBLZV52Afiq8J6iIcQPM+mUfalX9ZRZnzv0LJ3lmnSc0ToLO+7QWQa40RQWEEorpJ
55EighmpiVJBR9TLkrTAtEePC/bdLZ7pIUe+0KdrTaymPE/Bt0LYz+WvFYT2MXb9w8D7h0VjdDn6
hrYAl086sBy+aC7kZGS61mARIw2MGFYmfKRtC4bxJwPqHTgVLZSf6gD84moQKboZhs6isNu7TutY
928sNjxR9oshUqegqJ/+7FnFcQo1KzD06RrqI8x084j0NJJhOtHwpUwE2aES3Z7LwRoB5h7mzgcQ
Aw6o60zDBBo6Z7UQH5S19AmVW8OgcSY8sLhWGPnFTbz00nHFiDYDVDTx3i5L8t7dPKQXKlu2mAAx
BjctzKGOjRRfRXDvp5qPphAU6v7AVpSDRjTwqUkMjBq5SatteGsSSEXxJAEZcQp+yMixc4vtj9CE
MXgtFQt2RTbyj0er1dWPHUjeeHIc9gOjl3eAFegt9UxeLUnEpi0C5Q1bwDROJD4ynpHpvXUYEAMI
UV2FbRX5Kps/M2sWnjncUofvYPZyMGG04mokeH0aOeW9RPcRYocMASyioflHVoqZ6mXabWoy1EUF
b1ssHqymV19+j1Hisb3DLD1L9NG/2V68ivO2LrjlWdomXd2Kr6UMzk/y/5W8wuUu+gYvaJTW37ee
H4qTePyl5DH/79ZlOop6xnqWGHRjOGO6Nv9afRiJyHrsjt1Veu/73/Kp3v8tL9b8QT2cTtHxVjnM
ELGWvFTKtmNlnKsLfYofB/I9CUw3QWTyANPKASsgyYptKK9EdziHqh7jZvMAKR6XqYPRZ9E71i51
6Tej8xG2h9PSTaUXlbniclkK5YaijscJYfdPSite7TUcRAwB3DSU2UouaCPq3h48K0zb+f49j29N
bzZ8SVAS4oefr2UsCzVdBqgvjRWKczBaJNDNZeKvSn7Sp/a4L6Wy+dONhvkspkHgbm01iK60Pqqs
VhikmOZLrlQYGyuzoqiXi8xl8nx1pW/MBbR9eAKTK2sF+c00Gxit4Ii1ONYmEb03oUGBlZP5lL8H
9eDkUD7RlbqOFwrNcwdVBPw9ZzOOeOEP+zH18EQZY+nZQolC59Cti1w99dgO7Ottx2RHr/ZyaHG/
2agHLkdP4cGD/S29MqgJ1dnWDEtuxb5qjslR+JCcr3fjDKSyZASRzRh1EDvh39SrkTgaPyYEvLHz
DHVRDPaeZ7I3kSsbekbQlT/J0U88NHRTt05cXLtoNOdGR4keP/T8jjMBp2+CV+Dyq0Coui7jrflU
AsqCNI7zibh0kIixfEq4sbd9c6bbVQi0iYaGKvHVrF2DVMEaQv4I9OpLkpJKALqzlt4LkKDnTFEu
65oXAxggy2QGwboumvKIoPb4UWFcC7nreHQiLouhLEjHDpruae1Wvgqy9kzw2IcAX4hohHzlKlj2
Ykjg64vQa3vnkWSNFpCZKVzDpJDIiXk/9nrHoiBEqOMv+i2T15kfzCa6bMjJZXAdH6YzeI+PKiu0
fvmNeGyEzbf41WN+CQ3lv3tUX79xAZ3BKj1lMEyWc2DRuO4e5NxPC5aYMkRaNiy5h9k5BIbaMu0s
tCL9S1GK4olir698xmhqKvh7D5eg26AwUTbKe2yDp5jO7zcB5s9X42hmzrudLHncb3QkEi7CaJXX
50lZaHpkYfIlna5EjzrPipofeHTNeznwv7xyd354/x287orAsdlxhssJpnsJBS0IhXDzO1ZiEniq
23Ukwx8+x8LJtkE9XVnKdpbsM2p7WwxBXMIdLMlTdsoYPlJsh1m42ORywtpSbNxiAxGiIAL8ShTR
b5Z7xyWePyj4JEwGH/P6AjUVwCaQksgzRPMqaYJbUFnxsHq378OmscUFaDs/tbgpvghptUFW08RR
JPFASkqNpzu1tDLLNWZT1wolE5aedVeNf2P8Y1eysuWWR2JFF2c7TsACYuYavYc0irgZ9zyV7mek
B8bvvO2kDXDAxN7dwiEPtYL/lzv5chRc+NLRu9T2ozboX4fA3MIZCEQZuXLimCUKLGiRQEUUePqE
vE5t6dNB+2eISxsijJnFzwW6VkxWCsnQFp/SjSwh3YPiA+L6c3jyLRCMHtOZAfmVEbO1dBEpkO2p
WMaDHFzL9TVUtymKSY2trjgJkNOKGfFDwnE19RGz1x5vJl8bhT5V/bL3Yv9mSAv9vRqUpwSyD+AF
OG3jrmwUA3TKLgoePhKRY1HW/YbqqCvF3ek9U1DSB4cDdHlxDshYikmvnxkwMn9EFekLM/6JXVHU
it9JBDLjkVUh7J/CzEuX7H47NoACfeCMmD7l8PLTKlc4TxVIF8jK7mJBpzajGRjVzqDTKYxp6ePF
C6kTu+zIU7NM4gNeChlMXIjmTOzqfcX4T3N0ovbGJTUErSMwYW1uvShUAr6jkyGlN1tg2Ea+j5Qg
grRrjs41TJ5USuX9lXYTvC1FSuiM5r0xBl785W3RZOxuTwQBWXymzJdc07GYQ4xKbDqhyt0oe+9N
vROhoKdOZ1YGb0NzbFyexgUoFrbkcnCUpX0GZtwWDPVCTAKIr3QbDpTHpYmNLGJtlXnCWla7A0SH
FpWVdFiBkInhYZGp3ZHik3sEZBnfKDpvhrywu3EaIyssaDe9KFXFebkEEZTcwVofGYRTj/8aRM3o
JYtjCf143CynrNosrzo0OyC04yPTgYihMTTvl5jj3s0nyYj9HTpz5gLuj07w8vW+On4V1Bk+ZCGv
bc2UE9hc+NQBSamuwZjKpbjR7KV9hMrCVq2lVU3ecXUWzsFKc7xyrVWh1URGU8/BfkUz5qT5HTZb
u2L5AxnGnJRR1xGrZBgxwJLxR8YAOjpoDg1hemPWKhhO0eyDgYMa+PeVGKltauNVZLbm+flJKxdN
KNyV1dzpq1YnNmBHwlsyMAUMBpTmpjnhHTtnx36EV98SclRmQetkPxa4wdLfykK/FSCU0YkRCHmE
/1ZC2KU7LwazJAKQmnUAYH2kLyKBniRrqZ/IdpD5apBx08yCM+ax+fDOpxs+vMMG+w8g2R4TMIw3
gkjC/AdcUWmmeJyIJwvg97jLk//jKVU+lZusfZr1FiIstx1VfXx+UoWhXW/LEVkD7vZjDA1U6hFH
0itxUYlIBdPX+wZa5D2jzCCOxaubyLwV7BESJONwsoNXKIMr+DYWcQ0QXckTls6iGrNfbgB7tUf4
Rr0P+CaGgvubCoqoc3B3apYcDC6QnycYENr5VV5f/Nq4h904qCN3ByBmV9h1QPVRxC7IBmVg8nk/
judoDWnKo9WS+4kkiPfA7DmfAsTCu2rW6QV+KqDuyskaSFDFGMQTCW8wk1c7nUGClRXE0y0hSw4Q
9quvAXuN5WbuqweWcM9HGurpsJ0KN97O1PrFIXAduOMLlSutxMuhSXVT5UmjEFRmhCk8m8iGlYiV
RkkkwNwKkNFkTk6iJnqxGxUHQtcypDldqJgsKWAEf0NwtUeFky5y9kokYNBYR9J/uOe8Mysk9Hnv
a2KRVzAqiDYFJJJglduwbthybdqYjcMpp65gJBMY7BiJEZL8KHfVLZd8dRzW3mBqdCY8T0TWy/dT
HXQGk0Y7VhvYdWUhod5T7czWqKucEco8trW/5UwjGOrbNYipPk9daxaquG/KcFTfosB7TzyY0RZ0
Ex3eOIzVLjuQWMPYByi8hgo+ZM7o0/e8QBRHeQgBSBU2TPLTfO/D2OHFhuEFHYiwYi1jqeF8eZGx
3WXa3kTTxP0ZWA6ishxLhoqFtMXVDEmCqKgNZnIGX/SDiR8raPBSdxoO2KJgNp6ZNtsYGGYTes5m
sHyRfbrzKvFLnz/ZuOsSSfQhSUAFRFifY16TZNTzXywuvKZ9O6qtEIVPXQQXbekT/rP75XD2OoNG
rZcMec/3hHc5NGOxjMHF/zvOgTftzkCJx5VosGkZPEvAjaoEVioqWBwkt6UT6z0eUA8UmOmYujyA
rdIOXnqdp/gzJi+wIA9zeL3rh660Ps14zJJmDzpg2Pf5QfHIr19C4zT1RduHjSI0JshE1AT4fITq
uvIk8jhMdVJ1IcqyLyMfeuEnNR6KDzJsFCxoeke/aC8UMX8dBI/AEbRfNixb+DVvRMcU0qBG+C65
4vlyymN4dsVX6hRO0T+t4ZD4u9JjMDOrRzK9pM6b/PlReOMq/AYILl1YrL6ESjUqt1Lifps9vcWv
ORN1BEUg7JsGhy7RyK/Hx7SeNCFToHayzOUgiavObqTrY66eBkxZ/qHF945YvxIVw4uimnhoNkdb
BJ2HBVrPCS3aHKaohpkhvGMNTWKuXB6KrhMGNic+M48Yu62b54zI5FyyRYyArXEEY77lE5L1Tg8V
HbsOJ6YTmm1CaBxE8cg7TLA6weaQdkQiC1luJkqcs/PFqBgLzJSipqvm81Kw2mfX0znrDa99tW21
2GdzQaSUbsqfPnbQbPLJeDoGccyiCEy8XQfVvbET+K8AKls87LcACxuRsTrKMOsH+VhIgfkurgA8
aC8xDtnuj9jopwjakWqGf7yCeikmtyb1fOvrgzdFGONgksDndYY9mVtvqfr2WnxTlizVJ45P7paj
JSWuPmmzEIGLsJvVfMSBMFQqCyyZdJHZU5rs59bCcHm3anQsrg955r0tWba05lUCtM9zOzOSeY4H
KNqM2yjyDDwDnBm0a33ygiCQO/cNctIBh4CSeXF7DSDzph4Cd+HLWmitE3MLc2pJelxuDAP3QxiC
IRjiKrFSBOJ0Vhq8NciniamzK3dzEDcQRw+HfbCdQ5dVwNFnH3Lyn+IXcALuU2WODKdor1gc9zJg
zi3DCDzcrIdQ2sWUIbYKMgf7nhFcXnolfer4pH4XifcRYGMZbaLDo2JLPo3+H/NS+//loiKHkWVB
ftQ/t7mCk2ATAbooKYmut4De5CIQSCCJFo+PtEc4UkHTk5n/ukeefPKEEEwQoroCUq4evbERzwJ+
jBfv886ZXuPqJ5A3qrdxazdG+kquId8SHWvGRYJoe0iwPS+UcSZ9m54TmJN6nAXRVcnmG6TY6z1H
tB6++e6hIW4rbKcuCb0Sykd0C93DLjhVKpoqkVZvRmTMkhk77cqIxeI9Ixt4A74ABh+zURd2/cJH
TrpOcoSOLx98wuhrWMJAchUUXp55/R4Oscownx9szehwTw7QQhFRxJ/cF2bqM5w7f8hEKpD5L7o2
0z4F13C89kAaShoW/o/rDv7+KMCggQ9TBcahTBRGVUEdCWY8+cq+T+V6zbBda4zUWZjvTPzxJj5z
7LPhnbje9+mm3MlTzyRxa5qDotIFH9N9x8xn7EFUpI4QusmmmLpRh9BoV/9bLWebr7FGTuJWVScv
/iKL/sMA5nY2b3MOAYRl4KTWt37RFhMznLPeQP/k4fe+iXWKj5zdtbMSaRx7lr8AeZ6RHvNbcI0P
pZV9bxqS82TZrcLt00aC4UCPfx2mU8wBAbLVzSfaiF7dU2qBZyLggR0VnN6VWX9TiZgm0bSi9vUM
0oSGdGB0Xn2SYoRW2mHnDKNFbXKaIXi6cRArAVwaa1eBGgr//ldYlXRIsjCE/YjyRyozZcUfg8OE
BkqXVY0QBX9Y7p+4Q8rqRhH5Vf0L+VxTr/wfjqoDhXwK5sPxGL8qpSMraI71okuFzOgDdZH+CNW0
0pD3mA0gX0s4yzj4Bbok9lCqJrQo5jvYANNnV0wbXDcP688EhTqQusnLS+3YN9iDv8IzPPpYBX9P
ZTawE1Qi1EnIB/OnudB7Wo7C4mxK13mhvg0RADrNz23QK+x/oDCiQGxjIpdh+2EszMa78ZXZNiEl
3k62M+7BjpeRuD6jw0pX1w5eKxhWvSanb2OPSjxOg7rV8XWph5dsA29Ky7DonRZvixGm3S1bO5ML
WJwV3CAQudCaQKMIS3ixsh891KGB0bstPrSJWpF8S+91/CfERfguu8utcVW50Ws8wDk4FLO+bdIU
sThdztSDxbKOHQlfszBuSfHKwVCAIy24RjDO58IjuBF1uZ7XQRCtGjOTOd9A/kFzs+vujNWGJrNS
1w0VTeScSDwCHfwPXFp0Mx/lhWSdXJ19m70p39y+OkMKyiZ8i10pNn2B+8wW2uO1WDen5K38oNzQ
4XvV8LxmbNxyC3XUr38RePmWdIvzH2t7dSQdAbw/zP5B+fb2Wqi3FCP5doYRzWdy3deQ7cpaavmv
gnFKceXtfYCOPwKy3xAGEpspUOXklaPpb82AZfkBGppnjQosMZQqbVcfX//dAdE/CSrNUEICutib
frHXjsxaiSSgyU/7YO3UZ57nzTtTu3UXTrRgP5v6QOyDfC858BHA/omEpZ/6VIB2km26yJ/QjNA7
ZhQ3hnpQJSQ6NggdwXl37OGtzlqOvcEP6WN2R3JRRv/fLwpr/OS30cBFm7LlTfixr7yzcS7Yd/qy
5z1Zin48/p5zbJcXCkeS/J7TM3VjBfyGSFRIzFRsdsTdiNieJtFV8kau6AI1xaiZ76jqelHSE4x8
SH2ZHR+ZCOJmHwAh2X5DaZc642DtBt8CxZvUb25LjQ3XOFfeT4uNwjOpAfHuSTHy8SxgoQl18hTy
eTa+UOGsRxwe5Qmx0A8tZcfv0F6fE0WNJkHwUhudPDPsqfODpOaOZaHx3xfkH4GrDk2LOSiPrGk/
lE2Hzz179SJZIa1kKrxgHv5DYTPpv334GZaLvjXtCZI5kZEHDtdZlhXo34Ys13INLurGJ0ubkS0m
/O8ncVwK1D1qNH/IEv5axzHitbNIcXIts2/Ktvl9/emzoEDYwhiu07NhUjFSPq0A0v1bcpE9o2mS
ut/LwL+ywQkvN8q1/NUkD1JLmtNxSehbVYcYToJSisii6RcNM6fTcFI9ZdxxunA9BgITntomrnsJ
nmFnK3ZrFRFFCiDvaOgMjSGjgYWLOqLJOxVu6WEy9l/9G0ojQefLK8d/dwmEnDMofKu0PVBwXuuN
REaPrwVEPbPC5Snn6PNpWt0DIg82ZlTYW6ze0adkKanMQy5Y0rg4kAiVl3gaaWEg+02FQZPdc6bZ
/mYhKS9MtJDiAlCJ2pxpLTIX6PO7nye5DX23Pf+PpQVHWg8falY7TDxm7hveDAlZ1QaU7WYk8J/2
NgLV2CFTmpUlr9bjyXChDXE4BzPD+QLnUX2e0aXM1fbING/JMMFNsLH6ghvgUgl44YBH7+/YaBZn
Hjj7LLmsY/Ru+7tnG+/I1GA6QmK6sZYVmfK2zmMuqkO3v8nVDDT8w87S7IsOM+Zkkl8i5YVB6rH5
SNsjXI5t+RMermsib1cxaQqcp91vcxLvVaKqjDWAnCUWNkZrzWvNIIsGeMIGQXBXSNY4qXjHubKF
s4x+cbPjUe9NmiMXNGyi7yEQCaKQz8TzZG9y1OxZs9+BwxLMB/ENrVNEp4mDp9gvQ2mJg6TMMa19
+3DMLpgsu0P7408vmA80XXo8sKtGFOQYbsccZbL+XA9J+Xfp3Dkw27ml/6cG4ORXEI3tWY90Ewxm
vt89MeMsW9a/lq+KNjuAOAz134BagyfgdK3/d2F4lgGntOSswt2a+6NkalgH/+z8Z+wU3WiRsYIv
pOszHQafoePnYnwYxUPLE8YralAxfRtnlNclYUKWK3/jdKA6iZKkFfXhGQSrIvhkQOTd9qFfSe4e
HNocBAp1WO9DgannjkD5/gch+g8hpyVwG3bKio3zBPDyrwlYqFtuM/oOg8KhtuadYj8sXCRNhLVO
n9KrlqzeE697FcmtUqhHhbIqTaNDX3ojfFD+2pR2tydGch7lnQAFe7Xq4Lwjn2NlwvkhXGfMEEvC
Qmal0hjQh7LGpyJCMpOK3pNbF+SQ1Z+ytzVNcudwxj0uib8VzPrqO6RpDq8bxE9hBBdkN57MILdB
CBoUiq+0sOGVnwn60wYk22tkCGMe147tcLJCjMhwa6/z9o0okVmsk4iyCXqd+sxMRsQzC9cH1eMu
Z/X7HR5vnNG0D5ZkSp3OibCEfQW9UGrmOn0KrJCay9vkzDRRzI0DkNq3lIpLfipi/ExTz7U1Jt4a
o6jslGGz+yJYVklwNuPJSy9UNf0/vOuJ3KZ4vJm/jnRi44q8zypo1UNGfHPAbfmb57JqZMz/5Y+s
gu5zBZgfBaC1ngrUzBn/A6WQK9qXZs9qY6vXR6+OJeb2ok2uUNPFuHsH3vht4JuBxigplDyJ3CJK
2TAo9Ya1tVKbnLlZ1X4YnTaFkYsDLbihsbfO2Aja52TfjpSULr57fDbq5gbXfaj5sr3JO9XYINo0
sf/jgr5vF5Za3RV3Iqqrw1dBE4efpOqw4o+JO3sXBkOyvOpGfWI+NBTwRBYJdEK0w9inAMaSg1m7
BOVyk8fXX6n00yFCt0dStiJoPB4q/aprUSFfCHMkO763zLfWernxiqInF2jjqPvSYYnjTbtojVye
bl2OXIQ4cXYP1LYQmrVbok/GNQ0UbkTWvofCQlsGveSppknh+MV4jA7pvp0JDygAnavnG2LmXVRR
ILXeEmKu90RBU6PaNoCgjf/oR0wMOtLhDKL5QcTyHukp5P6J37LVfxhWUcitBcjBr1mR5szda4O6
wvbO+z7XZdgLIvl4Y1GT5vGvHQML/U1oJzRTbzz/d7b0Pq6ccaXp2paNSnCVCLxKaPMqRkyf0dVS
tBBKDhGGxpLyv/rPLkr3GiiG7vkXdEurntr0iYhTpnRrf0O0rQIr/u/IEkftD62IdEQLivez0Gp3
J8z964Ufbx7N8TIHbsi+55FQbsYte0XPoNCAM+bHpMY3je7lUMCDOvNeSOOnXzutZg28w5CoqULW
JU/XTJ5kZBH446LhbpqEfAshSTQUTUhvbtFExkZ/35jN1hSbfvBp9v07F2DbkH0uKRM4cLqU14tJ
S7KARl4LGK9qkK0xM1r/AZTKEkfNO1M9/lp6DrNeHOVtIilKqQf1G9ao90MxoJlt9xRMhtxehESO
bm/qIUYlBnCfIy63G0nxMRsA6qInx2C7v81LD/cTolDvBcmtEcq87RUATtr/TfioD4iF7GoXfvPs
zBlj3/I18VrxoexIqxo9jl+fBfBZOhcCA0+H18r35QHmsYu67lAu/kq7/Cubg4bzKQvcwcQthcII
3aQtaIl1hkYQsWDitMl4c8hapWmMHZphFby/1+4SKWxmQnrzWeRKExM9NlK4sZ6d1N0PzJbkTLhA
wE1ZIt0ePVxGz25Gxl9ooEe0jWeUsmjl0A0q8Zkscm0Ia+bnGGb2haEhcVprZzjOzSch7/hedwEq
mAzyBjF8iOfZXwqDQHFuF15kjrGv+sn6Ri0TBDgi6pZG56xkikKhI69ouQCLrKm0OVBeQZzWcb0f
N3oEheDunm7Dq/sH65fHgzufX4GOxG96BtJ3XqKHPm/LtAESrUtmfOw38RSFz8dQn5Xt77S6k7tS
dXNLqz9xR+pVu2cN6yXWzH6J5qihveZMuxRuP3qa1o04aQIAW3MVCQbz1QQwJklRDKxYlJF2Sn/i
wb8T2zpFOLZesMupTCjCVuoWYE+DOLRDQjgD9lyI9NyiX3eDY8pOo5rferURYzZnGPpMVZJWbqcz
JI1xGJhgiwqdqHIO6O8qCGtl9qM0oquDM6x3BFm+IVCyYTVcA6ZpZti1FMtgB1JFOBBq47Vf4F3w
KL+nGvWk2XeQgB4ue5r/Ns+X3dU4Q9tD23UVjGmuoHUkoVSp3Q0B+jgj4RgOmDdIicTyXmfQF8N9
RnLm9/ZoK/hVZUjCRqu2dRgzbvY5lTiDo8NrJxMWcTbPRq5u5Te6zJVhanbyl6wsLvea5FNac4GF
StVjDh2nmZm3N2Z400474Ez0KCZABaIogpClpOwg4uONcqKaszcodeUxiQYV/S86U2CFBGAPW8A+
4wssBSRhC72hRKEEObAVkhTH1+5I0wnmdEBuJudJeym/t0CKAUNYP6RhYHbaXJ/ajr/kCvBB6ryE
wBw3p0+J3Rq8siQj2jjU83KDgQix6fDbHsvk/nBbF9LmsfVCItw30Nx6kFTgGU8VPtp1BUEQ26MP
wCfHhpHzJr73Pkbkn7MtsHM7vswO0Vbd80yC5UcUL+ntAmWHN0PQ2AbLFxtGUFeiucg78HLb4s3d
16Ve5UEzLjg7+E6og4TmgL86ABpkOG65IomwcL8AF9u+0l7dL1O20ph/AdDUbAzkboxZ4lIz9tU6
kU1NBsatWuaUDk0jD3uNTWZuR5LBYlnJo1u+6VBt+SCGMR+ZGjisWPxlOE9x4VZn8K8fLh1KqukG
tYABTcKC91/I+076Qzy0RM9tgcxA2aXkNPxdV5dvyfsYNxlwgVs5zXCSmqp1s0IJN8NFWe8t8tld
/rrR3Uo6ceDijTT3LJGXM9R3DYdnrfBRUmFaa6pCDACxc0VjK1jkwTe1YXWyr19P2/b41XA5H9eB
hITv4jDAFIuOPw40qdO8P/qTPs97NHpF1ryhip8fpJKLCiCkgn1qJG0HWOIwisxgtTcSgO1JbH3Z
npIy6Oh7B1gF3Egpwqjs3U8kDSnjGDrkHTwumPzw0KOkABLwED2gMbacoehNod9T5kKubjh1R1Hx
+6stg8S32KsT6hxBGG3FFeA80E35VAYr0ltriWRoS0cYCjstatxotHIfFHjSN/Z/c4fLkhMgFmMj
SWLF6Kn83Xthz3eFeykJDEYdY5K9Kb5zsm8TVw5BBB/TAKt332AQmB1lFfhD8NZX4c6VpZplc3si
JjWmkOIDv2Kseei2hoZltFvIBW/GHtvLRchqRe/2Sdl1gAIsKAZMfQxjwcaqbGtoP6YIml2Ih6zd
taf+yugHjual0lCKi5glfK6zIFk/BIN6+WoKAaeWUEk+lhC8V8OI0JGk3c+258S5aNU0CmTGpxB7
+AdRfNs8PcLgkVAdiwz+h2v4lIxXrHO1nXy/geuMY3ydJTbngFqi6n38UbUB2yyDaxSnmmndHHRi
4pRSYFy9daRGndfSFIe2KKpbQxaQ3KO8KKhcXvIwXbLo8i0HJMLxD9K+jgCG+5KgRH153gMV6BDX
G5nxyzblgTocfljT7/oYG2UYJXQ/5PpxmN/YhYdHFavGypX1DA/eKal/vMYnIwEQCkPLswn5qJ/i
SN/+PJcdzeHCuXH5MfLOr1apIgFes0O7lJJE2J9Wo2SOZ4EW6baH/zPZKi+hIHVlhMLWARj6PIor
ILSRyOjf33aQOczSIgW4U53eaD2eF77tKQ8TlTmqIgqHKdZDd4v/KSZmPRWjC+DurbOIuZFfKW7n
iqOZj5MGm2kmb4lkOQs+iaTH/rBU8Vy+QJ09QPNQvvOcrnETdk9iIKx2sNY08d2wGOcwPEEXKRfp
HPYnlP59Q2x8sne+uuJA3sdafTg30EXH3y9K72dSDMHrhxzrVOpq6q75HhB2q8h+DnGqBciB/jVT
/01Mx2etK9L+SrRZZVzEfgmg7UT1RsJ+pad8peAAvSNUDXzK8kbKZtJk0TlEPgRPMVodQqIFy7cC
Mf0Ho0uOp6fQyauKohxeZ00CMN9+SPKkroJ1KuJvR6uaHs1Kyd6EyvutbLUetumeFB/vZyjw6TO/
cGhM/CUlhyuWwThVzMVmx9IvXqGfYCC4FbYFCgIiN4FRifyGMvwKK/oJIugeLw5kBfpqz5LKP/xA
o6MEDdqmBp8hDZ6YImhlHyFNLc4iEBD9ezM4t9uVlXJgcXmmw8kT5tdCMFS+imxVhzBb/nUlV4SR
kOARUK7BloDkbBuR8P8nTxxZ5I6DTZKtVe3rW8zwEgjRvRG4IIDm1IK6ZFrfT9XvzbmDtihzblOi
AoAVqdN+OXnOYYWZ32JC5zi2/ZaKtPIP2mO69CZkq+C5POIBMuOhZaIEeTf+J1Yn5sSPpoJO+e7T
hJxON8HMCYcU07RmjcunAojh6+qHnRUu14bJ0yzZ2HALEm15ZvIOWKs1GleRkm61m862nenijrdr
c6t8ppBnvzdFm7Wb5BA+/6qXCdYb/eqKvkQDA9EcSpgkxdKmYrP50l1aGNBlFBMNW7Th82HnLuEZ
VOfurA0mNtt5mom3JuTWgGtV2kDnaq1ZntEC6qSQqrQ6+SxH6cdKcMQGI9LEh5VIPQsJjx9dm7oI
uzGQcm0p7ri5bonOETwNOKye1lASFa3QS0lT3DSRKAdRl/jCl5+l+5m2JVwujfhwgRQZL2PrGVsO
vuuN0PYPbNvAq8YEZxQ1SVNbP6Tce4AUYOgzxyOGChyqCY5wfB35nAqUvDaRO62dBCp7CuBjCBBc
blxLkaPgxYxTxvTcCtEtiT9dxjhZmD6b/zeu0xL1DfTs3ja9rxKZrLAt9VzETcTRhX8j21yN1wCf
EIhrS3od1qliEBjd60vjpx9xY6sQhbyh6J1F3mlaw3NeFZOsArdseuPXyQtdixicEboqbvekgaiv
wh8yxg3+ijP65kbbIn/SuaZFnmPxNZfV+cR1PQwdfZQEEwFbN4J8jGs0LbrE0IZl764rBAw/ZbBx
3kwvZSCNkpLthb7rTuaLQBDeC04sBgjH23wTZFwzXzTx8VaEQ96hccQlb1DEEFKnu1HRk8YeFZG6
GRViUssD6iqo8MxhenSY4ojn5xIss9qnc4Y9gLkD9QbITDNNBT/T37p7haCwHfA+2ph0YwIZn4Mj
F+PhjS3UpSiN980MV5XpVIWEyIGdIiedwnYBte93b1Z0r/Lx+Gg9NKIfPi4En8MNistjtf+x/3Em
+G1IMw11UdFIn8aRU/H9G4Km7D1mDcjvgKbKb7E3urX7bAZz5yPczxbB2MnyYXMhOwjQbv/4AJg+
iPThyDG1io15QAWV4prL7RkJrEsNw2iLSPUMlRClJ5fRkyxdQPUaCMCQ9NO4nrWy8l+PSqRM2jMO
UNhxiVlkVC9ZbdOAhhl1n7dJ74+AVfeaHCG14Od4GuW02iPqMx10Lw5hxUg/7Nd6EYwSXfbOgmWA
fIEBJBl5Io5ByZ34TCqwQeU72PpGWk2KjQWXYlUB8eeD1Deib7hWlwFRRLPivZxFJZnBLLHqMbp+
0M1Bb7xPYp5/HaIjB1+ulurr4N+w6m/uMKrtJtXWO9C0z0u7vMCQdf8ak3UqpTzSpxeqmPd5h1h6
F35E1C8SQnazrjTRy1MVDX/Z3PgP5/PV2xeiWurHenoGw7SOL5IgkL50Gk0yhFT3Va1Lh1dToQzP
4UD4pmPl/qjuOEMZgbthSubBQaAt4Gf4eKcXjkGVFie6/8cqf6HdV5Bkh4SbXU2qweN9erRQ4G29
MnKGjk7c4tQjomdPD+UtsgKYNqeP4XdZa4hE7AlJKmEGBxxSIxFhRgKeAObXV3EPl3GZMDvoEiiK
i6zeQgu/jytCpp9FIyHZJm7Dsal+xT/An+Ipw183vAPCV2lhvz2AoQW4LOgdi3teIuxKs5xiYpkm
lvGuVYPY494D5PyskN2RrAJxiIKKHojpYJ4bNZJUqXM7Uc9BrMUKcQCjBxLv7QrCPI+1i30M5GSO
ChmynT8OpFfNB1GR35AOrY5m62GRSrYeftqUtnO9nMevX1W/nyU+bfFwFOR5AIR+h1rdFJ0ofpBn
/qYsI8Rxs+604vVedq+it9EMzopnMqbUsraIIYbo6DRzOrtdwwFgOTBI1P9IC4hApKAWt8TLOOpX
/vLHk03DywIv+nITsBK6f1ej717K79VHn2u+wEMN8+N+QAKGwQ0fT6ETEEVdn/bzjjjPQTa95mH3
a6oHPiZEoStPc84zbcRro+5KC8lugIl8eDHHV+OXEc3rIoSjrt6FExeIhhEcQFQ8TJ1S2WkDAHt5
MaJTyh/u2E+E29Le0FiDJavjmg/s7zuao4oA07LSCD2P/WtsHrKL7zWS51+XRiIP3rZ5ju0SoBAN
O6X48OLVhStq+snUcAsB9PEejG+WQJf1hUPiSCIZrXWFRHzX0otjrflnSCO6fkRFuLZMFD6IdCkc
TK9sFtULSjFFMbBpW/NqFUcwTpwkgSocl9k2MRVJpt349WMpIR6ytX+GHvRdlyeCGAkZ/wqRHuyi
2lYzgAB8FSuWujAlOmag32rr2GIsz1ZgImbab+Bzj20eYfBAQWGDXB03i7VKIl8zC81nmz7Xv2Rr
PTkmEXzlrUxXWSISeZw0errj37y7Mf/tKEslfBPk8LAzNF9Kq16Nb1dEn++p3dfOF1t/o6S2qX6U
cCb8mUfXt2IeNZ4NY068Viw2HszBhGo6cuc6CHUUOrfuKKrekzLF5CF4M/0+VgrVt1ObhOhBHDGf
m9lpl+6Spsf4p6XEBZBAH+6Gp3a/bEd7klj1J6O52c7pMA3nwPijhx2lO4OtuDbxCvlLP3X5MUVg
lLOZQliMh+YtXjqr/sqvPA7XTCLFKgVUNQ8cBMmztuSH6pbd5pnZpFpJwFnzZVdAEykl2A5rRBcn
6qgre1j2opckMhz/yN5EqErw6c+JaDH49hmh3+UZcp43i6QEks2g0i0o20oASotXfC5rA22TAdYr
CrdRaH1Wp1MzMsga8nnRMxAEejnsubvNzc/fzJ2JgBrG7D/K8FH58VDQXbUDiVr91WjhTjLdNVB2
z6ghk4IoA4fauZPZljXG2BAn8tqtCGzBzLEmRPYIYJEb1ZEah6lbKpHIP2VyRVClNzk25COX+glY
Ni5qv54kgD1u8QfPWIt4zZVFyppBM+WasnW1UitXnWi/B7gIROADs3INthYkvVIfp1PIL57HGsJQ
aNPKTC15rFGohZXOPSeZarnBmTQV1j07lddVF30AmLUAWHBV6TD8g9MbPNFBrbKT3Fw26FTrDpVv
PJWVKnp5FCIm4bqOXyuu6/lDYPegM4sXtSnQ1vhPo1uMdqJGuBNNvdebcw4nwjRnSgdLWKLMH7wv
VzFyzWnoA/Vn5jGOkZaEYO9B07NH4UXGSRr/H4jg/9hMGwUxZaGivvMwDBDD4dBPhsw6GYMYKefH
1BDzh4/8v+Y/KvRnrlRk1kpPjG67FqiaJHVdCvD4P4iDoLvjCsngWpRCUZ5RNh4cGeH5W0+DhXXa
ZMq8H5uy9pxWuQ16kwSwGJaDo9VYXCq3qNLvnuwLkevX8u8eLFMlAfSW+e5AKwpn/YZwaudVVPVp
DRtdLZffjzkQGqZvZRn9G6lbgx5kvAYRIVE6jtXwkmrTxNiXwsZLOk4ihj973a9swwmMyKFTyHol
w3oyWkQxoyALfjuRQN4QWQCalm+LDBXTqWZbXN4GJRFnFYkn8R/iKdOWBdt6NofOqlwOJZwLCy1A
okbuTbxzMJ9ih02IZLasnuzEF5d3Eja+/PbrWHLsgyY217EeseFOspJauVJE4qWPlFOH2m/8LKex
JeDntGqQPgMNT0nEYBuLVXJK64p2ZH4SzGfwG5JjHi4xCKx/xP+xtRdnps35bQkbkYTCOKiFyh3t
/7tRhclwLLoc04fW+2zEOauanv1d6pTCImksaecoBDfdtqGX1Ggl+KjJfxVGMYXfw4E795Xon/W/
Sno9bAwc9n50PuA7ZXgAYNH0fZS+jG84bpbT9H5qYuRp8Gr/hYKNO4cJ2ijg0y8TSGoJlAF+LA9Z
v8ejtiMRAmrz+C5Yg++5Jha1ewlDh6X+IhRBem6X1kVSySmLbtqvZR1RQY6sZpnaop7OP9INca/V
XNz5LMHWpzTuzB56RIuVAhEfgqMwZj2pvkBiWAKqNfFf5J8aaVWt3X3x6vq5pX0lX03sW5UoN6/5
cKhLK/c6K+w2t0YL5heRcL68MNi9eYWR4nVvK0INHaA/C5AlJyc3JPxUieY8zmhwt/gdlIGb6Fof
Tp/r79CSvlovLwEeBiegCuxdIdTfeDGbK4/M0oW/Yruvrj4ZMtBlxFc9Lg4d9ueCDMzyOdvttZWp
T1aCM9o05F8z8hFJDcuslTPB9bWheJ4QbnfTaxGmievJgy5BoPWzb8C2gKj1zxbasVHb5KGzydnG
2A0ep/tiwpdHXJfkWG5qAXePREYsuh4NwXujW7t7ROkBt09v8ifsfRpyUdf48x+PFwe7732waZvx
dtCkoPMpkJvUzN49kc5bTOQd/79nJh8+Yucn243OPDBM0SOkjTE8GhvFkbG2R0mGxtguzh/ioMdJ
oe13pBwO18F69sCQVpPs3SmUnpmaA+hE0+nSfllPo9Qm0Dan8vdaDqkBuyOxq2R5sKv2BrrXj7HC
bk3J2BTMtLe7MoxQTeMdD782HHEAtovPhf2auBtZ7KqTtmLByOL5irmnxXm2jIBGMbm0g8CqMZoi
N//phJniN69CfMe50LA+NazBMUdDXVQ9NJTj2f+r2innnZuKC/rqfKAQk1AUaNr1HAo9wRzFl1f4
xpn6Qd4UGPcQTZru9tR0G0xUOtbhwMlbxqzLXb51YDcfqZOp7zTyXl1WXY9egfNZC8eDH7TkNkWE
wO7mtxEazd/+ujVGR+tnXYoBG//0Z71r4cg1DOVMHSbc1L+/sAU5Cmm41P/s4FZAJ7BzuVriya/w
uxROsje4Fc6eTAWt5+SJcLBrBQfXIpnyWdd2pV46qzpDX0Z6hBVXbuSUZqqzTYDypJ/1M5y4deh4
kvZfxEvONwAJnOfeu3RD621afDK1mboC8kaeW08W9j47CQ/cC74ziNYCsflmPdy80k6zZka7CgY7
kVtyL8Gr3JRwoprAuWneAXrkaqBT2ddibYOOmOK8IDey8FSCi0d5CveAzvNxF9jBxPNORHNmX0mT
leXfLJ1P+nQ6Sg8qLBctrh6C5vVUmINK4/MqHO8eRDU2jlXRgBcQAngWDbTOVW2pi5dRkL78OJDg
lBns08J6pKDqQlX9hFnBYSuCynykvgDRuBRdGyrD+iPFpmdu6/z7PeSsCFN0ojPg36pBm38QqCUY
wqkh2POaQszrgNVbFDWwKklEy7ccSYFikf+X85saIPWFaAzXVv7Taz4UlP8aepgnB5xRM24hNAXU
V9h+BS7iFEjpZUr81DGs+8aQ9242EN0VdIBqM62b8DAiVS+5DUpkNR1EJMgff8+x4H04OXaoNUZS
XgTIKIUf02597UZk8+m3DlI8HD7BiBl9W1/p9INcDMvi2IpSKSpOjZvacqFgc+fvuwebVoGKrWxo
7H67GcJJNwJkYuG7zN25QVGp3ZnQxO5OQ4lXTSz9FCqVmR5IeEyLp5/FXY90/YipyP39VYC9yQZJ
Q1GP/jP+SN2xuovHkLG2RdvUl9aCCDHxj2Kf+rFIAr+qJNabb4OD0hUyKTxsuCJdWCZOoLO1yu37
f77w7wvTTN+tKVc2tEROcr8c6i0fQ7P48xyiK7KmdqyBHRPwysDKksyXAuOYeqvIt8vcTJrmtHZN
0E/GH+e5wI4JvJqaOVGdZ5qb0hHo6aGErCxKo5AZKhnK8zFxv8J+JN0cETj/dhk7OYbQ8PjU8k8O
Aw5b1Ovg3MzD/0L3iq88xs3R6nHK22+nBZT4cx+woPsTBD3EkdyF0mrkNlhfBm6QR+jj1Jaavq7R
yN1ZWabwf6AlFYFxpqTaYO/B3Sx5v1NWS8GWchmQVk3wdKmXAqyzINnduNghySNpVZ5MyejigPmh
UbRAHttmci1Kc5ES5/OoPtMsNdZm+ou/dm/r19dibslGQHMNQ4Ktz0Gu5iXqmHJE0LdRWlGLLrcH
wcaWPpee02ru7ZRQxIpXJMM8YwbO4k44mvEaZkVIgRu30O6pxnQBVA0JUrO+IS9w1qHDTJmeGg2X
wvEk9UrGQ5ZcWneUpKvWW6gnZAmQDhu8TpTxNPYkhA5cHn0X3oVmk8hIMl0wFTdTWXDBa3Ay9nam
TkfT1UgBzOZUqAlUZ4E5qMAYy/GHkNza5nvOHic06AGe6/xylJRIKtY0bAq0eJgLPG547pgFgq9L
3g0TynxNeOOimVfwKkm5DZLdptFz58vMy3zbH2RHZGnp70ZyFtkAHyn4aSOwxZE7MGIomomuFJd3
6ZwpTfeUmhv/8O5f/S/u4tYW6fxuRnWK8JfLbHHtP/Ko4DeGLtV0X7eXnKb+JmcZGNaJGVi1RXB6
yMp7/XWe/VJbJ9YGqpe4sPOYdC9qZvO+puCC61kVOawkFnUKjlS07JypYfbU1HJQbQ44IvGTgP6v
UAQtjCCeNW+uwWAlbGc8njgOhanLyiOjmRicxs64jnrh3+WoZxWcswdtW/CV6p/Q4kWTNx7Ufqj7
+a/Arx7qcFc2r9V1pi+vYQlS6Qq4VD5ucKa5h3BBT0i4yu6p6FV2eiZGRdS7bfglz87zF0sGd7ij
do3DhYm4OZQbOnJxIOrnwBBy4tgk83blYu0CUytZSh6aiAOIJIb70412pjFt9LO20+eh2YHmafEK
eguV/td7UBHplfewXUWjx2mw/7XkzvLOPui6CdxVjocAivM2KnItC1im9ebcwHfkxzHvwwEJ5swU
kPghOyCcpiHymTBVNQZZsmIh2ytQ+KiYbyi5GAx742e86XPjL6H66NUa1Pp6YXNjCEYfXB4nnG+r
ErZ0xJ5VKfxGuo/gVwJoth64+iKcBIvFO7zmEWDcY71W3k2hBGXCxZC6WEm/MNva/WTRdbM2TgY9
iOh5I3L6gSZi/xKU3yM+lWtNnoCkY1rrbIRdAyI0kyZsw0dL+dinTkdnp2LgXO5suJjO2jQ+Tldx
/u1aw8nMD+E233OWibdUjdeGOllltWbruFQwFBQfrO0jrT1Y1552PSi9uwtar0iMHqM7KGMLDj08
NzXMTpMAqqzu9ci7RHcVsw3JtE1bhpqqQbWlljJZ4u7/nTTxJMtYkkbgcmqW6nESH8ZH47sZl0Kb
bVIFB6HR1RH2rJvth8tQ2Tb788R7MPrCm7f+YSVbvWQv+lp5HqypFXbaPVDeZXkKFzx1f7xkh6MR
IGdB8A84W11sGirJXlY7qqsQqAqdc0gYi+/7P5vM4m7LJTHgZGegMup0T4FN5MJHLdQKR9D7a4qE
1PP5eLylTGhiiASgx5t0pLHhgDRVek+Ol6pshyT3bABpD1s3TxYsyv5z8QbQ4TiPOz4c2qWmNWfa
F7K+OdBBe7uswA5B444ZJ5l5g+7rkpg+zeN7tWrZMsCW6vwAJljttotinEqwfUA7bcPBcquYxkue
Z5OCLDgfLJxtPxL/BQo0Y04eVnPBLzgNxl+tDUUtH0jgdabwxN10nfoiyljDDmQORiZxQNSOTA9u
H4S9obKM4HFbW12Nh3Y824heUfsADHonlyuHATnmbV8lV5NCUCpIQsB1dHFb5jdTRGqV6uQT+pYo
pmbx4VVmlxmi6PumWlX9XBLzSm0jeb0EBWbUWQtovumMf39jtMCqiBOmyYHLd2GldpEpEB0c9GFE
BBatKz5RH623w4xHrow8GINOPXjWxNPPmTnaAAV6mvy4F7+Ns4s1WZphi+1m/ag0ubRVj/fch2gp
mqTeNbnnh0CRb208kAMXOTqXDURb0muNyKRQqv6pj5id+VXZM/54cDRp6HRqss00inTiitEczTXD
cYhnwTFvbVhknP3EknnwbzNSDWlFMJbN0MyG1YEJPfNnFin0zfJkJvBkL+ixW7uZPkNGoMD7Jzy9
vHmETF5JO4B/MpSzKiXPNSLK0gQHwFzWPkuTMRE9kHTwLJ6H8VKWZ97TtkxH+Tgg2NMGavYTSUlL
hF5VjTw5W0KyZrFmtRTJENdFZVfyekTxOOfhWB36RlBWtz6VRkI6Dk0Kp3Y+Yh0kc3saCdVRYAiE
woQs+9eaz9V/ig6n65Ay1GueCyK+GSN2D9UZKQQJuUfim3dDHsblgZwzKEltQA71QlEhCuLIazPh
iCATWARCqIs/jpllR5aHg6AOxPvs0IM4Pn/nbLYw0LEKRRouqlFrckpbDct1OMmuVdBnbM1mkJxE
8u/IvF61UDdVkAx+S0S93sKE3dv76Z6vs1bcL9B55/CSLw16VC/0HEphfMRg4qWBc2xNv0w/NbDQ
JpNHJ0TgyI6DX6y5URmURu8P1cpsKbf5x8oFHnGeloov5qwfRmJGb5o/Q54Jc4Sv2QgAhy7pwrmO
wTdJS/GVT6Wivm0mBYYb2htHMSxk2Z7N/nGNlFSA/pimS6Z3UCgbtHi7cS5wM3eMSBKYyTjJljuU
8fUpCnpX8T58/RVqVTygX+HrN9Okhoqmq3Ye7N09YPCdciPA2kq2Yq8xVSynaOpPXg4KvhM8puDv
gkw+JWPA8Lgr986UI8iRHMq5A+Jogm/mOkZFl8s3sW1Cto26jYIbZuq4kL7Slq18EfXDo/VzLemx
e3wlsu3IMFao43ZJaw1jmSPxwN1SNaoWMbeeb12SUvLI+wtmVvvLDf8TQPjqfGHis/ptBVPYOl0b
6r0PAiZtn6NICMO8cuPPPU7jHPFG9VV2Skr5WexK3UzjByFKa0zKNPpJfM9/tUcPoxju3c2qW+qm
+Q7wF7nPf2q8hChSBPnWtKrzTWIEj6N8KO++AL0xwYG1RG6+cCco+UfB/kXN9bnBVBKUb3+zzDUP
ZwmUMzw52lz/AMPb6sqe6rSQWVYPiL9+ReQIlTbig3mmTngjMn5pc2dnYIkuK+2FfiJQz8i+YRIU
Z7ElK3V1oMXrsxsZbKy0iFjT2W+lHAvo+TojYAGkp5qNa/9nzTKjoRDpgByTM0/RfByyYMdYsq7E
EnId9s5YUGSADZ9OK69VX7waGMrkUzQrMdVK6WbcifgQEn6Q9lrghXSUZdVYc1DEBexs6DXrl7tr
T3rh8evuykZ9LwG0BcS4MgOuRzgrnYjfJ8U9QkA6c9EGqsWeb25B18eacbeB3Ty/E5vZLzCpesR9
sEG4oFxSDNfNDVVKCGI/caJqP261BcRMS20g3bwysyhAiCGMWdvw7WmgDKRkaYguY1CQ2BPq3+Zo
Nu0YpGwtDO5zajwlCutJ3IcEhDbBW23YKli5Xsmf2k9b4KK1VNLikbXYoVyAKPVFgrZf2eCWn5mY
X6KQcoJr/kxAofP9CG+nxhUEITHNsTaHDCYAc+OE6B6IKMNrKhrgkVRjBAMF2HLo5Wd+WmyoOdJu
FtJlN6nsfXKdXg2MahilnD4VphVdpIW2915mBERNzXYKJdpLSPifMS3SWaPc1D7k4o+pTGfZnU1Q
CMB8HPdSBXkWsGQMMJh5g0GSeGHwAZbifUJi5l9u6po5er3aRKzhTNtWrRfvlZm4gNM96iZ50vvh
Js0nOlFP9+kiBJyGC8RlHN4jzSRPXDZS7vDPerjyBjFnhqeRGMB3uHFL34tNrYb6LfcpXe2ATGxT
sZb+xRtrs4uZVUmKT7DUgtSFWuCrm7bW5Ssvy9vI1lE9QtSN5MpZtI11wdpk4wwh3sBH6ubVxhVe
M0WX94gLveUACNmK9jAcrgK1wZUF2sTWcFaRdi4FiviNkBQBgbT1oi7Xv0cihWPBijCkJfaCqRsT
2BQcoPq7ZAGk1JujqOh2w3p0+zHeTsey5NDk+gNBTW1DYzoGxMrAhCxmNJItx/rAp9GCpJTxfC6Y
MVpyfCGZYUef1evxEuxisJPqSCmKqxJzfIcD6IMfUEqoK0f/GLqKoUBFnm2sznRc1Ush/t4cmMla
SfKmqZdn5iuX8eb+pNVDbdHSBTu8381uhnx7BG+Zy8dbC16iBtvnvdW2d+fJ0Tmijcg6ep0D6hdK
VLdBcx4/RSmrp2vw62cHG+CymUsKRLL+eigOMPgVxLbQXPq+IFcQay4ZKLGjVGvhe5AoWLbnaqGt
WeBUVTr8j108kEv8T3fbU2UCSkPtso/EhFQP0J8u+p4mEKeBGL2eqRLjxT6+mRg19lS1wLtyZ3/a
RY2VLHcznuWyXjSd3sznQIhx6QgjIcmqbGaf5ZIZtcI1Njxbh9ssIr8IUvoXtOgXJlM5N3j5hQv5
GfQPZ4Mw/4w28BE59TrUe0zyvtpurLVKu7o4ZkhDvw5fkQgevlLZKlK9vO1sRiB5MKb5rERwaSnL
PjEG+9XBcWgDVgCNgBBBP7n2KLGxmklu8ByaD2s+/7pi8kfnAa3HnVMftw0fYSKci7/Tq8MOtrG8
aJqOMCjWgnZtiQN0Asgx1mRmVgKCqhxLEqfat9VMo3WC+q3ONJmZ8z9NxWDSUdHHlqMesNH+p15C
RgxrNeM7beCkvZc6DtQDiB0Pqd3UGTtoH5MRpapzDungxanNES5gyd6PF9O4o9kUnw2v2nTLFRXB
9MT/aoJxtFxbEdUiZgiLWrq1dnpykpYPwGgyFMiozHSqE1AXHOOGpQ78GKy6apK8Hq9I3sosm4VX
uNkD/DMPEmq9wIDEv+8VIO1Xhuf8YPPIJRlo+aUHNX5zlraJ9UTfvsxtr4Fg32+UbzcCJeGkOkOL
qnyzGfsgeu7HqDmxL95a/xzQbGnlj5zGaw9DFXpQsBeh6mimflvgOYLc6lITyocTAO6QJpT/xu8f
H0UUBeIFF6kJ77Jh6ddv3137KcphXwP93+hsH9AusDWiFcPlflnCNNFgzot+j+hHqyjjNyNDcnBp
+Uwt4XLwO4QfiADCSvDSxE9DUHkOazz+IvomrLujoOoJo/SSnhhrdQElghEWsVI+WvaJ62E/XRdk
n4GjdFDEsNBaEB5/gp4bHEjJgmuPI4+rWQyG/rQOp/7Cd/M30OUKF0qgkOJ/D2mhSitRmt4t9wYr
RFPsVl+VTLW5O6tj9+TDt2AHiCI6m9ShHskVNML4Iupqpdqv8Mh3gfZevH3+sgNyzlTcRnlQqaqS
gnQZlpw/PS19rn2odfrxJFSjwND1Xa8jD6D54LyLq24rTYJsZ/y2XxaTfniLKHS4O6Mhtqtki4cB
I1a+3c91eVe4WeQuH/rblIuUahgYDlQeNB7AKpTxD87+vGzOSBLoIv23Vri/ZlQDI9AwOzZyZw35
88TGZHcCl1Uf1iYuQbkOXOp28Q/P/moRidaFK3Bpy/63KXt5j/z9DGbS8KPS6xtl45+MfOyHg5dx
QoYHWl5W3AlkxXVQi/d3kOheYxot91ELeJXxw2hzKecDDhTvLgjMHlpqwRVo+5kI8rR0jYaylt2i
l0hlt42asyuQdu8npunNqt9/9W6QrmCiXS7gkD/O1oNQRCR7/oZHDeTdsZhHYsPdApd+HMPB7aKi
+g12RwWZ8gC61BHwLDFkRXUcgbyGnDgMVum8tuwF5n5M3PKpSMmOo92d9Ame4BHgUdkWmOiu2NIA
zc2WwwU76g9FV1On+NwOU+H9HQfip1os5w8c003qXGPHBDagP6h/5QeVEsGdawGKA29dr8hoPuKa
NEhPX3YRy+cpqq2pUjpuN3BHbiF4/flAwaLc5UHl31hMAmNbtr+hpfqAaQYmKBqoHYFpFI1qUFWF
sY672en+fNaC31B5LZ6A09+gw6ffYt8CeFkWa+n50iBo3JaV8a/63kJOISTFMKLwS+ERZorlUeng
cxeEhrhZNkKhzeQZlp62/JXUid+p2LX82JyM2BgKW4225AcPNU7mgCAMGWVwyac80XEgaCAH8dFx
uHJPVRW2ajg8ItHiBGFy1ZsiQRP6rQnWLmLyeSfrBCdhKOBo8V0JeeOrq0DbEdYlFPUn/31Rm32D
NP1BMdHU4wU4qKf/Jc21oD8M9IlQK06lNkOu9eABeY4tA18HXMIoyjWW7vwrXg+1w9PawxlUpnQ+
/jxnhDPINPUdlbt25NAFmNsgs5AmWWbElAqacdBzamXAgCtzCSFAF6bOzzuBUmwY5cC/9J56UaA/
IjhLOUjndk7tct+5Os7MXC5+wRSkPbImxZcvVLMvsu4FwEuiXBKIPHrjEARsYeGUF9U4TAG5WI9m
+ZKcXTpJ189gfFiF+k+KZIlRM8MlgImYgNNlMJgYBzcJn9T1lHT4KVIX0XGVmInuKbR+V/meNflp
YZd9rPd7NC/85hjqu6wr3F1RKn+iV4gqqx/ySWzKEd0Llqz9O9Uven3QSuDrhIAVnSxY6UquPwWZ
MoQN25JkynOgEx/NpagdpVhAQdxXBZ40bfammdAeT8CCZAtXxae0yHF0M4K18si94I0uioonvD7Y
0nri0/O7bgESoLIU2qEQ+USSCujAROEOdfEe75XBl/7WzaKho85nmQLe0qxDooJCPaTU81rwoa4h
NJ2TNs2vZoW7mrlM1T2kTmH/6w2HM73NSu0T7Ok4aMc1I5WUe2PmpO01JKf3DYnoyU6l1cVY8TMt
C6v0VsN6+0IiMnzX9CIft71iF+sc5DeUQQ//efUEfMG2EwxmffFI9I9IDwqrDwfGv17qDtjCmzvU
t4g6sktULvjHUpMPHWrmMsaxm3MDq8fhQ1fOhTvL4W2v0cxTuxJdmc6/hF1kTV3Jxbt9VkP2Dlbq
ywUdonl/l/OfNJHZ45fmTnP0MdIisITosvfmQ+js4j85Tduidn2lhg3g+pNkixhUfPveUrTnkR6r
eFN6x24hAsJMujSR/n8GNUvz4FomzamT7lHddKLujoeUU4qwbDzWkO40mkBRcWwD1F8Nua6Q3vdL
E9VfS9GL7hCvt2jaYhsGauvYU5NPLhO2ba9DkwXE5zwK9j8o2P+6j02QlR3l90Arb/XbjDrtroaD
A8+fuHo5zgaKTD2XBM0WkwlkHTj9F9NffFEJMuIdwxfkvNBJHZZvlqqFRXlIXGfGbSAw4YC4f+1U
jxjiB6UXbRJO9PuSI3R1XvrxXz06bv8OGUp2RgZalWT0/D/o4rrCwOL0MAibNPYANz06QXPj0fdp
8w/VSXYyoSy1jIpTwsPAAbVNxrb02K+WKMGt15dwHgwCccbS7Z4yp6JmB0EKFsoLD9rXg/58/kne
Aj2gHwAoq+Swf9MQF2YOgo4M5PqW2t6faD8Vv8sN9WFi3WiDG31e7r0PqDJE7IhkWapuAoroIag4
vX4D0L008uBhIwtNLPS/ZERRBYlcdh/mHvYI3vrfaDrW8N66BB/1qSh06e9pX1zqRQ+O/ME6wXA1
ImsyR0dHUxdUjStxmz0EWLvANL2sZA4Eo31dDbkxAqLUbqsuBd9IsktjNtX7LXAveigHg5nCR0B2
crOVDNHmgx8SJE+AdjNIXSjWPSxijIlrdEywb0VqcEjKrkoaTePg/2yVzVKA8nScO7o1mV5gl4yW
v8StqneKfu7/HtO2fqe78uVxoPR2rEPP1x/qQhXbR4mb9sXJzncdtKYJSW/fPpGxUFBjC0hg9LuR
T+/fS0LkR2BwWF4t+beHFiAK/XzEBVh9660R2/OYkLZX7ApEZAcDdjkqpCNnG4FBY6CPLwpLrdG2
pjYGPJtIDpza7pjmfRzoLXdYomqkSiIB6zvhD3G0ti6dzosyaI4cheFjJ1HbJexOzwtK3NWE/KFk
Rw9dWSq/n2V3/N899Ul+2teA/9bjSEaMOPWHuIDMbZn33upbBpfJXLwUmKiTfWE9Ovf8hqOw/wXV
VhMBlT0ypH2lj2OOI10k2q/x1esrV/CnHIobeigyZW+1aI4IOUnKWWkamlW3JJbbYMzgwM/PaZj+
bHbMfA7DcNTawy2ikUI+i7JXnY7WBK+LV7S0VO4xudlR+ODoMylUm9J7ZnU0DR3/LcsEvLUCopmO
+gPuFpyQm0c65b7lUkHORmtacSbve4bPb7+QBhPYfn9OMCt7lG+OWRGZvJ5wQbc1+gMRwQZx2rvW
YmoAnM4MeKSQTc85g6FGAfHRcP0zg3hNYpF/LR1oTAAndePCrb3J5NAWBnHEr3Ekh2AnmJ0Z1tzX
gaXVbByAnRVHdSz7TTRV2hpoc9gu1Q5pKUERv70CZUULzV55FJL7Bf0ow9dFTX1R94eBeoH6p93b
TUKVJ06YsEgc17uSOQnigfUDKiYBVYR0+TE6bi5Zd1WftBCuscsAwpfHELikbraegrYby/BtzHgp
xMIHMN/jFS6gKXWqmUeMvDU33SIOYz4SzGvdBobeoPvs9XggSm2tV/NsbWjDrf7COVx7+KhOPFBR
7Tj3nj5iQZTa+CmGilZYf8OJJNxJ1s9xWNZGgxsQ3S9fDhQFFQ3aztsAYyLvr2Lr7Aioq5RfAH/K
O9t29ra1QveAgaJG/HgwnIrSv3wOHzgRdDFl+Hbk1+vPUBSE134WHMU6G/6zTj6u+Nn7r8DyZaKb
bDV95knPNeMqP/HMkHmXxHFawl8C1HOhkSFG1SaK9QbGm8AxOcWArFfgyRaMD69bruc35U6F4luF
REZLp/cjc7j0HnmvNSnltxaV7Y6KQzLL2xRnAz1/t13zSmhnbdOcqhd+2b+S0hFWwrMPMmI4gkcr
vPwy+Ppf3Uv5HxOX1tZ8kPmUe8k/HOZBt2gp9XsFprkawyuRf3GJgVI4ai7zsjUEBbLS4U+4Xbov
Z2M27jJMf00m79SGZz/Vo6pphyxJoHubfOjKfbKHZClcr9RWz/utg4rEZoJi2h0DNNQ2y+huOy0x
WTKj0Ns0j1D7x5XPU/KKV03GDjnAbGQA7EjkHVCS8adjkeuPhSlWlL/lEGYxaN++tTZOyBYP1Ume
GLN3jXTO4SrMxnBoM8CoxM11pT2M/YL1mdsXJtijofW6hxs4stsk9fc5vqCLbwxgES1yhMM1lg1G
iYKGrLEfN4EAyMz3PIzmNhpVk4a3iyFPu+9nhLoTx/65zpO+8k5Ig3Kha3Uss2PXDXY8UTeH6Tz7
/uqMCJYAjbSddpispTvg3ipcjyabAHSEUR8aPQlLuyMrI8ahgIWi9cJ1i7N4TUklnbHVuvWxsSK7
bqPA312d7zYb+9MfGvFG2hYpkDjOfaonzmIVjS/i41ZLGUiWAluDF5Nf8PDbQ6oeBcI/+gJc9cBc
ZJUZIm7DssMqoqhF8oB8eAt+CTSfZy31MCOx9egNfzoFXkhsqjL8ByKNR2eFt/VsbiRz0a918O1q
Xbl6qpiK8EsbTj4wDBYZNC8epJ+eMVihTo34vtgdJyCx2EC1XCzvmHMT712cibnp/g5+tz33V7CW
qIRxDWbhEOCzCO61t8dZY1Hok7zAIulFFS/2G1CSh+4jNMe5KVQp8uEYqtVWHJ3GRJbhuR6Bz6bx
gHXr9RM+NQCGBYBnpLFYjC32rg3Qmd0COUXTjx6zeTC808QZwyGKVjoFKtsuXpqbSH4WWUuoTIeE
nM5/Mot09PfqquVPXTNfQLLN2VZnWJKSPI+AE8XKqDkdUGFALg6AmpZJn7rqNYZWsQp88B/JYxvO
D+/47OPhXvjHVdKr3rfOG+24BVNsuBPGVKai/NNI/KPZQ+4d2Gv/MtnQKqA4So3cAUzJot9rK4+v
aGbeG/xgHGvQsbnlLIJ1Z0rFx0fad7t7S2D6ziJ6lUl7jPCtO0CILA0Ro5X5h7mvoAjZVohjPgEq
qKNBoveZeeDrkHrniQgWhJCmPUqNxHteKOADlvVmGHjY9TLFu7liSiUqpoAQA5TqZFMV3pJasTW3
tVn/DpkRaStPQjI7aQrY26S8bWFiipXIUslKrNF9zdK+NTKm4fSZTKAEEnt/He1P/bttSP9SqRFS
CXSGFh6PB8PHyrsCE9kiRX7Ym+3Y/APKvhEJ8M9X4HqFbhrt3vA2OG96b3XTir8ZmPRTNf0GGArA
yZA2pRVMQgReHdLhPHbkeIX25dtnn7N+HDbA59IqpW+Xkq0QGBq7awuZAHSvCeD2O9t3JN6wbjQk
4ivUx/dvWre8MS04ZmcNdqAnabtxyhr7i8vlo7n0ve1cJmbZIA8qQ4+S2sUPPBRg4HlS2BvFKU7M
LjOYhQjNWfhHxEP6wMvQmmwYXioPBCYk6Ys2RDsIgxB9h5ftntl6hLiwjyOfN0TWqtQ45oxfSz5U
f5KDUPj8d7O6E7jTRL15VmrineS5vSV2SoPB10mOJnlFuk35MJ0ndg1zI2EpzWibUIARqRnCnYYC
Cq093V+LLae/86Ma5p1b03qr8xjQWhpVeFeoxVAqPFYIQx21WjHk12SSSuMOzIOvVBb9W1xYqXGc
mtPUuXStkh1cAkCCff3LwnsItfGA9hyuu9Cdu6KAfFkuabpWmFf3XXDquE/GYTVm/eFK+sPT06LO
Wfnh3jdng40UJI26og/sLlojxLqsDiOrzFZh4SHML+4mczp/v8Xg8gbA17pYOpM7EnI1F0C6fh69
rIBLn3k2eb0q4J2tk1U2nc0zxKD63dD9i/Mq2kdL3H+nj9lZFU0wKwtkAASmbtGgTvRJrcBOldPM
dmrs/g1/Yac+0sDyyR7LB6pYU/U5G2IaWdhLb7qalh5yjQ+ygsH2KoMLrSZyX9zvf4AHlAmvISBq
TGOtrubKAUzCat3joMofBtIleyzwv8amRze2Hqf1TMvk96XXUyt7Y8M9m+51VXk3mdxDD1TaHEHV
7kdgCMMoU+9HPL/PWRjgFPsNMLynJoGJKmnv+sA4fvc9sRk/AoTiKbMvP3Xu3/YJXj9PnUWCo3Gr
FQwUkDhQrHKYLWI9h4//b0A2jyx18p4fXVMYcoW128RQ8SZmATK0XpC9iSxssS7qzF6z4tn+qQNm
epmfi81w7nKiMDVG+vmDb2MJubYO0KiRZ7utLsxXE4ve8gyXL/ybJig6akDn8R5IgDFX8eO/bxQz
a3GixnxMuGpNbs+wYH/DiearCG9NiLKuhrSXAwtuCLKRDnIZYCt1waC60B8xu8uEtIgzEfWsxCw2
lMSQpZS7ktSndF23XWTyOLjxGggLYbFWWyHKSVKKbC0evT/ij+n6/1kZCi9cfhvP6oFgSg7ugevD
RweBhtHwwvbQ6SBduHDIAAr49iJTHZzqiPSRsl060904nNopFcT6T078QzFkrreaiep94zuCkKdr
Vim9mi4PgEkVpgLR+bp9UBzB4wkGKq31tE9nokh4QHReDMU7VcrTL/5tkYDgRXQrqAqovBYVj8CV
nXvdRs1jJTDhqMXWR0Ws8LHK83JZV4yDmDY/Y5DK22zrvllt6r657MDqFpIlc8yhyG5Q06AF5rKt
mF/shEm1ZK0QHDs4cjTHSvHQRexnzlkXtRH5302qmOEITAvT+EUGnuF+taEf04Vj61Ngzfy9moJW
cfx8ysFMZSLKICQdUJGWNwT8l4uqy+gR6aHbix5WNH4q6N+Gvry6ZycOifs1p+45HTLh5xySJRFI
ZMDHkECTnLlzHz6Q97oPaTh6kORuYiElUnvPAYVEMk+kHf+IQXXIEJQmQluHraxYpyumYWjusMCW
+aiIAD/6per/+iPpClB9VcaRD9izPvKWq3GsTj1v2CwO5bdArzjGbv3pfQ7m3NBlsUpc8Ju7dd+p
p1vgSD0t0W079UeEaN3vbNRGF9FC7ZhNrf+M5rTHylUiVwu9hmPD6bdolYpzuiW3v+kLo83lwzUs
a9Vbkn9R11U6R/K9dHonRd34EMwurc6tHzWJxFyYp9F7CvOLl7hljdDaD/5jQRGSNZjlhUIabH2F
5uIFCDRmXWl3szRVdlp03qmQ9sfzV8pJCvGbOHSi7giiWz75CFj08XfPMFBv/3jewp61+6gnl91y
l9oHICLGGEEY6Aa9F7wDPDjphlJXee5NnLkHJ6WunTYRLeWDAVSRfV9Vba7kvjNinQXQAMNm68vv
m35+IBzTJ8DVtmECcjWGPa84bgRDM51792D2Ogt5ByC8cwzx2gtyRGLteBGkp9YAYXRPfXHg9N8R
3Bc2iAW4ixjkcV50bvO2pS/yK5//cYHxNScwR9R51h6rFBJdVlZBZZyyWzPL6j0LxCc+6EXHdfb0
bdafqS2xUF5FyeLbG5yax5sRGpFHix4EeOkuawJF2TcPhLcs5LVmSoCAalnGKGC10o8D5/bQSara
IoStlYhlRmvKc6ema7tYRxQfAzP7/fSJ5gogwo0ESgFaykmr6Iq/QPV1sWdEpWDMTUO/xHcwgA7L
zlDsOF5zvofz5BSYJBeeBzNjRh3peEXD6LbNW11vs19PCI5izYcnZ4nV+DBKEJm63BQrZHvBcqcp
UqcHKnd7T9NJGEGTk2gzfpdcFa9bxsZQQr8E67Twe7AcvSZe4eXpbco85n7W7WVVZs0T1qnbKmKF
V7P78PIYx54k8PSn0jfr93pOx53BSWLhp1cbgrKr4DtoxEwkx7+pk/Ytn1Bk75povO4RU/pK1JzN
T6sBi/XI01RmGMDMMyWlPZRWLRcwcaEQ+VU9GTAdTHUfImmX8EoEsTH9qa/Nhxcdpqwm4LNyNdj3
2wEmAXJb/j8gJumYcRa7/IKJgl96SbTSqUzrJUJuXk0+16SRsqduynLCWBqpk4rX4F3wj2yJ+4vl
TwZqJ7+WxoaWy1YuOOQloN+fpp0ZvpZHfxDdEZTdbHcP0NyGfOZ/aa9Q+9MdHjN8f71DZUrvgGZC
yiYX127aaQaBP5iklDFNnqs9PE4TTgIOgX10qNCwkuEQ49hgs264EWRsJM4dDz+2w7TP7dmXHT1N
2plbqFvclZTw0sFfcMz+H+alsLBHZGeVmEg3/GALQ3XUBWbxLu08sWW3P2G9ZHa382AKzcLcPqTD
mNmhAyWqK1ChPIfaNhgqjtCZImK+9/5JwPC0TI3uQR7DPHMsRLp+HXsbCdS1P/8bVi8fHsaVt4pI
i1AtEzkMdTfSBURmyuySTbbDH3DvLh509F6GRaK0p91T0rEdysfnMBzMtCl8g/jY+WoJ6u6SZ6DF
vPJbWoMVAkwxumK6VdgcktV3NMFl3Sk2k0N9EK4V70I23Wwv8ayDE+sfnx6DoKuTBSxPbKQ1i/7H
TTmnvNicfmIMYWZ88xQh7a7oH9H9EaFRrXMnfyOSXtzoqDB1R5RD6FYZd/A9wlB1hk4+3Oil7lKE
seX2DN8y+DjsAcWrJ4uEU70PmOPpcY8QXvdyeGoeXqfHX2DK07cKkcnhRrqnD/pvKFIY14SCJ4JY
UjuWBGWMHEEV43KrTcnTGmKGcobaiOwGTVLgzI60ZH+fmbLcOWGaiMpxxW4XRSHHZozO2paGneYN
oAeH8FJc3fK4mLpIHTbeSBD4aM1f1xKN6r/CE8Ynf1ry2OEIC9hzBlnjCpJvqeW4EJRcHkkGeNXS
Q/FLVM3Vo/TBjwTmstaQ8ktkO1Ti35eeZ4CZHm+Sosg3rjq1yUzRQh7OU5O3s0VhQLEYDz69O+Lf
oQm0OUKPu+nYol76/aFvOYOFsot1ZTHj14AMd8mrpa9QjPjwf1w01W+6nU3y/L1ZTUHMU54XfA3n
CuS/Sl92yYIc28pklH5yjVC9J6YpoqSw6hk9/Cr6zj1+TcqYt6aZwo6JKdxpu46taTmZRlsyGQ+j
AbRv2NxVMOI9jy/TOaD27eX1YvFt9IH8M/w2XgcNjJmqJ6LVqD5jgripUOXxPXcDoKMYNioMq41f
IuHuXLsn21Da3wsyniRqeywIlYSZN3C+aiPLqJiHpk98JKN3ixJ6ttBr4IPn1rxN+3A7h4/5KK94
4QXGv/ry/UNN+HoeKBQcJo+c2q+Bg7nON9o39iCkluQ76PjFLCKVElPFwijHAumXJutR3vPobbUY
5iKQtz0E+z0cZqlbyw8ovkaIn+o7ZE7s4TIJgL88SeD2DQn9uoRKpK1+Wh8kOJq6N8U5nJKBazI3
q0VAbLp4v5IHpHcq7tlqTuAUxLxMPzNLTHcrydeXeGN67FDjj1bWzXeKER+hLoxmfI948mbScU/K
gmlKpH2cO12C3LCveaMbIFbwPqyZlRyfMndPoYk//qkpkl8C1s9FmE6FTFhQQd9QBT0fd387PCSu
uvwXE9KYPZUv4bGTHlGPizLMaKvxdAmZQlnpW+kTg9f+FIo01cIEHOrKh+OZhzreeMOureNrycnQ
ObkYyprkezXCXbDN8SL4Hi76Bf1MKrFzkcslT4h7L2RNX0fd6F7TmWGSWAg0Vm6mM3jb9CQC4lZf
/eq6wKHZc3lrA7ohLIKmUDdLmlvOf0oJIaD7fZ8PpD+i1A5RG8rrw35d5RpEEdyWXoSEmJdpmdSH
2ODQdAS43HllnUH75QfZCVeH+dqo66em0NGvtYBb1sRwSeVOxlmizKwCpqXovM3Sk/Bv5/Tg9Rzf
jWumN1hTJd9ZvemtmKcFNzYTRULtquYSe5deahlSnJXwvS9d3A3GzJNklCAXM+xmhXbwDEotSmkP
cVydFV8TBtcRqL9+mRQ5i26CiCjltUYbrMAbZ8TTNj+KBNbQy98ymALJWWnjUMx0wc95nd9/IIlm
tAHLdxLig7I9EAuO69lsPkt6E4xeLfwUMiMvkV/vQWotxnfvntObQCxebHzha6FizdyMEmPlf61l
19jT9TUfHoBGcSyTbA6w6MzUEw7pZGOrTXwdFU6Iun/HGGr1153z2FoG/q0AaWxMBbST9ju8fUW/
MvOWZ5EprxiemN3/EhGUwigz+38tzhgSLdzVVFGcKd5JGhFjBEGmEvjNRTUZqhlWDfkrJ8vNZMeR
2EGfU109M5d1KzD1bM9YVvGLOqN1HPXzHpvBnnCMozuy0zq0BI7kjWGNTkwVdogdfAkVq0diphqs
GUTOrzhrXemK39yoGn6jU8z3yqDelBhrp8ss2G1FenVoTIz5GwZ0ZIdf611HlCfkdbzc57f9w4x1
VU4/KOqjpL4/OJMMDyVUrN0Eb/t8n0JjG+3UU34xkmFXYXusa5StnV7uUJK6tCO73BQK2tVL7G9g
HpLHjUNNEX1uFHo9Lc9storOK2vJST1s+gQnOOnTo2vSrZhfCs9VmLCT6MY3glf9T3a4q7vgdOYS
uMkUZTSLIguzRLzLFHGyrtTrhJwngHoPCn9eyQkYxH+yITVV72f4EoF3lB55yMe/bIMCZK423SKg
GHAdHsvrxJGhXuGi9uxWCpNO0Qgejl8oSVBnEQVYIZ10j1dYg19K141KhIQEH0mLK74Nb6oBqYke
88DWLkmM+GPwRV7PL0avT9GvGoUtmuj9VH3WsIupzifEhCmZBVsiz/mal6VM7pGpyOKipytvAXdI
3RyEFuP6jGsYF6n3X4eCSG1zMtDrIM3fF0rCn2bSd5a9uewQaTb/9i2pAk69h5h3iJ2XP1m2PCwk
XKljjV7pMJTsDb35hi1GQlt1PITa4ofXjr533TRDpgBGysqECEgOalOgGuNHEiQLAAkJNJ0yZ1kB
Ry+AECOuaGjBnOUayDTfQtvasQQNMDXTXc7Wz7D4WPN5ixNndkrs05CbaP+JHDuzV+5aTcWqUKH9
mJTOorVL79J+4QKOHMqJvgmAA0626+aGS6J3WGxP3J8Qi3R0G4jnjboRGl5ltW7zFToP4dKkS9Kv
t7HRikFgZkja76vKL+1+XidRf3ooCI0E6FsBiPhgVDJ5yp95/SfKLlmAJ8aN7aZXMsuhv58h7IxY
RyRu7b+gZScyWOGb0pW6OECX+7/8FZ2bTMjUzgFHvngHPExmiShAEUyB914Nc58hQFbNCGvjaTfe
8lp6IKo5Y1T6OfQ6uIVcfCMfdF0Kim+6C1aPjZZlfZmPmKGs/fp2R5JdEUqAznP6htMft8H8OupU
RzCP/auF/DLGBCknliWFx+7itNon4IrrxOXaDhbQcJeQPAsBbn6q+LrDzZVioRAoTzY/4uoIydL2
VzYIBow/fErOltpaXZu/TdKzDb0iKmOHkPUE88nYtUcSkbxfl68wrqDbvUMniZxp2fu0QpQj65DM
EFNy4mMFYaE0TJYSuBmFRfKzJQXkywefPnvrUmaj8KlSUVXOoT1t9UjOXNWd00PbFRI3p3xiM4po
gpLn9QW+6Ekc7MhfyU4VZ2RMqKmWhRU/VyF7INcf8vcFcs68sQj/T6hnpX/NgSW20FZhGZ1LUjhH
FGyC0AugIQ0idVQKzBhRH9sjcnx7gDKgK2dLlSyNYbXAO/rqRIIw2zf5h4+l0J9UCG1W+Pn803Me
ar3Prxt5AnJZ0fZ6K89h2Bk5V6DujwKwaCT3mGAzR2xwdQ0IM4Y5pAWh2tngkDmrsjUi8mOsk94o
yYhdfLiBXljVGrV0xm4KvxYCTAZIioFWuFL+UXZgb0hFODc+8iRP+eye8RzWxDt7+IQV5ksUUjFE
NvoeWf+wg24qgd66cZKXOCR6Fu0Pg54+7p00kEmwqeJxs89meuDY+fes3D9hL1TY7uW37I23j5n2
udKUIcrtTxAmKi0HkS5PbSrcsgtFnMqfzufR/BcPECOBz7ypO7awt8qEwn52syi+tqa+7zxhHjBq
aw4i42vaHyzXbFeQFjHAZQJHT06EucYilLsL7BUGo+Vfu5RF65HhyR1CvIlrTaZnPamF/TIFgVpP
wCYvKm4Kw1glz6XDyrt5295s4WV9NtgX7mhni2GvALZYigGRb7Flr5AYzWZDFqJ00sf4NBUv6C66
DnGb+zDs4fV0F/PNsu3108ROL4yMhOJ1zw6qFeVzA//H9HqYVezgCaUDfDDgq+xpRQKS41+P78+j
bHoHpI29/jHeFrAHeEgmWTHjWUYMhSM30Lsffls5pSlHG8tfPqNdyS2eZlC1ho3xO4jjBykPXYr8
6PHx6uW27HkI5OWqyttzeAt0wlSRkrYGJ3Iz4myaR8D4kPFoN1BUbPmwxOehdqIJxnORb57MTL+w
jKi6H9LQ1B0c/LDiyXsCx6o61l2cxXA6FD7WhD18kPkWQqhjpVTRSZFpw3vuhOkH1Ut2z9q7Ewlx
pF/LTKtjXkm8sHYMZ8u+/btrkz6dqWspltsGAzxppBcOyfxa6kCmmnDPHWUzbC0JN8EMRIwqDo0/
SZYNe7tvk5SJgUXhrL2+u7lgTpQm1gSg+hFA1TBNfOPXvQDTlgPWB9bgWJW/CXvTPglV76OnZ1i2
bnKDZYZnJLMDU+ggTLur2lna+x2uz7EOiUjLivPf8OVCMov7od2pSWQhJlMZXIoMhZfK/tqt1h9w
DgH+zvESXJ1yqrsRuPjknqvP7vFgUdPv0Q3pPDtLPcgjsNEOC1xFcQhDUxVAuC+prazIvDnfp5bB
R9o3fZSYBP10wuO5y5DOA1uIqbBFv8uvLuFSbbfBID8o9syyJFXiWeJEz2T/O6Fkq4WdIWvSY9tK
+V593c857wN3XJfUX+u7lwpZgaRAKf/UKRj+DY8gio8WZx4KYH3+cMc1St8oZUeTvKj/sbkZWFM9
1Bl1FrPZ20gXNRUwveVqj/IFbfZjSV+7SZxm0fGrOm4TH2VUx08J+tBh8EIo9RIUbMlJc5+p+OGS
ROx45bXDXgpKsJZCMK40OlBOwXX7Rt4Z3JQfNGXNTh2sjz/GqgVFaPrBGwGyFcslXYMt0LIaQ1oH
VO5whAYXhvFJzkjMC7bWSiFdvAr38YaJi3sV3HZGNSw+jWgMLXfUjcpSurIliqs9Kqy3BC4kkIdY
hRaZyV8tFDtVqN7MbqV6icH1HOOTy1c9kQT5QjG4vKYtoMc9npQ+gaZXuSGvfFnPBLu0HLQ9/iLD
aOi0Uqmmf45SvQXF8nqsRUxSC2364ekoulsGvJRCxoTVLjBLGOnrE7b8BSXv1aJkWrjbc8YrWlsJ
TETVRiaEAnP8P5S1w4dneiM03dOJeojhl2u3jz5eRM9RQzz6bxY7gQnUnaayvbVlVKGQxBitTZIi
/gL06mjaqDndMpY7/oh2R+OHH6cL3lepl1vyx7nfykpV4P+1eHc6qr/fwEw3sBH/PuXDV6v0AKkP
Sk17XWP+ORje8FGhjdn/jUJnCY2attPQYRFUrJm+ln9gIYe3tAWsRdH21ORPeQwO0EyEp9txPWDh
KVD7kEFIYWaA1FF9V0S7cOGyacqhIPPp20RW+smpgIrhXZyQrTfi5EbTJ+xOkxklLxvl05mKsL+t
6g61//WC1Vg84VNcdkEsot3V7QSjFCwmv/fumq5ZOafvwRrxy47MQQiP04zT46mG0U99pEDnHw7u
oFUM08IlSSs/pyeiNCFEpbsm5nw0xlZ23klwaK1lHDYg2fcIsHWKUXZKh4R+PvVCJ4nzKaDVr9yi
kOu2I2MYr1w8BI3UuJnjg9Uc12pe7zcglpegVJFL/m75oF+sUE6eOmSBMQYdnUkRq9aIQwaKtlOf
/kwQ2s884wXFvdi20DpB7vWcRasiEgua7pYTE6SRchuhTOlcO5N6wYh0btes/kjQ/g+t41zoPKzA
JCAEdvMt1Plm1As864BFCSxyULYnhkBgqWL8l/urKi7zNgeT1pkS6czFTlJLRrPRU1LI0DFJFuZJ
5o6aXP1BiZ0uNBt24oiwzfy/E0Oh835VaqiBhBVZFNON41deNpoxMv9VjYajaWYbmuEY9jOoe9is
X1/yk04g/gnAB8i8fwG5k/NYOdCJesn2amNK53VTY9XQDP8ty0Ip5wQ6XK3SNCTpU7EU8h0zfjF4
bH1QaqDG78Ms7ag5icbWr+nSlLm27zLGuSCpzfeWwbA2taLmlP5HROZrarMtglvsephZRu+bIZml
HSwXzIvURsYvz1Y41tCfhFlm0ypr/c99ltK1k5Eq37ypJUBwgt5wcAfooA+odCj7k051ubWIkwOn
DSBEYp/4vp/NyNA7UNqi519b5zhNYyNuVMhNm78w+3Sw22ZXyGL82nO7exyGAyJ50TpVxLB/O2Yl
8KE9IUeuWDT4cvkIQzSbNNQmCFHdcURmgWu+uelIreB129W0hzk7KXWZ/4jQVQreOg36w2z/lywK
xwlT9slMRc7kwQccPAs7bNCwjKwd+YRJotYZOxFKyWE+/55rb60jkadJm1Hiw4IkFz97jUPF/Z3j
2esR7Z7Si56y/sBh3T/Y8ELlko+VdTw9HgteavT86GtyLMojIoH6ODPoOg4syH8ZuCiuDfTj0wh4
lsASKA9VMLHS7/dlcHvF5VZVOMSqQy1MSiyHb++gwOtQYVIktxFNJGustZldpAUdtirRZLKqBHXa
2TtDPNK/KEiAcPyEZcUB9hyBW4uYPSfpNcTlLIJ3BUnkvG65xYIrrJ9FkDV2iq+k46oUvq1zoalt
DqqXDH8asSqxuDR2+yjufTb0MOTuhdR04o0hJLzGuoP1jbWn/k9AzG2HORW3SQOOarEuMD3Z4vKj
B2QGO6dxBYanjcDdc7gPivF3xAIakk90LWgRgEtLDQtOpFwlYQ1jL26jTZGsF5NzKFx3toZ4y2pP
E79L+TB4DgxMXBeavAfp8abO2IAUQCxEoZCEex1FDA/WmH02rUBd/bMg6L7KhlO0UqWMEaHyHXpW
PRHKfr41fwwlWOgjoys47mj/bdsO1gOjOtcEyzPwHi0GIvWnjKRjGWLzovUPmZDFEX+p+IXb0EKk
r8KMnUOnMhITKh0bgXqkDx5JaWgmOYReSCl3gEi+rzHbSie3l2wqpwTcKVTwXKDRxdOYLPJBqB1q
StcWV+N1HyKehJHKX8tQKh5BeJABK9NLwwlie1QGPe/aLKmJEbKwerEF1vOI6DmgwzUorjRDahA6
SZRrIhroJqmHxgzA1vnMVc+HIyFINeqzDyK6WJi7TjMVrA6aUvNq/0i2IMbVeDQr3QfNWPPJsIY9
6W2YenTNhqjdSob40kSOWgZ8AOymUZ3VKiDpWyKH6ugJAX4E/6LQlRtHHl7e+b3x3hg+JZCoRMfP
XBW0o7QFToxx+2T6ZWhRPTV5ub8htC3B6eNJAAmfZKZBYTUQ+g/h1OI2rejDEuJDqdrgJ6b2VS6B
8PL3+ONpJqna1GmwiReRS4daKgrg+AKpfaMuy+xMkKThwibg2cz8NQE4/jNBeKS2USvrGUWmesEi
d9IMy8nynIA8sUO58/Sekp6x7if3WMY7POFn7wYxkw56hOLvtRSIHCTNTAUbISglWXrrXJMm9xJ2
lxBkjXpy9+mduky4KQevbBNcc1wMJU/+9hMzlTZiIZUGS42dzBGxuGklbSJgzw3XwcJPQkERvP9e
Bu/B2YWFmYOxGJvK4p5z+SWE+u3+qP7KMc0A3bWphgdydhTOgkTJ1TL5lexcth0Z2QbElvdvk195
Yyx9oADozFJZI3MoCFxMACVsqXdRDYwdYLrD09YnJVJalmwhebHtE4AfXThcXtDWM4kl+2bHCbHZ
yenYMeZI82gJij+1N9c0kJEpVs3x59QsoVKLVZKE+Pn7n2Xhw7+U9wkE1W1Wc5udpSeM/ek9iZVW
/uS7hKY/a4K9MNw22h+ij/5sHlq8mQQqlPRw9E4MlWe24X/PtbkITzW809thR0tI7/Vg75JQDETp
V7WErRouKokV9BRrZIHIN4hbvL5yiWI4XTpwpiHSxSZHpNSKRtiPzgUdvL5/9jH8Y043YLw7o5n5
HBi9yOeMQc4W+ooZFa7O/tXbmox7aFBFrM6y+K2u7R7CTw+YDf3wORjjIpUfUjmdBW6TzxPrVakH
V+UQl0axSnoifs1PSTEAve8VYl0ZAZcwsZVLn4UFhSf3xy1qOBzVNDeqnJG6+lWvEEk5yJG0aUFi
pOB5/YARtb6BmT+AAFnCxQb7T95qOTSLjN6gexLQscXNAEWplvVKgVhbi6wVdjR+JfPbBxF8Ity3
quUNW2aj1RENqvirudvQ4SqK5e+fdNHS1vda+9yzzogNd8fzKc6MxNPU20yWaBv0x5odJB7ugGpK
Zg/7Rfiy9fwUU1AWlIdNQonBiOfIFkylUcCE30KdDjjrnWmP/m/wH7wh0iaZTk8fwIDv6/urXoUC
3sAXpfXpfkj4+K2la1UUWE5UDdMImEqZa23wPkahxyyGs0mFrHkOhGXmvEyKc8bAhovOMaDYiHVm
Sc6chrS6PKs9nMxz3OVithDH/3TshSNiJ99+Q4SlJ/n7nOGpig7bJ7N1B6M+NwRR/6xyRt8HFaEj
ts2c7KPh5cP5tvf7dl3s7im1wMqahUkAv9rUxMZSkNJok9SGVswiMuwUMaZROx7IhmzOL+xgAIfO
tMKDIs/EhCXeClwXtt+pyqubg2TBwhLH9KEZ+Sq2I9qaWqRaNY96rX1OGrsmaDGTRQyZg4FMSM6Y
TNbcAYGrp7+tRgm65HeaJxBUz0H34ItD7qW7EXnmesOQcXSN15c/94gkG9du9cFzNPo79NHWb+CG
h5aUYWySwk4oXeSNIIe+Dchey7JAmIzjUkLITqQLAVDqRds24CJkQ1HK0QymS2mPSAB6GqgnbkEG
6zOHFQ1FTFRi/ZwHxiG8k4CvxVqsQISew8qrR1ZXf13aavCKtyBVyXileHNJiiU3+iwxdsIB4Hip
hQI7QZ4v4cIO07d2oTz4H/S6gCRNfTu5Za6rsUps0BoXih9vc0PSCbn6X/us02/TmtAFeYpBvm1P
WhAKPsEc0A23YkYEidug9fT5dyVgdUfFwYnXWk7SZSDAYVHwtpmvZpLkHbRD7uZeixcscp+W+GtA
MOYFFopHatEaRj0wCtrC5lfusVuvq1X/d6AJ0xG9pA1CHKE9Y1Ksbhe+v4HjX1mApIvIhZSdipZ6
QIWojXs6N3uWs64Hc+eUM2VB8saJNJfnsIorGF+yhvCQCmQcTxPworgcVpUzKw8m1UEfpP8Dt9lW
YECCqkwtZyK4cEDzDVyTdIGV/lasGkgp7N+EF0+dzx10BvEsRQ1G2iCASZT8HgfdyHz8bIkpcbry
jLg/UNTLSG5d14620hG3/kue7K9AgR6hc5SRQuTyzot93pn9uhPLxYHOkQ7XM7HzzH+AiQ1ST9hy
yvXR8fQWbLinqs3M7jTXWwGrABgllrrvBbiAA8/shY7b/pCtrnDO6TXfmFn/QbagfF9kuAzEZ2YR
V/3pz1h4IbCS43OLk8WLweBm341IzEKlEp1yQi2xom1R9HjktBn1tABWfdUyI6MRrjC5a1IziDxv
DqTg/ZFo22ajeQPMEHzAZCuE4EBXZaA4+zFE3k2oRXfpPR+zxfxg1ZnZpN60gWFwn2Zxpo9afjfM
TLiBbn+TEo0nXV/hCwH9ys8YLXUPQlxVIpsf8u5xec++9n7LFfN0GBLNi6CVE1dHzmuVHMq3OMoz
ugHdMdHB7yMsXrKptXC6ejiu8i03+4QfJsbdWwTd3HVkwwfN9lbriU23EHZZAlKhcIFeHUBJTq7O
4K3pyduuFZ7JUhn4SAPI0wW7bRU2iSEZ0fYHNsq7zDGzfREbsqZ8rqr9AFq70JI2Az9g0e/1Pp98
myD+kheojSpm+vKxBwEIF3BLBYSyj4tB7FdEzMixjK0uUmBpicRDyl+jf7PKBhbYE34Q05AkGiGe
bXPeAxm6wWiEk4Lo75lBcf3EO2uwxhg4rpeSf2mlJYroD1vw7poZ6l3qX11H5uxXjH8tG/3KXhaX
GOwfM0zL/PbjkE48IKJHBcvg/IKxXYGFYQv/X71NErgbxOAciX0QS5a1gDNbMeKz2vAzAzgExl/5
GrxyRDIja5h/EtavLcNwHegg8r+jN7zCpse+TMYHZ4TTojuxQ8pji2GQI9m76OQRzXdSsLMpSJNG
ZjzgLK2BlpZK1R+yoz81JKPl7kvWXBZO1cvNO4SLFgDS8M98rfYboUwQnOOdDwG3ZF+K5CL4bhET
tEnsUGrvqIZcVcg8aekmiBCObtumDR8NOwWrb/YQiIyM6t4/8w0/amcuuuvFroAIGmedclpPzoIu
jv2xi03vNcwyig98/syNow/hzzdeC8lrMr0egmkVgr8UrMN2MhXutv7eVRq3W2AYfcZC07sLCm4e
CVWFrXRH0Z0USeiqj3J9uHhO/8xb2taBTcJ8aBAupmOOsJCqKIOA+1N2c4aTk05RQ9H23+ERtuhI
EK26zsJp5mdca6CPf0CUKAL2FON983CZDcW2cswv9tsAvAE6y52PkC+lb1Mj1dPWWOcKpXrpMA5Z
WXBfOxTxUYYnZDjtlYRR9AtvmDsOJOMYyfs4A0c9lP0ObruYTf2eUdB2xPLPaNqWlsGqandt2Iwm
0vNgo2UgAq2wEdu/++NLtYZC8D1/5iTxJ3Qar5n6MrqogSxrOhnfrfr/HZ/GelxIxSfPaCLaySPl
63iHKxa70gNizC64cvT/D2DddJRUFpng9MLZq53DX0wc32PWz8thPTGNtcGjiUFPvGE9UpybIrck
SIoIQ4njI1/T3UgzPy2BmDTpVp6Ynlh6HUParsTZ4eVpNuhtPLRClyqbmb9CAFyHM2tMX0DBQrjh
R3SmXwpDkPa1JvKDbknGK+GEzbVGmI0tCY6oJ5oV0Trl2e/LcRkawOdgJzMVJ2yu0u7+vX5fPoM5
gyDZim84nZZV4zHiH1/e3Pz2PU8E0VFMc/N4y2/wP3QFBZ4UfTBTGLtDmAwGmVjOYMEyTFbwIEeb
Q+WRa+B4S1y3Z9/6ndPDEpH7A1sXtlzie4oSORNgzyjxhtsg3qNN/s6LpsgEOoTcc3EhUzcQyYWN
L3yTGok9cmbBkeRDblOXlngYIdZgPUkUQDgBNKAvPDVsYrlkbbG1n6vE7NUY2XxsiAhLCDcUFc9t
DBGZFXAX5WgtqzLJXs5mXGBJe4EK4whsetVMgHtWkzVxg3aw4ZL0qgZufTi1GmKpjRZ2Esg6Se6z
u0OBWUd6YDm443VSFa/RqHPAFJuDY5BZwXbFrvKiqOtZcvYnm/FJidHbmSTvk5hPMksPq1GUS14x
JLJWZBt8konVMKnc2D+pypxM1uL61ouPAB/nPgHpcnq5+NHXtN/SBlYMDsfKWCyPHiG2YJVuRj73
ZruVQzaTXRERUNOvtNTG9fPli81zQc4HVsHucdzFVo2B0CtBDTLYc5TRVGq67Q4l6u348YleMxbE
jZaYGZKrF8mJClq/zz8pUXrYGp8lHP3fY0IG7Z8JVkQvxOo9+UuJe0jBqEB9j7/Zdk4lb6yy9QFq
NNFH5xBVr4qQFQmvjOmsLsPz0Kc/aTyPbiNY9fnli0kHIPcVtecG8Ug57caEhndEWHTbMY79PbDe
Q9OLPwubVkGcTDmHnlskIIxdMt6ixt5oj/NR+Grk+fAWaTqeJBkfLsrqUir/1ljddoGxlxO/pvlS
wTivWadLzErXMnQTpQ30eDeUNDXykGFyw6AULHf884w4oSJRNix6mmESOQZqq3bAwOu6fi0U1OUr
jqnEEVij8+3K2HMBxoMPvUzKxkMRBuYXW33VFQ3ja6dcDOYLtB+tNs9af4NaPvXiSp28z2HRr8Ku
m+ePzU5ByCQD7KBxwV5Kt1FgrG0LfmNNz0HC8WEO1pVACqGl2mflCvjwypmK1wMoNRBd5JYxWSt5
tMA+3+03mwI0G2JAJSHq5i7pclmvM+8gsXU4K3f/WJzFugqbC/4xPC+svoOq6LQnsC8uKMmb7YvA
vvkMr8FLRbCNQpL9ZZY9u1OhGiMwS0BlYIikaT+dq8HmOxA9wclx6Y2mNeszx+XnLtgI1KlUzinU
PQyosIv6F4/GwKHIdJ+Je5a2ijZDXvmi7tS9fNfMXbx0SyMLhusBz3Y2MI9DlIEgujsCpJcyGH7g
2b579C8uzR7hGZaiqlo94xrneM8/9eIOP7C9r4u6NyxfyQOQyRbU4EipDxySZc6m3v8kVF/2G0b3
5pfDjeJVH0zdsciy3pA43Y0CV3miG3FRaBHoL7OdZUQOe6EwRpaYwyuHC+UVoeqZXiBVYhs98fUA
HOapacmPkqMhl64hQqelribI/dIB/5TV18As/FLBX5m9h9RHYS9/J9ZX7mODCsGBSAqT33Neo3/9
BidydmReh9d68sKjRk4hQ5cTOkHz1VqcSZ4WA5cGr+Me/xS6A7YJ/ur62CEwav1Y2qmCrMy3OktI
d4LJAcXiMEiBLGyXrjSiKc7RfyqfGUTayQdwfnnqB2Q0mn60kUhRhKbxijlPiRhcBCwkc/TOAKKL
cPRe3yrvD0V2UTC/vOhcEuVajKqbMUvb44jA4VIAY5hv+TFqLYxqWHTBlkHQLRsquWNBdLbwrqT+
SK68vKn3957crW6YG4dyL91h/CGnySfoFMXOD55cFRC6jEgJB52wIbsVocKo6ATdBLXhs3QBb6C2
BO+NvHw2AFi//FgI/svK4vERRDsKkC4vXfLPOJh7kI88FXXLp6L2JODhCAuC15uhVc4EXptYBfJG
9LND0WNwCUujdrumbJ9cexPF92Lko8MDzRZR1D8xlyGB06OBdq6QO3yvakIIYCio265CZytA6Z6D
FQbDVmFr0ypkZf5H19eAkyAF+f0+FRODxU8bQt+dP0IxHQii4dgbCbWOjzAWpRKaQz9Lx46H/spS
OMkGWa3Pb3Bj62lxYClwfbetRaQaKWwCQvVfw0S49XtAmfsuqfR1hgaoBsI6XHOBmvREJr1qIMbS
mkKFLMtAnf8/LqbmH28zmwAl9bqKb2AYN0mWSikyldrMxblcb5PyaPrX90Ebs1Mb+FCNu8pWlbzX
b6QaI+srDpUMKy9NmS82mRABhEI4cgcjYANaIWtlbjNTgvFIHWkBgUI6kCUO8zQEkEBNcOPUFN1r
Txrk0otnpWhj9M/H6AXxKhpf77A4WzJt8ywwh9T8Pv3MmjnK8aAg7MZz4lRaeExXIqd2RwckyP/l
fd0d6a7zKb+FwGHrgs4cSgZmyODKuUEkhA4ySUEiPAX88YiAtW4SghQahCMbj58V8+WJz8JjtKsS
+iABQ1/+oZqss22ngsAJKX2oUZ2Ji/45T3vnSq/NEtsEoCOIsb2Sa/LY1sGUCtFVegTW0wFO1pNk
hLU2znZP/gGY71yey5poKPCfYEtDzY3C2PNFngBUkiqm44KgNNLOhxnAZ00TSGbXccM7Jyc4gH/Y
Do3NAaesvYddsRojsqK8wpOdoLs4i5xQ+goqjPWKqOZkwP3SdSye/smWMZY1zUR/1QXkApM3hyqh
xS0GqLu6XNjc6R8E9KkU/hEZYtF5QyW/RXqzQWRdLDNK1UtfwOorDggOQF+i1wLWi+fx/FET7T1p
GxYblXVAvKubd+5XR30BrlSqQgzJ1pMFgXtcqI+hNCNQzm55YrUalMuKQhxGqjMMgi2K+5OMtMrR
+T4dohzqozQCQxAeop1DCjrhKgbeD2e/n/quVUyrhawe+qyx8Za8qmB+zEBKPnrBvGnRdyQ6T10x
fGZN+x48/uzkWZ1XWkfL1ImTY2jiEuYZMnuzLtl/LXmyoZgPx3YJPnAl/R9+SRdIKXKbeq4Nxwpg
OM/y5EU2A2aIhOuWSdM+nfZ/uuMGonaQ65lePJdoRMpWkFakPSEUNppf11jsMDan5mfRvKGIydnX
fc3m3tkZIUnLTFUWUCKo6xVrzcPP2ejHJVl9dhfo5QxSowsT5/sNRZZOXxaX2dtDjxFag+6cJbrG
OkZ+kKXx83fH1bU2Hh9dtz75ZhQaMqIXVPeZ90qsEtpougp645QiH3/pzesgD2y0DgEWUjws6UL3
80PD7pWFulI44+SYI2Mf3qhWvESJROAx43tqDAfOscKJzRMb4v/UavZ6ETeAK60VTAchu8pM0Iku
kbMJn6KaqCgFmyP/D+hjoVeWa/ATCBGwp9zeb0KoezsZ23hkUcehUKpFat6b/3XwVcsTIVpOHM6Z
ZwI7eOYf6c0044LABG5pTQFmRw7VQlcJZaCo6n/QaoRLF8mmWcckv9gAfIsLQSkPmwSyfYgR4Xr6
iI2YhTbzTDxeeQI91w/urBPE1a8zEm2UmSRc/77kVqYFoC2D0qgsPtER6A+y81EjoiirzyCQ9IOL
/Q81OV3z0rkb/Vc4lGbCXJ8FF0fJQVJ8ybzYFgiwo9/YLQpnNx3f/ELvK2uaod5MA1pkGe9aJisb
H87jtKsbUUIqdDQtwGIoJe2PinXtz3YlFqzMJu9ezJKCVZ2CaG35umvuJsI5xB06fFe6pjeCxsER
XlmvlQ/JrkfYcqpuh74Ed5IGFTMCpSENH1HV1eQSnnF0bwUQsti9saTNAQzuamxIxMWP+KyJFkaJ
2Ko132ZyerXzKMvHSFO8sUZlVgTKINSWm+AIWvMEArWDw/OQ6AZh7EpUiBAGhLt18ZHvZPz9b/KB
VeYFXUgPi340v1kFhIx8fkxkm1SfdVNr3AtYVuZAzZgveUvBaGkE+ynT72CXJcaT+GxF+ktN7YfQ
lsMIx5RbZA9pcxZor7oDs1F3uDK5FTyZylApYFKYXPTTWvdP6IxXAE/vJfqd9so9qeKDjtn7K/Fx
cRIDgL93vktrZVQX3/v2lwz8bEy7hJMqvcAQF8LsMB162KJwLWnSBE147unKjbzwZItTA4b7cVTA
Lnl1DvO+wlZr8sT/vZWwS06pn1Shd+ZxVdtQ5m6+cTUfBoMhYyY1AjmT7vxIJd6k5yGHZ19wW4Aw
7TvkIkxlxHJl3vyXZljojJoBleWkfBF615LaUzM3zTbl8FgJj2XcDiSifi7MAb64ef5LHbUrYfFL
nxtHm28BVYEPOo2xRFpciWTaaVmW0z5wNhYIZ7CvcbaWTjUiUe0E8lUQVp00MixEbCNjooZgomrO
QaMw60PmCm5GbImKi5n/Ba7hh66ab9lfMFYUXjoc/X1uPa990pfZvXUgKEPquw9cmvh/Ru5ThjJh
d9bLSbpNJFrvAX6ecBjuhPOf2FFsQIJNlSKahR4aXiaGhoLAPZxYMN1b8SbZCJHT2Hsz58I1WBX8
0LzDqZpVSyN1DAfjoKDE+FKP/30grxzw80O1DIThbffUdjubLXxtipHXkju+4GnAcGZW2lQz/FpD
KRfhxkkfegdipom+ogHr7S+FuWIiCXAHegOUF83tre48fnrJFANVkXCmHEKfmtzSR1uTxxU8w2gf
ml/FWPbbHjoSuIvZ/tkaOYsHbl4oOtZHNt3sP5kY2G2f35axPalFmSmhMIVdeiWcRDSwxcIY4S/q
4Lmu0pmHN5mdDKfalNoeqju/HuDrU65OFcR6BOqWLAhgnaYg6+DpmFTvAZqIVh3D7cs0jALcYPI4
0sGMPszh9/0SeUUG48z4hYqCy/phfc21zAx88KFHRbKbfJCpX3pH/+AjRqLAn0LINsH3Gbc0Bemn
+IfamYCOvNDkuG0bnkCJKmesWP2rVCyK/5ym1KKNNqd/t/ZmY9514PcvYKKnLkNEJ6sV/i9iFbh6
/zA4oGKedoyMQiTIvlsrum9Bk4CinlYDQyEQj2k2OGsugQWMe0wM0rXQSyqbZoqTDA7zlCk8IwC/
Br5iyMShve5ZhoArTauga3w4kIzc7fMj7PocEhbt/0lld5jpLuiT/wygkUjLB1SpM9GVwmTeDCZD
0qYvMW3rryJ3Udga0IeZh3Y6jkrlYJHG6lxFbE/7QUNSVU3xNKsCs9KkFpr+GP27fClEcUmE4kp8
S04mObaNrSA2RsVwZ0TW/gccTWXL4sinqAgOrIX/oTD4UhkqQNnNOxlkAWxurJdH5KvP3fnOLwLs
dkvRksp+vYucjfODyiMkMld5JubbHhR7pLPdkZc0/LeJtvaVUqJRCUCfrlXA6TQkvxct7vVsePif
xRngV54JcGFAiTSO857QKfwEuZuFrQRUheTUO5MgkcTqhHl4KVVOTIw52hwyPV98x6lMtNhOtvvq
Oq7oXnszoaWI+hl0dBHiP8vTW34YvRoDhJ034efzcLYgVEIA4+QmFTwuC4r2m+2/g6tGAlPhoEqV
+ylALykbnRvfM7wGc5LRrDdJ3jDk7QCXspfUsakwXvXdjL32tgsRumUZvOkFguLwam68XCBMLTrg
LWEl4tKLdt5knZ+5o9gBdBRq4Si8mtZpB4ZjJAwG69tBq92Bu0EpGTEpMV1kwRYqqEAmt8G+l5tl
M+MQH/e08T17jvlxI9+AVA87EDtFuWQ7wM7MAhuVugsWuqoDJDbvaku2A8WHfW0pXP9p/EswOAvK
40TI+bK2AFxZOCjinjwxHQ1PguQdFkJwzhAChdR+eKFur3oYPvvgrb5GDVkZ5E+NhXEU4rURDWD0
IqTZ1tLmZtdxI7bQIWErsylFWWIVi6dUY9jN7azRM+Gt71heMm1kAi2Lb2PF2xmivvzAeF0l6psC
LJD2lA/ZgxbikAjRZRjbUc6iwkQ4c8CJXSRuI3vrNrtlycfdGn8MgPnTU4nmxs93sygNronaawJ1
9O7huycsgC2RMJSYj8MWTW0Tg9noOAK7/QxutItttz4e+kXn84A2NMuvOsnRBoaCN6WwsL4pA6s8
eeHQ36OG0UiIFOLDXvPYaCwgBKOtZjDllKvGfMl46CXnKwTAObOmcjnbVFLt9cyf2kABLuIbC1C1
RXzvOrlfAFacPKzKq4A016DIXzOWRlHhiCERs0x3rxBXdLHU+YHL0lPZuMTMT5tByRGarMvW4+mR
zDHMSsdEr3PhFP7bT/IHCqLMTI6PVXwQahHgwAIT6FC7fxkIYZhZ+QwxZZeFiRfFUeR3f6X2SahH
Yk3I4azar3VCvP/nZYO8W1GugM5lCnYGbpVF7j/+aLg3WSjYn9Yddw4COSqDe148ZN91djdUB3oR
wUXOJRKnSoZqRlNh25zuU23Oyh9HVChn3gL5+nCLoaBnkhzjW5WpyQ7XOCh9iMASA/INnpc9Tc4s
Z2ZEE7bteMNVGkz5hOX3jWbLZg8XqG08nbu2mDVf1IPbR5LWxvqc7+DiPzPbeh+pn+URdlivG30V
ifB7ViSThIuQscb8swHBYTKbUjzF0IND+hU7MzLhRTVws1bRDahA9qwTrkYeuBUmnspsbS2lb321
+ASXqOR1fOihC+bNu3g0xkDPUBwBDhC9lxxE2z3te0M/GzLraBCF0HSxUCHfJiYAarOSlF/FJyUa
5mrrKd+JYD36AdrCpmzc839Z25hzRhyxXEcBRrjVJD1mDe+gNGu+VGgC3KIjxxgGpH1tDkEZOJ91
9u7UFWrJX5fLlqyEmC+UVdnhb4N9VckPBBJ/HuRzi8YtGdIbX+7sDK/re5+pxP5V3+GMgEr1F9fO
sI9ir/JBJmM4vIxJsLO7eiuecAxGOjkOhnyNdv390gyBlokjUZ2BCh86AHaguAOqXggg3Ojn94g6
bC4VaUaqgSkGmuAYsmEY9SOr3RzHNbJLTDYrrprgVm4jmxpYdW4/moMhEnBmwHwdklCzUCc9oVyy
A2DsJPvCTVjB99Ug5YH9GgNIqg4IkEXeZU5vQ5UxPmQwR6brH0/Z2posOMNUv9MP30QY8lWK4GnX
xhj8A0wIJkidO/2yskHdD9s8wutEr9DBjevAgxNvV4SzeRkFI7Yw+pg6frJJdHLaYrmpHpgmtl/4
06847fISB6zxaMzOHH2LZhPbbyEeYZ8I63Yg2emDWsQy5817Ajm/mQT2PDHlOUV6SxmEoSfhabab
Tc9j7f/25t3Rz/Zm3fZ4MdpQClOXDvIxLW3uA6sd2bZ+F6OS4RnKiyYWDqMsCm2P41Za8yjYa/eQ
CzPzxit4lA5/BJfO5YAwK21G11lyZ5yITOgv58MND/dRbm7fL5vsjfRIIGtMfuNe0QCMZgCOMho6
RAN1CDSo73JhKOIUk9qqVU+sQJCUOrdZVnyZwF0cL6d/jTFS6NUKYeMws1CJH6O2NKjcIwQCiG5q
r7SPqtpmGStwu8hUfgJ4SEW92K+8az8ASzjRy4ntJAYKjb1F1ovRKbmYPwjWua8XY07FEE4xbH/N
0ogzwj5M7/9Y6I5lGPdUNXHdTKH/Nl6tnN3g82b5SDwBqurywEbjwD54XRdEFrj+0vWR8/3h9S0t
TwH6kIf/yCQpvlsXUEk6Cadc7k7W9od9BJ9mWcXI6XXc8Qg7ky5A7CEIUk2Lfd+zi0VOLcCd586Q
Di3/NinsPMo/CoeyMU5dol9gbhrNq9mwbt4tnBIxoYVbLUA7pxRlT9haqPGG6tNv2elEPjSd7Dq4
oxW6+dCKNMK1RjjVBREcTV5UsuFHs9VGo2ANMiVXIP4TtuydDdHL6nZeP0LIT3AsnTkxEKFyDtEg
qp4WEOCGZMw7NHoH0GAxyGpZyrv0VmLF/4ga4mvRYA0CMthu7aqavRfmFD85OZ40UOExCPodgOXN
y2hinuTs5Lb2B6lQdF8D+w3oqnldqpPKSEqR1Oo2pDtKvYy9MVZXLmZMkC2al5hee1/TmNAgSF0v
IAvZMzUcAPyTtyGrh19bm/D1GRLiKvkcDw1anYSdjR+bZRkuTuwl9QQ1oZm7F72LZ24iiyC9AaVg
7ubbTKEFn5gIELsDlEXDhffD3mkZgSxNcdX58sIF9gEmRDzk5MV7yeBjfQj9QVyhXKLFjP5th49p
RSs6ru2SflHpYN9z/suTvVSgY/zJLVL9stky2/UpZPti2xwRNAbYiAoC12zANbOww7ZMG8W3Px4h
zjNyGw+iZk2wyYLWYteIMAQSHjvcl/o8Ggufbiz23ccZvBngclBHtMutRdxKaWGB2wz4J0ASV3R6
vx0B8vjXGJFKV2QQ646tz73bi1LM5+BWq+EQoahmRgItct8VM3iybXC//CSyaOy+xAecrjO45YgT
WZy3LEycwt/RkJxOno39uiOWbhsJOkYnGKAeulcPrNXh/4GxVEv14FW9zUxO7yOnSajjfAS3Joqi
7RQCa/N+tizkLFEYmAJsowGBBS/XlkcC8IxUwNdpFqBvSncg/QClbMNzj9iwxMgYLjRebTi4vXWS
7hZOdWTKFPvYq+woub/MGPtw5mKo6GC8ELJpTWPt4v7e7YxTv0h5/gqYI80RovZS7R0KcBoqwBKw
V8Jev/JjNnuYY1kyuj1Lkpxloftn2cgyF5nEaDzD9dC4fhSplBejra0Ra97l1A9fDDiyz+iIVXGo
Hd7yDLoUeqk+CLKTPIMtrd5k8drBESaUcpflV3QvTfWYHp/uKEU6FVlu3qsLODkWurwi35OWPTBD
k4BuPxtOf5oA+HQvo1GsDAl4ZHNCDwR8ZgHfJdm0+E+p3wxB4NOdHy10uiyQhtAgsDuS4N4TAOsa
nCZ4jne+XBwM5e/qG3XgIAsWHRVeSppBRE1Gi0c6KNp7Xi6v1IbVcxkc9Zc2PXvW5FcBNP51E6FF
YZGj01E8eIb36P1VdwtEcqsGXzBmkfmgVIhspE+TYa7r6vmpyGdOpa5eMT+Sg7oFza5R5EZ2acNS
Cn2rTm+g+n3KPfuXJtrsUuWOThNb01qd0Z0XoWj0JamZA0ZXGG3PKEWdQTBBN46AoxabMyBN6bNx
LRCLwh+E7XdX25qeO7ioK34Y+ih0/2ThsiPFm/ByU1P4xq4bI4xpJwoAIBobOp/SgJkKI/zereBu
xigssJdys+pN9kAQRPqGFnv0UhU8ozJeb4ZmAgOxUGZW2dWnJG34A8Pah93jvxz0R9EaBbKxRP7e
XJ6CdtCkYiDw7sh1M7AOaTrmefPX62iIB+Dr9W9q4UWmkxfM9PFw+h1E0oA/6g5VPiYa9BjIovk7
84brMxOPqbYLk/PIo/BYBffOcOFCmgR1H8W0CADtJy7gxTxjOfzQqaR73uGMbTGKc11eDqvFnlwz
e5BidklpA3j1/s+9rCr0ToAX0VqwTGXe1uGMSLs7S+F7Qv0wZzmcP+fiv9+SSZHiq5jRyO5q8S8T
nSHybLO8chR80t1e5n5l1XoHFRBElAHncOAxrDQIwAVrHfubU8AKoOrhtaoUqfx+kj7AsuexKqvV
L3k3cuVGoEXFA3E8FId4coyD2nUHXXu2DY1oTl4CrgMJ1TihxWrQomVAjLoSfCz0nYxvVi0YBsXl
9d+jPOHOyyK5nEkSlSo+sXM+drQ6GwjjoW3IYwFNuOEDZ9EPz+ZedT7ncv4kNUj4da9ibCgv8WYv
ZFTx9rvYbbnRU2p2thmTk4xpCnN+Che7PtN6CifBORfWK6CKRV7qUJF/OdHqe3F8eKs+RGDxifBc
MIa/+PItF4aJEuNewW1gFy93+/3FmM+Oko0JV+v0272NJdD3OoaoUq4ylQu+Xz0cL9bF91iSB8y3
PX83crOBy7Ke15B121HMTAp0KlfVBgcL6N6qb1GkdPWL3GlDzt5gscCoFxRecxifiQBUH6TiVyJ/
5N6OfdsaH3qnF7LZh1Pjs7OE/7h1Gh4J8Pbi5PRW6NcO4xAmrUQ/2sWiyzMIRSx0TJOnWTqrF3ZO
C8xAbfOGKqgHpuXvvR1q3FhYt4ZIVLGN64j0Tv6SOh1f4QFKXB7TChPCxEqsREQM5liHSRQ1limg
y3P6qgJcEpsQEHOjlXwspZyWaQ6JC+BVshRHVdlH+GY5fJeFHj4csS9ZnsHjHdiPcOMrQ+Kg4kDv
UveLX0kCQC7faJmJFCeDJODT1aTcl6Sebi6eipWxS+2AAn8QKoblA5h80pYmXtzenfK9CncTckD7
KSyNFkUkWUr5e5AFd+4s/AD3sZwM/m/gJL9+6p3B8HslfWTsu+n/ArSfz4MKLibGbddKmpQEtPj5
7IZjMf28NmWHi5OGbBlGJOWYWj4fZmx/bjnrzgCF8RqkDAK8KihBAmZkHS2Ju+FkgEcTJe6A2Tp2
9G43NvmX9TZEXBZduLjBGEeNKlp31x7oyhGHM8vrY2JScMi6J3bWdTTwSWvqv5J9cTPVu4vRThto
BpItHUtlbuEIuncO7YPfwijVgvs4hPZNnrJDGYpUUimbkQHy25/jaRJvj52UbhqENvhtVMs2McuP
UWQlkoCbDbnq2//QEgWQrIg9H0SyozmnEfBNqi2AFWjZgDx7MUXrA57nyOy7VhXutoSNszty1YYE
iq+TH37YsjkwDQPZjGgJojxOy2qGLrOgfCVsuxN69MX74dXWam1BART/yI8Zr0YkBDS0A2B8rC6Y
bMJkjBljDw28zpXpPaYHBoOQbyxeExfEr8VB1Hh+kjKH+VqIqWca1SzOi5lmnmc4Ac2WKq7YxuO7
TqSGPxkYI5WjPQkiiD01/u6lairInM/19hhllHVaF3uwko/Y/HCCbOzBQRbJpiYig7ZunrkxeX9d
2wK5rmrNpxgJHoqL8rsXwAp18cmDOItqpwETE2n59aOc8LWUhPD5fd9YQxrkn2FVsdN3HRaKdawF
F+yxLFia+xydJ1sOTexgYYyjs0crIQt1ef4vY4Ttj12ygqijq+v+9IiQY5+WNf7xTYQKGNUX7txE
r6JBBmn44p35/VCtMzipCtNJvtuT5AHBsKg+tzwhygRVMNYy01O2LWXaM45/olUP+zs/mFyzIQAh
9VYfIxaKRZTWC7hnsuJLofJK8ZMH3qgq8hlw+w9qcVVneL/HQsfd3gQJmSVUyqRZLNI8G2Lv7JP9
vElcCfxMWN4huVfWmpqFKqAzolbp3LhmLPIvbdVIsIIbwCvbTkvPsoaK2rpcT6zaMvTOXSqW2pun
htFBIg1OS/31t4rt/9Y01KWI1Yj/nU8k4IQAtVq/l2N+1p3PxhGV7TDPsvmcUR+Ym5FXNiZn9lwx
Pg1feHNDM8+vLHRclW6f8Lpzaf2Vm1ALlrLKhB6e/yKw0F7iLCqo6Uz/y06/pZpBPtuVrwmL6kZ4
IdghYjHJSS/SicKEVazcsBH4YcpPnVUZa2+lTDFyW8j/TjBthwTkpbd9NODOALOgMINcyM9m4oUx
58wYs3N65s4N/wg6hPdKHgwe+xwWev/TtC4jIrNvJmvI09XeJmYr5Kg6usvodJvLRlU/XHhXKToD
W060/i8x8IK0O4mh4qzXJUHMtUR/wrU0MQQ5WdhNbCZaKke2kVQj0Lk1UHY8fliC/Oc9XZi/8LXR
pwhNmkQnZ64sbNoDDQ/orA+oBrxHo6IKlCpURrHSmPlaYDB8PcjfhxyvcaiKsuwFSRxVlZO2uIa7
8VUe+UdPqA51DJ4aJ0r8elsfA//Qer/NkfvsVQZS8Mkua6LhSvpQMtp0eLpXMnv4JxVSCyxg+mOY
wTug5/3Zoxd55acmQLtoETl1+srS6v6/u9kHRVey2lrhcQqWnrmDTwkPgPp2OhP9iDJttAaFJAUg
tAGZSc3JwceElT3xAXz8s0ZKztvtZArvQt9TEcmUl47J79vaE+AGvSwTJeAz0Whvq9APWJ9EPwHf
dcH9E0GUyquWyywIiXHObNjusJbN9d1qlQUdvSYJTtzmXGpXHVQkUHIGhH7BFSEz6ySB2+04YRjK
j3rrokwIfiZFD6lk8OQmZf2UxbZtetT94/B476qyR1gx0sQ4pU9YQJr/35ruacq90Qm9/LaYAkV3
gputcwVhd/UnArBLOHkexQ0zzRdLu4IFg1P2tNUKAGOh+05oYLOw3oyyRMIpxSyti544Y6ZHjcG/
g0T1qli9VB7eXkSHReoVOZ5LkGCeEy7GLSkC+q0AmU86fX3XDFpnOTuOxgRTj8DIIvCApgVee5mG
37+qPYVuwCnV416LaN4uQj0zUXwEW80sdPw4Yfr/Exhh9Bm4hXWpVJ0g+EqDZcdUvD0qb0Ok4nAb
reTN+0kE62bOi4jv3l5i6HlrtwKm785I/5+9m9TiAQMAcCljycUCxwTkzojVQqClwZ8/EDH16MkW
rg4ojOgyoJ0Ud0qYe69ugm20J8TLrgTB7/p0a6BUNeS6BrHF39uXRZh+qs2G3MXUFLBzjtKyyBjo
sQESMNHdpi0Ou5BLj4uB2xBdUTo9Iazw94M/i1CcuYGfAi8n7fuVg8iN1dEDd8w+23jiIq1NMYL+
egsr8cNQvz0mEqnfpEXaar7NioK4yL8jANdRZbguTzoEQ+mE8PGTruhxVf1X3QHbw+nRjDzAJjYS
aBFncJPmk1PiUSxHGaaeaSTCtMkjFx4shS0VwtR5binaPwsuCFJJb2aU7Wmg0OMExPLpmLr08EQI
jfnse6xAGWdvzAWkQV3cv8856H7CRa2zw8tWwnJRfpE1hBGiwGihorDcrCjbRlM3baRVSYOicHZQ
bqspbVrlbN9EGJrO13mCG5zfUU4QrAcKKN+BNx/FiH+utIwRlZPfaQX6/KGb9LvDR/wVKU/GMQMR
gnhCeXmpwrlj/UXLYvFpo/hLuz+VouetUJlWqOWnzb6eGsMHJWxiCijO+TGP5qZF+eq0U0lwHeGh
IWQk+YGlw2mOg788OoRF1arS7K+2wlo68fARavVVL3suE1YdGUYPT61u6f1nAk6sth/DY8JHfHsY
6JHADcdrlK+wNHUV+/0WPdOFqJJzv3dgi0kRbGji7W+aKbxN2MjjtLTFwgnza1rSMO5UBArSYmdc
8JbudZkYa6tyxnSMg61R82lNJA5mp24VFHcSHiVkpb9rOhFLwrAujTT4NOYcPM21euYWut/kBqbc
mNqRgxNsXInWYJEzH9UEqJ8Wva5RRD0V33AJWfBAvA4RN0WwiOzsJiXOLGDM4/MD+avozCztXbC4
VvqQYVSUyoK6Wcp6B2Uoybvapn5/y0uMXzKg3+AuV5biLRMsCQXwwYPyD4W3qZUKYC+S2HO3Exr3
7LfRrij6QZNFSIMQuFehFKDde80CnUh+5+ZplS3mFCMUkjnpgQ5saJqptFpxJlH+fJG2CIsqhVHO
kIsZ0KYpuNKwxJXyNHJr9Gu2bOBPBAi+y/YFBXmu0f6iECto050SuLSP1IAVnltrWgOhgbyrbELA
rBUY8O+qDBLfQ0yv2UL9eV1rJEk416vCc/leg31pFIgDv2nCCa2qOIYHCIftIMVfRQFsXhE+HgI4
dP5XNOQeL6k7awoqn3elVWBw2blTWOzavCInM96pP0kfRAa13N9DhOPSmCLEOMG0i46em/o7yocR
ExhpqnT7rMb+kgGhvL/XZbk7P8+jli3HaVF25g3C3t+dzVDW9ABVJKly9Ph1Id7p5vVHDNfLrlhM
AzOVV+w7FFLLHHJKXnSwp5P4dRVgY/aDtVbGA08tHYTJK3WYrlNKmOOnXr8iwm4BsN2wc8o2ECWK
bGbTb7ZLi8tmA47mBaCHb6TQNdKfntxIQBeM2FrQz6NDw3iPcbW4V72/zcR1CvAqXGxKLsWBnprX
sgPDCTcThI/0eDHL9PFGpvpMgg4A4dN/iblld4nmeP9U27Bwq0rJu5lVIvkKge+kjXAhfZlxJ/pk
ET1MNLTgvbBk7R8Jl/J67rzHw9ZSddk0x/uhAd6zsylgrrvhdPxZLMBoUlnmEo4SI2fMCECYt9u8
13Y2NXnAvNlINrhqbVT2VeJ+sqlaFuQfnsbnu3pFThEJjRBqqgmBxFy5HHpltU6MTOUnSkAmdaDn
5zE7k7bMXYVNILiaoxFnQJlln1G9R7UrCRE6oHlXtG/GvRRip6xxYffO1pfuKImy98J+fIF0Qe1P
KAdsPW/i5iG6UMNX4GenmC0mPkwidjbazdf7baeN4+i7Ny8tFhVWkarBS9l3qh1gWXOwAJIxA51i
pbghb0W+9wT/wFREMKWrT0sjHsqPpqynaUg5lnjQNvOYuFXX9Ny9FMY0rgFZDyc/dxFENrNIcDf2
+Pa5SlSE/SXUaUp9WYh/nsOhTtqoRrx05FrpyRg2q46v6Ps4HKM674B13q6fZT6o4mVJy+NERRtB
5WZN+qBIP1s9eqea6jiNRTC4A0bCMEf/PbwP0l99L8XMvz64f23QNexeBLTdiVRzVPkvk+MvwMSd
4yuEn+eu+yAwrsS/dmiNVVVhInHrgdB3yadB1sW1DxDVU1CnbUG9MxDpC6DLJtT2SMRpYPIG7TuS
9Z0UYcGy3xZTN+9lihWuQiXmGPyVZMs7WwhN2CmWyqRBVCR144VPNbrtT/G2sMFziyMsHWKqs+nO
+RMFsHtdOf+cAeou3ZAvXVXRCDNB4nGz9JuuqkDUvez3qLf6gpO93IAhhjVjdXF0QmtLQ7mvHMKz
yAU7VSpaNlvit2FvMEXmuYk7GVmgl7GIF60w9rOGzxJj6lg+gEEGZd3/5KEI0xAKdHUSFkkZAcAQ
QspHRUA3OWoeFJvNo71sJjlDuVcQPRIW5SwFzyIvwKGHQX+IsZUOW2AFhPBKQSz12uwaT/z3Z+mz
ER9H7xEAHTIvuHnu8cC/SdZqPz1u7Q6jWTq8LF5EtsNoKSWD90Q95Hunso3/xNvrc48OOkWEIctp
pr1AViZZJkMvHZ2rvFRmtDX0tbCF1AwnqQYBFAxiFnYdOlQ71kOoPH4FQJd9y+4MJNHVRFKATKjM
c54M1DqQMclnMOCQMCtlKIo5jUnxoWf5+0gl61nYLZULsErzZDuzyxmt06IK4iSOtNoqNXaYAG5A
sCHrPicn4IQSHHKCnyNWNpg0sN9wDuanPihTEvw1p1annOdoPv6chc/h7CazFYvgUQp+ccrNKTNu
/K4F8cGdJMs7oTJIhoWgK2JtfYzPqSCVZaxONZwyVUinZ+DCJ039OH1AJKaJc9hLLF/+rqEBzvp0
tyURJp4EPjL5CNP9VZeceDVqPcJghFI907cWOX3mtpy6fuKDGvkHL2Fb+B+WM7Y90UKTDvy4pbGW
ZY+iicsPaWDgbod6A53vpli3lVHLyHFv/uWpDZcWWT7l3xkHtL4X2zulfDnzxGeNvktnIje4+8ao
5jyJSKwHMCGWB+fdYCRDjF7Maw8Ezf/o/fXvFGZnzgmSoTPCe+i0HmA+gN8a9MyHTuZFOTt/qziU
9bqZezXv7gt4WgVa8y5+f6sD8Kdjm7t6K6DOEpbOtwncqEKiULAm2qxsk7DDu8NlvcBlmaKZuItV
JyqO2KcA0n4jWm5jQKLVM56jgfa46Qh22Tl/X+9c0H+O2mJo40aSoKS+SYE+swJCZfB/m9vAiEYN
QktRI5HWqY4FcsObWVUIFTwD78uKHUKd9K052ucaBovsudsUU21nvP23SAN3pRIn7oGXl8bU2l5o
nNJskUDbNNWjHh94QYQNeraYIs7svd251BRVvgH9kkqaGR6in31n62vcHb2iJtzKBHgbBJ4gguEY
ZM/uo9Fni5fJbaeUdZ/uBKbfsy1P7H4EDcmfS2AkulLsiWNTBAyBt4s/KTJkWp/W283cVo6UfgyF
HbqgR68CQZPJYeVjhBbhOeKPPIIMqj+xDbqEs62PvWKjzEgCCsmjaZC65Np3sQgxMHfcZwjZ4ewd
thWYMd1pTGXTBcfOeVSoYQbDfWZmGt0Dxn+FqcKAUw6ECmcEdkongAEcGl3QTdda7hC8tnqRtkrN
69t1C0ni+lhbr7vDXgpeVFaX4l2Tq9W9CmqNnkUNPyW05F2/M0COYpUG2A9SjTeQYe111yjUlslQ
j9EegcMZYnuM91AZ50RWtYBilSCHpW91vzSQ+MRgC9XFV7vIE0lpJo1gQ596vGFaFnrkA+AcyloS
JPYmnBr+dFHSJGngKd5Kjn39ZRiuSaklAOXcxCH+vc4rnrtsTu8clSekSHCKTUYcFV8BhA0IGfy+
4UCN/G7lkhfBMLHM+vel4fjV7izaaabQl+pjUHk8gM8tXVI1RRJNJW9tWN8MI5f/LR05k2q2hCtn
JN/sBqVLgMQr1FWqR4xz0Fl+hLSy70uXp0MZdzMp1QZshxsoQ59oQyOP5xW2aXXQFr0xFBK1r01d
75mL6oqC+oW0d3+wMl25KIlQY+DizaqNkK1J5NPhWURaRSiM4UfJ5aL1CReE6DTzhOXJNC8SbF4D
qa+1QoYvDIPF2OO4xlSL3Fr3HInhjfXkRi3tBeKx7VOBLiE4LLoqM4LxbS8s9UyGBwYFKwUZ6YzB
2LcmEJANTzHDBhutkI5pWCB9SxezqfB/msW/icnboW+9lpAndU2CdAL8upuhzbstBEuVsr3AZMOE
y/ZDBBfVJTguwsrVMxqnhQ+X9xXrTySsPNokC+iSQO5nimeTbNYNAvssM6/PSpcFjvO4DTGI3IMi
mD6WdA1xQ+y8oKNtdvDvXsJGeuhQHJQ9SDliXf8VZXialrbk1SrBGfQq0krf4g7FfLd4AsfdjvWP
82xF6AWg5f/9MwMrCXarE8XJZSTRhQpiBrIwJv5cMg1e9sVwvykRW0vb9jMsYiqJjmf6420hhd1S
R7r+4GCPG1QoPp6TqshA5Zc/0p+jZG1/yNsn4NVVf3uh9tVZRjjLPnE02uJniZXeS2Y3dGyUBK0V
wkEerMbS7KmmAb5EaYMarFZbfm2ryA5YskJ8FtcFm2F2ePEghd1KIXUewqK29wN8nBppcmoznroa
qD6dtG4TUqCeVoOrt9DNhvL8obDWxtDOUfJ9ew2B/Xl4enBYPfXes+j5NbGCI59UQjNLTkivgbLX
d/8wAzwlmWTsYTXYRLqeJcsqhs/V3ygWi9eWSz5BftmwFbIebF59sGvSKRVHavMAt0gf8+Mee9qF
a+WQHqsA3VrnTrkYUaEt2t5WoPJnQHIN/LgEIT5ahe6KLyjNWvMtVtxmruUADyuJVziQMKcz/nWZ
ZcQoaUxsKkP/VfmENPhF/OugZVanVS+kI9qN/6XfDw0BcsVPtqS8YU82TMZ7gnldL3ia2GN1fRsQ
3ee3cD7sn1xqInaJmr6AfR9gCBJwOKaCR2hUJaEIDaXmMCTTYvb/FZagZi9HOH84KkkjOtylkCTn
IXZ+8jL7CJF9c9bIaqbv2S/gNGEnbmONP1b78zCxhW0xAPL+VsI0dxzRJ2TMJDsJr1DrpjSikjUv
28iwRqcVBH6j6MH6FP2EGib/OkRDxpt/Z/jrlSIWCAa+UPLbQ+X79pWkpqS0HWxn8hKKecN+i0/A
dci5LlHoVg229pxMgby/GbrKtnhawcoj4iy7BHGFfPGQYxfu81+Xi8zCL54JSm168Tpg85n+cW/B
q11rmJ+bigqtpBEvln4CzTTFgMmISATsH8tL0387c3rFsDgRYECX6vjmZxuOSr+VxdIJullrBPys
uvMzpn3PTwc1MSOBEHJ/kgkL6qxo0xWytnra593ZS0rPBuLoL+567U4hRRTPgDdzuiAFAUnudeZx
Iic7iwZt+jycLNgVG6zaTvne7eBpbIZW6T+bgvuo1gJzY6RYqBFYgA2i6Tp5aBiw/O+X46QaZ7VP
Jc9WxXZwqpxR9UH2TmJCfGBqs4GKMpwcLxPshKUXUH1iC6SVAI6ZaXS+2kRaI0MbpLB2fDVwTWU0
kXrY+PdaxNhuxp9/iN3xzc7qrBJJvh1IH3wM/KarBMFJulGAJQR2NUiYMZiidVi6uTmryk4pYVGi
fhfPDUopiOUrKlX+7668+XGHwCZV171EQQMDD9EMtr0yPyJbt+a8Si056DjP+UVlSVjk8wRs96iQ
kJRi5eOi2w6fFb9IQ4atlHuZtCtXuOIVQ7vMHPNUIqOhPJQ8icTCboyfNLxlaKVIjI9ztMy8WXtI
oao3jU6bXWTZmQ2/7osnAc4DX1hxfLxWrq1GYcsRzWfda3hlcw1P+vax9I0vtQOa2VKErVxfaN57
d9CMm/GrJke+qGTeCaXISNXT4eGAg8xUX/7TxrFwmRQW7RnkLOwOodTp4FB2z63l/zgY/xZJtnsf
vtSbKap5FoBUkT+Q7HDGwZOWanimFhOQS6CAq+ib2U7dKHFMidAcpfKWWuTYpsMGqbNEpgvpvC6F
cXNSrGcIaHUF0eHLsqOFOsQBCnx+l5Zb0158RUrNEWBVJRZ7qkZXpZTJbsqKtoypRPbnJgSh8XTZ
9VLCZxYuQJt7c5DFtb5fmPnBUBmYz3HfJh6N9J+qdY/tPa5emZHblIF7IMJNi0ityTps3JIUAWUv
Qnhpa1KZEtJ4tx2ag7V8LlgT/kIcs9JtHFYzgXv3tC037FOiazi69/LOiPM8Jj4+rkBm9TDJfSVh
CIxva0c3vHfpUZUxB6sbVvdC0KgzHUrlkxc1AM16BOqr5BsFeY8KPuBiqrLCNjA/s4uJM0LfPDAi
OXoQVDjYPGQHE706xm4HS5pOAxqfKVht6wLBnGus7cZ5j6H7+X5l7sSHndyemwU61P5jqOq6LqdQ
6tzg4fhrB6ed9okrmVe+euwY7hWB1XNvZPgyx5ugXOgoxd+WP2sxvjIWpvxnREgfgegF/FxTbuoK
0lBhXhsq7nsgS4w9YVqiiXE3dBMFJhr9KQN4LuCoEsQLU3TKt9wnW3ngqEGPWsZuEuzbFGDLv7Xz
n0nHCeUQcWmbCiPo8W0w3XSVFruSh76gYk3lAAVjvBP24okvzPr34dN0sNoW89BsCBgBukjsu8a0
VoZttSjVyEE04NFBnBNMdP6LkBCwd4H+r9fC/yg0hojINwWSvnCt7NMIJSTMtkB2Pj1DnlIAhigb
JXUKsfSWHkTZeJwWLfqBbZEKoJHhDQ7W6S8Co2gS//PVtmbnX9qlBNvb+NvslhbKHa96YgEznkg5
+ErZpjaaTXHuTZDP6zDdPRFFZi9ASZTkyCvWkqwDtDRRDi7Z7KUx9XGePxNaqjsbiyEdNSa4a8VC
WipqNCy0CrqLcQdFxwJLMCTUjNWQu7xzt6wLgD+l4WJqiWdrHR2ThUbN9+wcFh3WQZNLJAFpIS5H
0eTepAM2EVZDC+D4yniZkPSZMjR5vN+USUcBhdpRUZdgeOxe5/tnvHk5tpacVt4ySgbX3CFmGoYP
Z6KoD9lohkX4foyCyWYzGSbX/uFrzn+20hBsDXE1vbeoUYn8i9/dDC6c/cqHExzNam+VcHPVAYAm
CrEYn/J2ypxBxz9RZPpAk2icXo8tyfJFHYY6nVdYykspip/kYbqRg3XQikhyXmAug4eJam22gZ/I
hP/8wZZsEcg9K/io/Q8p7H6u751Ij4LvnXMXzlEMdxltgBfobULpoAsOEwWPuYV+pkz1LLNm29xi
CuV6y+x6XcA1S46eSvpWK77VkG2jHAqPfEsXBUXjaW16wSQ85LThG08DbNHTct9EYj+gh3/hHUqh
ku1yVUHJmEQyvsiMay3cLZazauhFh/pGD3ZJhFJtZhhf6qiQawex5Vuk6LbNlZRQCVhEaVSTSU4L
R5N+chUjPsRh0tAXDZRV2FDTiTgK1pq9KkevSV/kcLQmDInQWYRaIUg3+znoYgtF8hyavzigTomu
janOE4cMKQ8TVWAvQsd+ZCsSWzHPYnep8BClCtQIyEQaBglW9ULGCbRq/Q1wdMUurtXB1T+wP80b
C3ZQ2vXEBYWY3MApE7k6YOCVBYYEeEXn12CFSdTX+/VLIC7Z5ugnc/kRVxr/0FrjBO1msO5b9txx
ctG3qAh02RQe469FOxkEh6ENcGrDxTD/VcHaUx7C3cDhj9IB51aKvmD0czlhBRB+abn6H1/v+Ccm
bEf92RwtFFFICaV+XyiZzlE+m+jnG+Z/Zw5MaD5fgaF/UhZaQ7Ntf/UZldCVr3PTh1vPecq25Hrv
xLfApgHv5JQNHSthLi75TC81xkAvvI+j58nx6t8bVfX+PmvL36iMtQouwyPz0VXp4LT1mR6GJqZw
NsAW9sdPHYnSXULQSiccK78TO/vEQgamIcel2LP8cMwRyr8eBh2UtJL5H3N3I2o5eE5lcHE/vwBp
aOwy1ZbaMdQ1sG3FKC2jEzWX4o3c1I+KI5f9g7IEBARI2kTuWJPjl4mkP8nRKHOIr1VUKvmXqB4R
VvICiC5dUXK/00XfgtvORzzBd6d3a9/yYcpgZtzzv4/bw3qDDVHOWMDvJPMzuXLqnVkbvgyL1WPW
a5zasheSYNcHxvqv0o4X4JQoQgmj1dynw5fjzIKjbS82suPo1uiAfCQbmKdE07EC42R2THZ5RXQq
Pe3MUXdecUHY6ioxLBlKs2lvCslTo86iSoiB7XVRf1Huzue4Aj0CGw8ETbJm4nAVXJPOcTaJ96PR
bkZ2j7x74jIC+p0x/zCQ5L/88dTRbSHcrd6jx3EShrMayUTolG1NcQdUb99EpaKpcEHjtP9uRVvi
3FU9NoVShAzOfv5Axh5AwqEBiEzsy1ytLxLr2sq8Jc1Ra9JiBT4YleQn0OxGrXdsTcRM0Nuy2ptt
qGP7a3jMNN4CPfCCP2xo1012kw1iJ1WTPRABL1QGAvYPtGEl73RDZuTRqsBzOCvXMQkb4DSZshNI
98qN46pC0o09tOVMJB1BI6uWsyjcueebFpNDMbd11pUibdrKmEsVljCh+JBxp+1BPcJ2EGWRCoTJ
V/3mmWdLf3FSY4sx7qf9HqR65gcWoHhv9Bo3MyXHhLYpAg8rleNgkB89oqhJNR30Sn1hvLbHCvX1
6XX2/cAaWW6s7c/rYKtIuWTf5OrmvIO/0c5lhPDltv983ELVkse1IqQdpQ9sUlu0aAuzPmLZmdbi
ySeMpY/veYnXGG6IQ5wscZ4DqXNnOX81FTbnBfS4uWGBJJFFH2O1/JOfyOUCm9eNCAWC8jU+UgXz
+/Pr9MteRHgbpBmRTq9VgKsysHVSGIVeDuHGlQ2ITzepTYQXQkbOELRJCOgt7O3yQXUI95catYy6
vsojD2us/c+9FRSo00/PBevRCkSPIydwKe5dhnu5StpVmAmQkGLszmUtIE5k3t2MMKxr5jV3UDeC
m3OPtjZnTBFEjuEOO2Prs8VGSpdsowqUoqt63Clf5dNg4alRJ/mwbqXn671oka0ZwmOoX5wOlaLG
KZcGUJuEPlxwcnqHommi80RnED8QlWe+r+kvOEbm3xW4f1r/MNeOAh7TrcUZEzxANkCEcA05asO5
kMy7VGGOjWuzqvtsNb7BJ5PCys91SHm+RpFpBYUR3PsEkaxppw+lnhnjt1EMXan1ql/FY9BObitC
0bHaP2t2O7UyokFIXdE0xc69Un3NtOi7paQ5AT1cuvv+yH+DVAwY+PUjfwpYnzkHOsA5GaMphGuy
7t7D65FDqu0Lq1mB7AaIKZCPw9JGJyjGQFNrk2DVgnGjUwUNL71t5RLUH7vz2WnkTPA1jPFi7QZH
6WFwAC8f3W/NA2mZGP1tzv1ZnTw9w3pWFO/x8Gp7r3M3WRilh61V6RSndcat/QL9ZTX9gYB/msz1
EUhixvzuO0QpnQxABUAKkdZDha6o0JqGrWyZV3mihtjN9MifLNvcOUjXAelst2rCQU3AkIDDVkhP
mR3DAd6XOi7r09voIic6TtQaEBNO7KXqpztn6UDZ0u9V+aQvqxgyHosJC97xll/dfOXX2yFONYAw
VLXkMR1ylYS103HUDCbkiwZuA96ozMgFgCnGVKNKTxozdyYQO7D0O1qC8JWOplbg4cHc65cbpd11
ZbYS0d3Xes+RQlxHC+nu8+sag+748gcKmpNJPNdV5a8ymzqNN/hdJToGv1F3STKnsk7/jiSonW/8
JTx0Ry3rSzjgj50MzZBUmk0+Yqx94KUo6DUYTUfIkQaMTLbZhuzQ+Y60lBcvfdPpDdF5+ndIJy1q
5zpOVhAguXkg1d6IBcl15s/1+yAu482Z9HJt2QVhQBoP9M9OQBdafdx/t2W9WdLaRnTzgeea9ZJ3
iWGxOWBt+PHU3vQtWk7umriXz1Tywt8j+DEFywm/q75TNd9NwMLAb3wGcPZhJTG2KQYjJ8b209JO
gpK3Y8WTEw0IoI8PAB21Y/ST2fhIV3bfkMJbD4+rinqpjwvYlZ4mqHHmpGfNDGM3GQRwUG+TYzP9
kM+kukAazm8OHXj4j81qyGZLBSnJ21Cd4E8Ol16Vo8oq/P92i1/KyRzqjuAwmFKGOmfRZsLegD6o
kk2jE16rtgyvX3mJqCG9RUqBMltPufQtCCkAeMfkPOJ4o8pzOtC8aJ2upXNCWrvdg03bgBvOhgpm
QkASVY4nMSr1wxRxwGG70f2Dg/p3uL3fxI+0zN2rjKhWaLx8YkIXTkgB8is9tnIIOprZxRg2IbAH
MREwyVIPuRoY+WiKbxopEKJOtzQIVWX9ApbR9VVN92Nm0WM/6xMb/XEN7QBLRYcQiMmUlv5hKd6L
dPnS3XC8jquJ8MLEtlfrZL2cnHgpsIWIZbXr03vY/XvpN+I3xaNLbN74eSuGCAsS/N+00pBmY9wy
NVItbK3SNA7WF4UNEqbrsY098zoL8g/nO3kd3sCSdYH71IVdUKnAp77e5ix21+E/jQMQVBlO39So
3ylqQweHJnf5geSm1jWnOhPqjJUK66+SgdGp7EW5trzhGzCfYb8qiUEu2QzgeCe0nUCbDONPUp2/
QKJtUCDBJpw0bafScXHgn/AyoeVFKwzkAnXrF+FOufxyrhYNQvgFD2CLNQ8/Nd8Pw2fxK7wQcacW
Vt5HqMoOziL7WOdPz3L7B174L7Kzb4wgHhoP/QfFB3Rm41rofzroH3VDwAgcUV3SSybk7+VsW6LS
WRxUnivCFYzf9Tn6CcfdlwE+0lRfOOEqb9TumWrtRx3rfLkJbBa1TcqDOQw70EykeyLFfVkN8kRc
XVTnXKUR48kZQGjmLeCXZryrdWK+T77PQGMyZPWlOCDzekX+LGWzVb6SqkFrcdq5q3ynm7i9vbgw
jlcZQZ8WVJAvGtPdXvQ22FZYr7SbSAlrYO3dm3sPvRkc/2hmZlbXpxZBs1tI9PqFj8iK7kT/xHej
m3v9tRm+RK4L0Lh/n4GR9dBISW0RpFDt1bEf3XlXSHHesgOYCKvpCrl3kZHlE61BxFWnafzPuMwr
EmeLsKcRealekrqhzqomj1Tpi9MuyKGuKMucQPrcDaQQ5j6TEX7vtAV3EY2Tum3h31zZN45wWGRt
CVwJkWMWKjRCowENVL/BEuMiIjmVia4DZrOdz5YDRBZOFsVsesXXCb6y9HSz48KROIApw1rVx4Ty
oQwEHrIAxRiigLVMquEgoh7oAOU4DiL6tJxefybF7CMF/VNYeoG8YUevY1AolyLxN2SvFMm28zpT
lUj78TzIAsnGabLhhpGscKHVK45GFLalooVAEL0+mMnTLYV9h4bOjdK4DFr20dyhf4sB5FSAH6/y
2MHKWdZcQHXbM9Ga/8Zpji9G3IisNG+QhhRgumn7LtGUxoyH7EF25D/0BRcRa9OBxFB893vnZP9j
lKti/uhJwvFklD4+0IxVV2UQEsC9HBHGrqL9eX2rvre9eRFbOtyUtEf7oQwapunrfMDZAafFjumy
xnkHRmmCi0s6b8BjeASHVC513UupFaLgBBf/vMgFH7Pp3ts7FyQ7VRHu10lKMavYpeIg88EW/cUr
9GvQi5ZTCsxYWC50qSj3o0RCfpbK0KhqvvgG94DUNzpWxX/XwQQyHH0i9KBdLOK2CkWW089Uj/Og
5TP6kvw9avIvA45028h26beNwgrph7NogTJsqLczF4lVz+J5E3ckyeEUD0wR4zXMxSnzSUb0YkKD
2Ha3tnfB+bnt+C/ZNXqDilIqs4W7dvIlOTKYt6Ud5HDUxtQ1/D5mL6KS/SHmFE/aeWZEGdpdts3s
w4AByP210KGuSwJinQh/rgvE0+rWdEonZiMZyZZa7vgczokmqB0iD4I4dRxwS2EUaNuLXFwk4ok6
EWvwsbfJl3j3OpOKwPM7b+44L5cqHbmXVTMbuv4jLGjQwJDxr86L8+LrZ93Q6/2CKBgmALDtJtDt
U5w213DkgM96GSxEBwIaRhMgpkdffW5eviqs5el3/Tzw2IjgcFTmRf1eDrCM+FxyllhKx+3KufgA
6V0evWoHDdYy/P5JDWgsR1BpIe4Q/pZk4vhbvEwxwmrTMx5E1leQ9fHkMyi8n+QdH8y2Us/cUTkh
uJnRaBnMibts9VYmGog6tlCfc4MXwKDE5N1/MSrLzD+kbYB0xM50PK53RV383ZLzzznNKHUFfhCd
j+vsEaKGicubg0IbVKwRTzfzw17xxwv72oodkypYT/vsve1VW3lKCNdhaqfIOB1il5varRERe4S1
5OLpI8YQI1h++v2DVWMMxkFcSo+ePalZi6/A+VtRWcSfW4ckd1zzu09B4k53+0rJsU/ArhL1+j72
gZhPgsQRrsM1HeCHiL9/m8pELhfpLFQG+/vhYbySMGJfqDl7OJFNek5YUBJT6uyqCs3NMD9hl5Jw
DkP8fGYAjK4mokjiYNP24GjPgZwIZ8ssHLGlL0zSnfWfrYPyE+QzxusgbL+/jXDen22IDT9Nm/fW
47orWf6LxG1Dr29Il4Vb+OJOnUlhhmeVZORjRjTC81bEp6/G9Iu6ofbFZFW23qfvKEPEYW6aAyew
gBwGv479uUUhmJFZh+7vEd2FlQhAT5j0rBKuYyFBM7ijO642UDGWXyv3HINI4LKBPi7OgYUCL6c5
Wyh5tDd3vVVI3Kul0ZUE4s01TdvcGngtupIlyb5j3GMBA5L9PqcDV5tlvQcy+grLAYMFuapGXVMG
gVnM00aFC96pX5D98hjsJ/x6gtcMN+sPiCySrbn3rmoVo+dAvYnSZ/oGF2WrK8wWOR/9XCAtDN2V
vsIUPusw0VK5J9jBy5Dzi5o9Edw+yb2LkghUgUFAMj8/ZzFGQruPS/lUdinDso5UOVyYMyCYUu5N
GXysv4pImzBf1ckz3DoctlaoxAYQaP+Lumnz1zAA3NLB3uazwHrRY52ITquVmnmMoUccjNs7dwNh
CdcqF04BdOxaQc4ohbZtOnskYXHmSBv5Xm0SkW/RRJh4TSgOEQ0qh9I4wxPe2FQhD0VTQVD4k7+t
BmRaYMJxKwz7qwh8LK+AeXFLUbFdNDQ6Kzb9tc13ERBNzqJ62BPY3TGld+PqcEK+GpIz/7rds7v5
XBF+mzn3HSN7wNd9O7yQ8VpoOXbfEX++sY9xkAdzhPc51nxXxUWpxJJu0gfJwsEdwIgVkHLmaLlq
QxNZ61azONha+kRhSvKfASalwNsXQifg64j6cZH6aBSicHbA/GKpVKpMdM/w3Qn7fas/t3J7erah
imDMB12RVVf0KJec74Bala4f26rAgtdXPaN0abuxYUubNV0IzoBkMdJngeRMjCEtV4BMUz5rg41t
fnpIwoCfk42KzMyXVSgqBRmI8WtOPhFQktAVWkY8PTCCIKTrxxf41wdzEuCBtk61NmHz5XkvMeUF
j6gtBYX8Ro2ZuekhMdcVPq9Z0wGWXpTvbdsaasNS/uaKZGwl2lJ/GAV9pL3EVNAEcf4ttMLiE/B1
mVchkgUnd/ftHX5ksDcjWXTb6UWFw4LKdY6/jZe09BaS72S6COvZrrlC5a48t3HtFzCtL5tX8ePz
mznzjt516597hZFRFU35PgS/CgJqHm+ixn8jvDnlbxEPgSYtig0+Wv+6aCpY+LN6EhY7yxQApR30
kSKWBfmm2o4OxtD7Q+q+v8jpGAvAIh9Jie8jLQbG1DpxKuBjGDRSLbOtH9UxXF4RTjiL6XljxAdt
AmcPY9/odbd2Fv+JCz/Pi22amApW9D50gtRIE7N3J4t7T3lKOb2CBsUNE7igMgmQZ78CBTa8i/t/
718RXiamToBQyp39K17yTk4ehsg8fljkhHeq4urXW9QqxO+wsjlabVGdvKJpwb+tWp8D5alvMn1T
ePqr2WTAD82M/P+REFAQWJoIeMYlaZuWcAHSfwxuAucFWMIQ4vq8U1p+ceRvvqrdVaJgpyRCN0I5
3DzO0aowGcQ46CTzxPOOZywPGy97orY0kok8zTnHhJ3SwxrvaeL7riBo0mgShpWy8nmqrlSyddR3
fxbFMDpISPTPHhdShDeuXt/ANc0lhEFPpUZMogGJTXGbPDhHIDPVgm6VbSbm/WwOzOEZQq/AmWwt
MCdXfUFXRtJgxfnFEjEPT93zV1W63205SdtJhEy+E1mFBJi8wrgSdXkm2JMLlDKkyDtpQU3jlTrb
OqLsHOw63aKsHdWW6ATfSf12O6gIEHEkmCkD7bMt1Q4eF2Pr9AUzBGekq0xTI7lBbW9RfIEs6CQA
lZGfhvmC3RVjyguiXp4Gh3tTJq926T/WbYKTfpHsiAQgFcJKVFase+hVOhY8yR/sa6ffgRuUOZBz
PORJPB0jG3eaXx9WqgMmCaKfp513nd2Y+TshDDU+/47/Ds7ykuvXiT14+iv+JA4dv1EUW36A5U5Q
yRuIueGy3Iexz0XxVW4STGC0qjukmrzZKKAbNAJ4kF1O26j9utFxn1shiN8GHFk54s4deKgrz5zH
2mmW1/0OF494WSCsA+Xxk8XicULvai+V0h8XWxEf2fJ/IFslExxyH5fYF5oFiy9CLkl7CkTp3c03
bLWe/3G9qCzLGAiN1Uo0jZkVuCu7KXk+CVqIURxhW8bJrOLyHA4SvF0bZcHCkq7RNV62xmyXDw8n
7UHK31QIbsz08SMYeIYh9JbATkmbnuwY2gVrfeEnpxJ3gdGGmHAZB9VhM5mZSEeQJLHDmxrJ+vmr
5Tx1yk9h2sE33v1zcxKYMUvY2ckbRCEgS/iBrkj/PI7kKrElkKk5O2coWfbM7SnoKqSh+u47kN6q
1wO2jO6kcI72PMO19kue7QVBt8P2Nw47VN4bYXt8atOhO09NsKZALhEu/cfckMXucEADisdmhhgm
QMn2LZqTG0w/vpwywyQyowSfx48SkLUJ6v1seFjCrh5wzGJlx1r4T5SKYx+LuXlFdxl2AB5m8pZk
4eaS4SlrXcS9e+fJAe+VJf5VCzwZaimEB3YLYt0k3dlagh7adGQieDTjZrSdILUwm+t8ak+1s+QV
3ex9JK5SIfldE9zf1f5xsinXnKwwxQs3C5sDGJf6Ehz4RgK//bl3FysrXSijGT/z5c4saxWiKfFQ
iTqJpxEE6bbK1aOW0f0PfSeMUy/5Vx+4Yae/HmpbZ3gOCyJYOFOBOQfD3b6bVXs3wzHTWch0XAUT
mCGl33X8/sFG+G1liELZPrf/COFgNLPiQ1a2UZKagEVaYPx6jUpCGXYXZaThU2Mfr9ZRHATjn8bm
BQ7pTKptDgPn0J3UoAaF+v1iPLEgjZXDndkkjvIcCoqR41EsFFgx2xUD1tNe3Blp9heOIMfI5Umk
WrR4k6SydAYz1jhySODXzuQCHIR+vB9JhTBWHQcZ9tWe0ij3+SipJSkxkXzFVMTOLOZGcrMm1uq/
C3CFwmAs3t5W+Ace2LxW5lR2QvOMwFyezbCQ1xjAPBkS9V2EwkIcysyR62N6KhP5ZvUwd5xDSUkF
GSmUmvAZiGKEBPEfp0DOaLwPvX4fkrdxHyUGmeRCLqfO4kNSiCn/vX1sM35snwLZS6oFh5Bp8hmC
tO1RUQ/DZX5mT1Vvgj5QOiE7YGSYsogqO5hDbmwrSBXZjrF17h8wDtbNt0SzlKcKEa/iJ8neQ9dK
/4lD7aCwxDvyO4xTvMi0Cesq3iypEVDETnhfy9Nsw6lr/1mUOBo2kCek+fzjr5fvNhYeP10gUCiE
B2vaQ+To3MsLZfS5yBXSxQGur7kkMYUbkyA67NpPHl4ac/gk7UtovTqMJVcy6aR7BpRfKbCznNHb
MTBq4agAsbNNVpXPitVUMEtGuRfhaMARG1GGS8aI1sw+3rCnrbspe+fclC8xtgJhO5mEB7CmYbMT
kP0CGztRyscKIxe2HQdJkS/S+iCjZTUhjqW1rcFLFbCd5UMJLgRz9/ZuLr+4NqHaW25jNMceL7st
VH8d+ZLsoXMn8LvnUwNij075UXyuJTAHXxDVxFjjE364YHw27KmUXvJ9swQ+VcD6hRsGH7WXseeI
pL6oHDzVbADb4tFwf87/bUsaXyMINzJcTehCUQ731XNjhP5kyLnmGxOTAZJDMoUa8YM/IvViE2HC
jI5b6e8nprNNE0CmIu5M4xj+fimH6BprQ1DKqPTP9pgNNZAsqetYsUtzaUB/p2/QSDQ2/nw7jmwK
Eh1KLVG5cWWxd6XFD5ub00IRzCcTemHkyBG1R2Amd6vVWekyzctjkPw1xMcek3FwwAN6BzfxGziW
+vTjVsizFwwKtcLs6liS0QCkHmr2dcPsRLHOHE+QM8J7CEIQNqQ4TYbLX36Y1y2ecZo+qdwNCSyh
Xdo9nZeE7W5LpAAUQxVW5Pq3J7ZNnI5i3/hgUz3kwV9e79GD42Ckq66JwzUNBvmjILeVYUR1gief
k7QMRgg9HAQotGRTt6iENxohA6SpqE2M/YRADq2nsv7A0CDf3XSoUO1KtXRp4PCwVnTtdG7BfLxW
aPSZLiHVEsTT1D65zqUzh65+/dzV6ewMiW3pLTKXn2Dy54CIh0Lfk6wt9GpPvCt3i+B0Nov5Son2
Q9eXD1M0ppOwi4/GgtGSkOfg7DL4IgnPch1cMMV0NH7JoPv1lvmT73PTsBsywoGcNxFrV6n7uNzz
8u19oM487w0DRQ095qpOmWwHcd5bw+Yb6/MU7nx+xAizC7UMeQWjT4Uh4l325BD2VHPwJLdR2cdp
Mp+EpZcqLigJgGlse6JzND811pFpciYvAv8guZpj7ZUTcnuIEQA8yebVj+vARKmc4YliE5MTYIo4
UnPF48YWBzRI+Z1LoKgX3i4PB3Wku/SEF3N9lzV1Kp3++vVz+hkmF3qaxONaOgWEyovG/nt1hCOJ
ynE/gjIbqcj5rvBsle7KDVei2tSr5dFEdfYMOv7kHGotcE1oclpJ+adqhKbHXRjgnodz8LNzdy2/
f3Qp6jYekHQ6VXvxEcq6q23gntpagNR/YoADcyRCpqRI/hyz+YJPXvU4zdV6xbGcWO7pdYMx4Ggg
SU/NKNCw/8dgU65oSlQkD3Vc6zSJbxRL5RbAPSB8M5naiT91AHqCVoeFCHT0SiB7kkd7w28lezWL
+8EhhUQiuHiA8EuetEOvpnTaeLU4X+w06wYSpxjpkurxworLXxBMWryPgZu58twe2uRnh0LjD1cx
yKxJeZYHkk9aQ+6Uw6iuV52v7WNfOINSPtJSnF96i6tDTX8JN1ppBWjIKVHJvuKnjkQa5+HT33ID
NSxe6brHl9ZFPImQ3qzbpd4NtQr+OwlTHOnQOuxLxe9cNL0jM+UycOIlUxh2S+5f6bBuaFC7aH4t
MR5G/6DQPhCRnnMObILLen6l4Dak21FzIlxUDm960ArpQNybtdURIqJlO+GbVmJaWEuRizXJUwvC
Qvzr/lsBIptI+OMyj6ZDnEtNUyDCE8DR2TyZb4Ndvwb9KlrRXAXODkp14vFI8vtFOqIodjjy33se
3d416HeX00FGvX4hgzS9zY0iYWeh1+PxQawhpc0yPajGnmU1oMMWx5Eid5CQYgQ9X24UxhwnokDX
2JoUT1bIVxiNpGlbG78XrKMWUk1QydtC3KOmUC2JdMdI0Ha+7poyb6EGAQfY3yyt74bsotNK51jB
oSewsuShQwWal4aG6o6dGlP8HRmGQrnDZCBKPW1YVwa7hSWJY/5YmiF29aPTGbeRWozzLFvTe+fL
IzcgARQLc1obVk0ZpQbHMRrjLJo7pc+0j9uWb3iGeZJktpu/yKssTNHnpnYbEGa8WvLD5kgdDt65
zVzojCCgrQfPn45+5I4ffosHm0bDsZR5qSdIdLFtxQeAqslnZfuEm+WPTIivcFmeh5BWK2S1qMqB
ohxg6li81GsZfaiYmE4Cu2DCAG+3QmgTAggB00ldsurqGMUHy6pvsQLdh1iczhNAIQdmVTmRXWMG
NCQRCEwl5jSZNTAzBolJW/G9q05GSWH/hMXNxw39HBxbOSUo7hc0RDPtn7t3bqpcaecJj5P4DZQL
kJgR/Lx24v3FgNZKoVATWOC9noSslN3w6x78vJzgzhU3ZQ3gr8v4sEu5bX60E8eA8MtytOAKMUDa
Llx8Nsdtkol3IZqNG7K85Q2aULLFslvnAUfBlMK/crDDjcPhoCnPte3NQCotpvBvRYR+gH8mmmHk
l6KRP/Um7qVH6ZWxJaY1f7qSE57wa6wJofmgSX/r+owvi1UO7pXM0TZezgdsd+A5IUWVrwoMFCPk
6puJBGPqrfsHO01WNZ2DL8Nn2hWdc5CJJ2+vtLppGFZk8XzxG7qwCDe97eklQlFaCK4PUAJp8VCE
snrgz4+SKSll3AI+K/3+uATfbVJUoR6cVn7OKMKF/nEMC3CEtjNLslB6d9NlsittTwfrfQ92k/d/
GquhY8WCOEZlF/tbR5XnMRNKwT/g/wNPbEQffav5s/Gq8jZwgbbnDPyXy0fvLvhhmku4UUGtc+zh
NCdp6H/zK2az0Hu4AHqzZmbSC3hhWW1UuCi4z84gB+lJRQXG6HZpwf2CnAOJj7kpdhrNoaHb2L9t
bP1e3eHQ1scWIrzzzWwQtRlbgetbZNcOv/IsjDpAG/HPK/GNsorp7HTfwmg2SmcPAg9mQbW2Qggx
vrtp3Dc+7Lb20Aw8XT4HgRINndLUBByuwul82dHoKKq1fS1R1DxblDopPunHJbgVFCL35q/0gQ+s
6BFRDemGHKv4rYX/e9EhgmCxyEhu3s3sXUGnlD2N+rlh3WdodsBAgUo46DsqNfHOeZcVaCoRzqU2
gFpN8E3kddC/qhYVf9QYk2ZbVsxNd/inBrVHn6CiNzuQBawsdPM4cNJbxjeKQSUmr9jasMeTKKnW
fQKoO4Cm27sOkKRWQ25VkV9ioXcbvrriQgztQAPyVwxvbvIKihOpht8JaqWWymUUXazOtctUklbM
d5CbRgGquMpjJRHn1jyUUnRpw+2Kmx+jiygNOTfjE8nNfZwmTh7D2YB7qKB/IJxwLjPd4OQOjKm/
PoNErP3iPco/wvAXOmVRUw4FVZUVcoeZs2vv9DnKUd9LU3dLtJs064HPgx7SkUZILM5/91oc5cqN
UdJkgrD6C8MBawXfKcwFWoSNwloDlECLelAFpRnLrB+XVfUKKWyVQm2PdDVoSm6fdiPAJOP0mEc7
gFDbpheGzoSiEqjVjzIcAYTGdaKKguTLTHVRbB8YBeTYyGdKWc6UA5rxskeMvHtQtRiOSDCIprcG
WJEC8FsBAZk6C5IVQpn49XKzQzWzOWj4Elj1+OR6pyEmS/fi+7bZTePi6Qg4vzKhePkJu4bThAkJ
VH5O/zNbvEQmIRdtCpmha3lhowVEBJdQLvAKqZnsV0X6V+eHw1bKnz0YZETmKkCaqU7E/8NxUyuJ
pFyi8MRaJm1TCf2jsot15GEx4H82XjJdtR/nUNBvnXn+bPFujYn5ZZrVOCNFp0lqU0f5JzttiJXZ
XDdPsRp84tusL+zVLMHeL1q+IcbJmGDuEGHaT+vLEkyoCOnF50xM15SKeB/A20HCcuN8ZcRMl4ga
AsRmLG1pkJnahTvqW89O3yrQ8RefrlKSM73cLArWVBEGt0ljTrMLBYbWrco6SCis0xY0ojW6aSJ3
b9L35aNh9eVvMwIZFI80LrET1Md04ibOkeCPZUGEa5YJBbbSHXb1BRwScbiMUmNQZqRKIVajrYRd
6PBhjF4YsG7zcmtJ37qiVWbDPiw6nz5OyxBldHbmnbAOfIMfvCMBkhvTem9UWUfN69bwE92CB0me
/+uzWtMZwbZRX7AGjf/Zxzw/d8Ytiijg2Hzs0X+VnQyOKiMUs+wXc6lxVbcSl+qNKIgZ2W5SxrgV
DsyPosxD1+S7dgWZaY33RuuL3/AaSJzVSuisFsXHV/62HwlgF20fDGqy/Jb/nsbHxOCbPcvhzo4J
Bg+enAOCD/1Gq4t2hwic1t7nQv/MjunFDa8jf5Mmc0GZH6zn54ImBHkb1YoE1BgwFTdIsvOTzIXW
XczWTx5NmyUOmHzwFWG79ZcHj6abG158+XS5tdr2KEv7KIIIdv0DKpifrMLQEq5gccjbu3hMdul/
SgqtXU6AuHSFrSYFWts4zswi3goytYdehhxPjVCCKuOG4f50M/yIh79akxPN/kQcAHlZXjjxSCGi
BXXlJDbHmyrVwg3oYNFyBfUkEqUGirtEcPm6WpvqBKJ/jE3konqO/kyO7SLvMRrPHkqo9kJ4IDgI
0qlGLzr0/V0nL0M2RDFpfsnoi9DSONoHa3onqEpnKjZmcdk5M44CM2JPRvnNGOY2DTsxNa3QRqg9
stfE59D/Ek3celmtHgZibT4XNAKwi8y3zKUajPKlRfKaR1mGv4l5z5pB92inch059R7b3OL/Luvz
ylkcxsXAhiHmLW8JftMgrSLW1MehrMKQudE/aW52+2vQld7w/EEmR/0OacU8uf1dyCnboMsil7l6
PF0Fb/2z3RAadoF/KBEHD+ntXaah3UZ3crsHnxVvB9xh/gkxs6zNkDOyT85YA0RRvRQHsUtbPQIj
7VukA4fcdE+lMwX6/9qlwsD5N3Re/hANcpKYIODWaAyqHNsg1puMX34YAWME3XlYhgsUhE6H6XLK
V+16f1HBFtdTK/FEQMvuIdQsniTzFGshJ2GuWEloR4pv53D6Nh9TAn7bpVSfPVhAwXylfy8fSxks
3sV0QeRkt0HTSNOA8KdHSg9k2O9+Jm0QaU3NS384lFeC5Lp/xNhcEWLj7Z4SSQ6DXRjXZbJ8+jGt
RQqjIyBhnQMsD3QALkdSXImsIcXL2Y6+7gYJ1hq9krLFJdoYVfiWVl7Maf076lb8ZAxX9t8q+CYL
didlkt5S21VEoEXS+lPYc+KCgvrS8+iKo6lIk830XTdrtQX23q8ehQOqPaD0OSMRNfi5Y/yeL8b0
eMwYCVetWfNdm51QgeDMP7DIaRR1jAKeP1in9B8OErUquQ4hll3uKq+oLWMU8ZrKk8tagkx8GjVa
1EdowYOHpXUg+F1x+zP7Thv+w2Crd6H7szRa+Gygdd5DkgQgYd7fqKcQV9+6W2cKoUtqLFJyLAjO
AnRZwHZCeDvDlgzoVloskvGQ1US8Kl0P6IbQoIaz0DDAdXx9UJR6kJadAK08ywwAN/KtavV4vT/i
IUSkT2llt0LKj6Lz5MPYiZeie/lH7U4CeQWOEsgtW6b8rqhELmOr22FvBypPt3DjzZmbm225SVFH
YaiQHYmCb/ioWsCkeCXyq46cuKYRqOx/kTyFTwFw8i4CYo2X9MvBWGonz+Uxn4Wyjf5rLEcQJxfl
tCbW7FaY1CjnY1ZDYUu6yN8Y60zRRrM57HWi3ox4uTeEsLj2cEBcW032dRJssByzDadofGmx9Ap5
EqAwXRfL1M0wylfurXayCVMgooiQqd1u8y0N5xt0d8P/L+J96QgKm0rYL9wdCEKN52EdpwWFcpkB
2uE9awV7OzXL26LdVwEzwy9sbVYdcmlW9zoJHqt81Hj24Y/uTIFWkMKKyN7aS5kH0CetWoWRLKWH
C9HIvAR9zWOSEzWcqkHK9LIFMIBSAAl6Eqb6DS5m9jUaNccAhg09ZCumMOt638nwyMtFvBTokWVo
+zB0ZnkPeDsfAmYCLbYOBbDca5eh6/R0BdIfteXNfnALiXh0cAHOAOnNpUZoxhzAKMnewQn9LWjS
MqbTq9zKlHAJ0SLWqzCEGFaXI9cQlIXPSVIktTR24+uIladTHaK76PBbY8lF33xZF+zYLo0H6STC
NvIMj8j8lEJJpuXeplF3Ndwo03ncMrIuYrGA3AbM6nM6HYprtQdKbkAPLwxpnprqXDnuNtDiAiO6
//FpkZs+KAlY5MvJZFNdrg1lYg7HQEOa2VADvMmnrGvZY6KyjWfqvWhyWLEIOHrnjaxUrozTi7JS
bLv7QpRD78nhAZCNWHkmXjsVRgth/fWY3/qLPxjG9jctk+0cXtfhcoLUcYhurWVhXZ+En52no3sZ
AB7e5rEzi3w2H9DXOcET1vjMWgVd21r7L6IVtvSduc/yAwQIOUXK2oCnVlQweRg838Sa9AuMbaN5
c3xfnpi02ijkxwqoePintmvMAlUsRF6Yhd52vmQEk85TeAu+NWrzBR0A+Y+ybYDhO0QAWj+1pJGz
c0QAoWjl36zdlY6Zf9wm6P60GfCEu2WvC8FVqgfZzeDlOH9RK9fhUhrOmz8sN9MqJ3eEDUDfyL4x
/x5gtvP0YKeza71jL0eWIm0Q31dLVOVe6U6k8fa+Ma1J6CkLiUV1uSGLiH2wiwJD9UgumccX15o6
6EDdtRIglbHRHHk1ckREH916+N/YmY/iciN/pbKqybz+1YcCG3H8QPKDDykwXzQXZfwNYZUBIF7l
MXN5mNrzq/rsMNxIA+niIoGBDH2yCjxc2JH67sxIghQmFhVlCiBiLZR4GUu9Ms+qOQGS1NzxpYtz
GP7vX+A08T5Eqw+N46cdBdtAw2rTPFabRM2294eZtYgx7Fx8Av9N1vM65vpXhEWWQS2sOLkz4jZS
0Sgv72AxlKwuAcg+AAQS0DBrIiGoiapNy3Ut8x91yFaznqGlCyeZonfHWIVwYs0DmWEdsKNIf9hP
AjUJaiV96Oh2V9sosyZ4mhdBipssUKurHdbQbeMmxz3XmuCLsZnNvAaDHVbTz3CIHNzG4xbgGGEc
PspKuo0guWpl/U2Gbxc/GuNMTnohAccXauQ054NNsedvvX0hn07moTq9KN63V0O+t7+6hv4r21zK
au0ZENtgAsi1XEYV8HDz+sNRKNq1YtDnWx9/ISynzElnbmUFchd2I0rlfLwdPPMgsXoXCC27TNdS
eDh/kjXZF8fnoDL2VF0PXa7vI8ZwJ9I1O5590XydZNYMtdtLtk+h4SfiriquU/BJiGROhjbcpXsL
q3PxeC1vKR9OP267SdyRz8xtL9fqh3DxDiGycsf+6ZzBqYaVFg9JrXucu5FcsD0VGB4eDcYAoIwD
lWYjLlW0j4/AxIvV98AkU0qSx1/T4Xuji6pwirpvq6PiidNauLWfCsS15P8ZF79QkKddam+KZifh
XaXS4nHx5n4U2jpmqZpciQTNGvifca2xTqlfupo3LwgELkB/JZnQneGfDivyEntBEl3KCW6h3SXz
y4LOj9XhzmYXFULSq6F8MjwvswOb3dNAqr5wtexjcdy+BJ4MJX+ahIsdi+ytqmybGW+R/Bs0LRBH
mFT8RBzuOGN52O8dh8B/cednNLTiUeDIkcLjhHFtJfLm+3WQfyMkCO3yDWe/k13bCei5B7vLIkcJ
x1bR4ZJbtdq2oz4U1gGEw9V3+FKXqHAs3+LEoTrWWQaMAex5hB3dXiIqLypH39BykV6jQGkPrTjC
mgoD5VW7CYVr7MBm2KFHVExfozw3jEgv6PquwzjIgVGkmhPixRisUnWp7BpaRojkW/VpsKYbBwQZ
3sY8s7OcAwsffc8BuFn0wKStYwOXsDktHTkPyVsLa7YshCsWFlXf2rR07FimGcNDr9W1EZaA5Wx3
8iYU2oh4i1yoUmw19lvXie5qg2xSm+off4m2ToYyfG8OQSnThH6UIDyYliM7Z9bHc9vR1E+1i2Aa
8203CzNnKPaBQuTCVVEZN+KmZqV87AyIi2wJpcWwqAGyBTAjsH8tgu9MKl/rR/L7Ey7KUnf+dqAM
u5qDi9r2oeHuMYpgSdFrG0WVDHCVa9ZVeS6yy+vLHOYsifccyaBL83NmRb9a0mWCTR85RfELVB4Q
m1oT2fTMdXcRfmcvKadHNwlsAw6TwIkt3NARmTSe90dE7oO4C3ZeLA8kc9J7rvk/HrN++FA0u7kV
bgkbgkz6BHnc7Sh1dv5tN+3H/KFMAXiiwlEsCWtTaEixNjwPyboDYp62I/thQ+Erxdeq5lKmFcC+
UsCgUZJ8Z5nMUUSLevEbfHniAwgIeIjL5ZXGrdKqHY3z6+W3/IDT71WHJvZhJ51peNhVsQWNnZJw
dl5iAiDSB1fwTSvU0KhCmG5w0Vw21Z/u5DGR+snjWZn4AbIIY7KOZw4JfKo8wKYegZA4CkHGaECY
w+RpDhaxJsywFRGZIVYwNwwjbhZplIa1wjPVWg0JfFJZZRAZfkz8DVERfdjEAyWiKVLgku08und5
nuWayWPcPZFK4lARQb244wCVUp/N5/NnyYC9wU9Z3S8Zrpx9/psP8gxVSGXmoda+lNxyRmAtCqQ4
YkVkfT3YutNLes4LxgLhShZqlh9se/VnCCKeH8vHE5hfycR5AuLHEnnvLdAqyuwN/UQ4JbahU5Fa
M7CybnckUJb6IZtpwBKSQizDnt0HM4Vhk5a4OQrQ6LeFBK2LihKvw3ezbVRzAUDeTKNvdLn2tTIp
mHZaOkfC7NLeD6mBVZbZ+T+rT5t2X77gXbU4O3Yl+YryLs5ve9WbHHmwBFxTG81TDs6Bq/B22wau
/1bUJJ+B+oWcTzWKvQ2A0iBiQ9fPPRXZL/xTHBwAUJtryabNB+24jNxcBHq3HhD4Q7GdI813XbkE
35+12DyJw4HcZUzAmHRA/q9pwT+y8X2hLtFFu0OrwPAPVW1HEHUDA9rX0qgIpZorJ5Dl6gzB3CRZ
6LPDj0x8UvPzmmu4ULP4QqD1Isa2mt3+9Od5SiiyPHgb0WOwXa/gBeX/DfkQaA/7/k82Sw122DcJ
Dxyjvcd73Bl5PIQZQn37KbJo2oxDO2U8J1bQu8NoEK35lBkAzgaSsbH2slgb3jr2+VUxnTSOUXN1
qut+/eDHV8fO/qCDGRH2G2pcZDnWnzVvHZWppYxrxK1y39WD+ghj3Q3xN5qG9egOhAW5wfvLZXVo
Cl5qgoFTRmdcs8BFvCV165CKN5mi8D9If3zjEGUhUncwEqJ8lbGSpnmyTeeUdHgxUcbxhgv3RKGn
iYVMTpRdFkDRhvfdyDK0ba0n14QG2ubDIHv83VYtZbnVw71gNY0qvpMDTJJBkoVsrXiDE1AJ1dRx
mf+ZcQt5QsDxSGOi+uMOPFtVU+Ax0ttzqBMskRk9owMnlS3I+rhHei2HxX2lW91+Q5dQQXeL1Ani
1vX/9s2abRAVgvmYdKs+9+KPmJ06Esuu9zctZQ/RnSo+Hgt/2zip8bhaVdccVcfk6DG4ZGRDxCgi
K5GsRE/elWobxy6sysi1pAV4U92GwOxLVxhEae26WFbG6MvTYzJ8acmVH5RqeCKBqhdFRiwtsCmv
qv3Z17ucCMDrhH2H5Zth4tjKMmrIqt/HPxI4VXKmEKjtW8V38LrHqP/rhRNfHF/iiIVUUGBmBfcu
SmnB2u2gLL3AWw1EdeS/oxNnyFhyGCaoaMDaR2uB6IjPr7LU07NfODvtG9OXaUPcC3/pFkRhfR1b
oBA/vIB12YOlON4Z1aOFkrxXD9+VCRRXhAWmVybSR2Ga2VO8JtNE2ZWVxnqBAhl6BLsiX+/QRunD
pzb+mdqPGmgGzue3uCqzC8e7fn7YH9eNh29B3/8luMxEzv8MZ1DnhK2URvdO3BCZHqDjtgNQuKjF
zydALn5XgPcFSZNfUYEeptVyMtn3QYPjY3F9R7vHWbRLAPFZi9rA8mkkSMj4uJPT2zUkwIrMZCvE
OYc5XHj7+/7MArMZBj7CsXquDlXCfGRWew3hj/kvd6iuBfUkrsHXQoO7VBLG3o+HqiWbBjNIGkbg
qS/BXjBJEaAsqct/QZumbIEDHRDq5MI33umFBH4TwkxxOuD3MiKnWcUVf+jED5UmwxpI9Ag8BxUF
C4/Ao4NdQlI+0hlelhBWuAh1K9pvTq8rZg1Yg/gaufHYsuPPM3L8m/86SHJDHnUqnzH9Fs7j1L+4
3fF8zGVdcJty/+vUvATcszlum9Ot4BRn4Z9NZhhnQC++GhKW4gWLibqeyJZjCEH63hlwKLAg5O5c
F91wpxeGbl2ECRSQuqZfgUiCbqHRoHZikycBfgK9iL5wMHLk7PsnkwjBnhef2BGhVUxmrNq80PAd
naD88rj7OaTO4aJSx/Lh6E7UwASEeZquQHuYMdglojdwc1WrodLE791CeqahExMmzQ25UecBao4p
7Vi3mgv8SFlhcy5UqKA2EXMHGcX7knJLZf/w4muoutWj5nMK5I55dxt/NWr6SCM0gICpYGwjqYyw
mhR1MpCP2OBT6pji2Zpv+zSDBim4TEtLSOvwfkl6f2d9EQa2d1CUyXKyqoFIcxhL70QnEaqsAdjS
Tm2BIde39NQT9VEjF6FRDpoGbcyaiVHqlxkQn7Izd7I1Wla7gSzKZfU7z32CRGPQNvxmTpfunM+/
RgQRONIe4BMyERHWymg+v3nsqOLPqBNt7OGN2PE/UGxTMoZRNhnzxKBpE2f29DM12RejdJRSSTfZ
o6iO5wlPKBxMF4yAf3m6KPYFt9qGSc+hdIDKvwgTKuRWIt+4KntJb9DG8ZP3QopWSgDcsDpkpGYR
t+0JtKe0Jqrab0BGKySqpaA/sbIw3YIJ1W7OntoLrnGXEqEuBujGNfz1qZ+GVArzlshP0kbyB86U
gDUyBG+Kh6tfWbGRXu8dM0Vw58GHUgHnHLVtm/PtI9JlN64xNiyiV1/0Vuog4pfwDSY2pGfM09ni
Q45f6jKWP/sZrZETsigCm//XFVLFYot6/lGf4A/lsE8vN6ThZhhVEdWZVWeFpcXz4MVV4Ym7UVAw
0Wmp2fzWeCN0YnnCyvM0eSpiiO8wQi7KEJX4HWM2MDSzehGO6W9hHm6iv1eYX+pdOg5BKg2clHnq
PSCd67OUCRprokAyTT7Xa72WpGVlGyUwq8F6GTa9k/tQL5gpKJoCT7174fsRKPP3T16YJT5JqRUp
6SEKPd/4FZC3F8vN5pYjpXNd+qJDM2D7w1/8930xcApVVhheyuPr3vMQVdPjqT6UVYiJJOsySzzT
iV/9FYXoj+pIkPr4vVI6LcI92RyMBjOUlkoxzzfo2Q+7STGM0tLf6YXfZibwpPXCHDFZ+RHeVYP4
NUzaq9YMSgMX3gSYEtZiObyZQsH5eiEjmH8znvjELqVMLb2nIoEyV0hLBlbb1kfZr9X5N2EW5lP1
3YH/DsHMWHEjSKSfwB8bQV6Z7+mqyBnGxB9KyJ3WfwocKWwBSGip40E+UAFA88jeQFyo24pM6jWy
j2H4aJPKRTQO+EeHxnn7bS01xDm04ybYatXo8AB9pCxJuz/QVadHUGwThxynVipsUOxuSA4rTpdC
p4xAXTqqalggDGvglFRb4dQK5fBgJ9eHQ7j5cTS3/GGLpMLesSrvQgfcRvQQ43MrqLfV7NXFwTYp
71XPBzT8rcjVzTKSAi1trEljrGYXlmJhCMIyyt7qewhMPgK6YPB52gmZizjCdDcGB1T7ZUA66wFU
u+fcActjUq6BpdAyZ+aS6BMgirkhr3YMiTSJCtycCFMoIwHeJDfRCp1fYysDk5iWV+AnVC0kaHUz
454L0+BDZ5xHttng2lF9CbX5jzbXj2JJDoNPlsGHEEfMdaRO/ZpB0ZqoNQ2bIt2Qphkz+uxXJOBe
5OfuofveBP84UsmEbesRUbYxjpF8ntD2MDNRFK4bOknUWeE3phjSwvS/wBJLNvaFBUuZSTaau8wY
YtSFH8Jwxg03EgYLvwl7diqhTIiHvcNLVe8BLx6wBaho2LAGGKeKucqwj9svHwNXS53NqKpNw2+4
hvlaiBYDVZy3omV5lC7RvD6eUEvw9JI1NqpFF6+mwIdw1di+W7Xf9i0B7VSYCuIkZxZG9gmhYlzY
3A2jouMuy/4ZBsm/LAQSLFQ3lSFl9gapqsPSwYYcqzYckhVHN7nQHMRbYVJ6CEXGppXhwQ8bJKq/
YfrUsgI5h95+mb++Wg5sATwxQ1roc0f+oFPruAi14FyTB2w66pQ2WrB6VzQGoWJ+UP4DRSBhVirC
Xpiw6bY/XA3luE06VfqQyUkLo7RoKtrq+B6zAHIMuf7BnKh5/IOMmIUqVajgSUMMzMDgyzK273gs
sYm/6ZMMap6Xng1iW/b3zBk0yQbw11pFdJ3gLJzpgXi1+qZp3HdA8BAyvlWRsP8j/s1M380I7mtw
9ckpfQONSGCiCHJGXoP0FAnl+9ZzcvOXNHcZAyCtejegvGFEfOBr25C/IO25k3JQVfZlqiiQynCn
ToiWw1ECRElS8pJgSU/LPOabVKgJ2ogRHMrV2AyIoOZI8Po+H5+ytad9oGVgwL/nnZ0hDM3f6nO8
jqRIGW9exqM2wMfCEFv0PfTJz2vzdJEaw5y+IL9yPAk6soMSuJhoTJ5dhm1EKEuXTdhmpb0tHhFn
Fwhw2UX31FXAZRTI0E+HDtqH3dUTF3e1nQ1rRaykPKb2zUTp7Ysnw6YilWuHUqRWcL1E4ynTHPM8
uMFB/y/Taq2VU1c+SGnra6BYSzUtLWdLa9I7ehavyeEcf983Quwanswr20lm/jDM4hdvCftlkajs
NYoiRFv9nN+dabeqmQ6UGLgzA+vFcu1dZjdlANGyz2lPs1LffY6Cj5QUi6E2eoKA7vWphXEp7OgJ
jIgJ0aybxJvlC2bxFqpbr609KSywqBfdPigLfnS9Lveupn99srJTa0y8dY26x45lnknrD+R3vpjm
tvltz+SpjpWdg7hkvQknHi+xcEjNSFHGCdPPKm7OTt2X3KA2IbYjbF1apdA7qyc3AhMQCkD7IWLn
QKsWWFSDw3ENed3YOkDQmPKVdjZBc87K5wFhezUbDqvYPQDVBIs75/lFYRWGl9W9uMofM8Ds6Pib
Jsnkxq+9zsVbP+gvTSxC8ieSWvOT5D6PMIfDO/CNtwqOYoExD5oHFaOIIcM2uSdblDnVYC3U8ayE
++J+MFWBrGexxfQjKrV+w7ZUM/VqBVcn4Fcl6jjtMu+UPk9bpyYChzgqUSzQo5QxOd/QKvL0uGwW
hfnI02+u3wwAJEJ4lI1EKlprWWONGd+ZXsgA9E8/rU922d0DAQomNpypcLAsN3UxldIGankrRzoU
Lo1Yj15pWtuQKzQzdLy7ZCbLwXaySURezumejZRmiR+YVh3ozuLi1GH/mq/7v+bi/I10CnwnP0LU
sBCZoIdRZapKetM+qAKMOzfJaeILydnk/fDG4A7jzUu36GhW2mngQ7j4sUyfcw4viRmLV53zyZq7
qdlhOADHumO5ZwJYctwsrvalhQLLZvQgZThuzoi0VSB3X+868g/3h680h3ZFNupdzU/Sr5MCtHMJ
ZXtTjp/7KV1SeC6UYXl6rXbx0LApkZfuzPEay5/c48VGc4SrFLyv892puajfylCWa2fcMctB9qDI
/+ddWSoIkYpLsgzBLV8tZmaw3baEx244oaIOuwDEi3P35y7PI15fxQhLcC7aePWBxHb/lz9HjJS3
YP4diohwZKz7/8aUKX9fOz0wPcKTTL1absTBdQgNLDpG92nYwK0Xw3Ju9/mQ0lgg1Zp4balk2mUN
QzLG6QnVUwuJYK3ssHRSunDcixH09SYVYbLdZ2Xbq7pQhcJbwPCAfjxkPAgS/8vXBqRQv9igoiE2
FE7Mo+FkzSRM9YuEaERt9eUvk9gmHRFZxjX+54Fab8LnGJluvtsGt6UL6NdoMedrlxgj3tS2xOLS
CK91RiSn0h62zQOtASFtiACJOw52gx2EB2JLiWtrZq5MkoiXl1GcT4K1X71gPc4GZFC5rkpVnRnA
su4m+J9AaDaSFYR6CoBaZTIwI+x0DZWUsRcQu/KmZOOPKbYZXpdhHqCRskgbszTvcnRXrxQYo6XT
3RoyGCMIiUa+cQ3G9ZUZF51tBXTDfZNo+S75Ckvn5ju7fPhrHeyGOJObZe7CDQJV0nLC2nhte/WG
mE25JDvh+qtCYYoYFAL0A2hlBG+BJqeex6alpBRQf20SvqSpabmoi6X+25k4oFjpR8p55hBpkuaA
FxxL+Hkn7+xpE8HMWoRq1c5dtZJUqRLlKnW3RR7vI+doImy3rp8I5LjFeDCzlUZNAybIjubDU6qr
IGw6m0S7EdaAHexAf5oZ6EsUX4QvWO0vtclMCAAOCfpa1XVWdqzhpwi+2yAfNYPZcvMU1hCkcUw3
qao16loMpeuc+lOygFkR233VlsnaOp8pcDH+xJyR78Yua5gESXdoBjCj0NTeItog2LGEZWyWaGE/
5NCICWA/6UiCCg0sw7vJIPi9pmV+2vGHG970U0HIZ3w2atZUXRc9vyczld8rFW7jTf8WZiZxbcGz
MVtyj9NFhwUD2jjPhKY4XhhSzIhc7Ec3C8UJ5quS5Oo7lIjJXqF+zcjTBk4xRzgt3t3qI/FX4f68
cFj0ufd7gGxH0MM6XXGMvRMHlywtx2IBj+ixKCLL/reWEX31luwTSuU23wqx2EhA1rMNpjMmOjIV
lvIwMJvVAjHKHLV+rhfxlWwgql412Z1d6fRDsYL8zeNsNDU3Ll7dgbiMVNllmfSmsLo7Hi42fa2B
Ie9ANhO1wEGHzSU3Up06j1zeJys0BQxqOtsWY6T5C4S0VD8qJgYMx2Efcxs1F4sM27H1rjYCqBGm
1P9Tt4rxCVJRINORycC5ibNwWKtbEJptooEtPg18MBmmtF+/7FaLl3p+qPBDWUSkqh1yw2knChfi
g2P2Z6MxUgC/YPr3pKtaOGoHZXHe1L/RchBSS0Wu8tkJ4ROH3gUCTH/xjjEfMavEzZnPlc/CCdUC
eycdYlHxxIffVocSJhBOOSbttOG6cAikplFx/Sf49Yf13VOzA5YAh1chTuDWGuxB54AC7bm19OMQ
jo775OolZ1BQjdzHt1LPdkLQhReZUEmK8SQ9ZH4fSOi4KULcNMIWGvH3rv7tqAQ1vAQNvo6/ZILL
U+hdeWeHVMA7gQkb4MsP7/1gfTTHBR35s7L72oG0TjHBwBgA3r0J6VLoveT/NBh4KEnY45oe85pU
RMk8A49i2Eezc1qc5gNh0FI8NnA7nJ7b7dBAj5WL4dFgLyDmkvD6wMqBM+KywyDiOQB2L0wGs/4y
vLAsNL6FfykQbL77vzY2zJYoDlPL8QYbvsMaAA8Od5M2OM2xc/xs+8EMULeXaZkXz2HY53USpP7+
Yx0uDoex++osW+5oTqPy3irMBJKQlJwkwcnti/6XdK62rBcX8DDHRzXag8ZCF7I6erKEcKX/K8Ov
SLXBfj0Dyss01umBX3L51PCRavBiIGI5oAIX8yAugZhlkpTvBw1kUinazYCkxw8OYHZQAFq5+p9M
ceTUUzEVs6e3eDVOkEZeJYQyAJtK0DMOn999+goWR9MXP7s2WxBz1Vx+m06piC1iKY6JrKER5Vsf
qA4F4Q3NsaM+49Z7k1Zxd5tCcjL+xY91X9ZksnO+WZwiSjipam7/EG021nGLGbzrEFoZzfqflEdz
/tuTdak32tuuo0FYPRz7DMKWQg758yHlBcEp/Noyq1tVhNa2tRdWrRPm4wqa74mpkD6Ak6GCRfvs
NLs5g4AnOYDgouaGU0lTfCIgmggukQVcSLfqkK/WWBlXUVRLCdv3c+GombqkRNYduZf51NOXNOvp
cW/1GgFm7eFph3QtCFd1FdddLMC5yaQRzS/bnJDemNUk/J9FkHcX4O2jlg3sohDxsTpQf5+FYwx1
VBTRye0emzFScXbXViF/C91C2MnKv+kzGJKNpart0MecoJnqCdFOX/3xpp1B/lgoPd7p1bR2eZlf
UbOHsoq0xnqIrHKmqid0pbM/W4RDPY63vWSgmySMnale4DPXdoMNAViwdJ9s64K7gTyUxtUeBStW
AaCbCK7zz9SelobLoeBewt+LnWqTEBgdeJIpXeFhyE7t6IElVFAtoTXWS1m8JIE3y+nobKOZDJu2
VT4foFufS6+k24j15DnqNMBJGudCGhH4XkfOVmiXy5KsdR1mNhqIADv/DzZEnM/kNvb508xhrwgU
ztjfEB12z5zQfONyOUWNPeAgLsEH9u5UX3MumLGLwreSWwtC776sgrVjsG2lPdc6TiMES8BepRgZ
RnWZd9stNC/g5csrzyGiWCWUclVXEc3J8dfVmX3bUaSDVizd+0LcTTTKd/5AM7nNjehY1d67GR5K
cWde8ydf7CF0mI3cOJWOVGHZuYvq72Z8dxi03pirvejUsQt4DTTb4ScJANKJCzbXzmpM8LcuFy4M
+OhMayIs6IHdCFKm+Ypg2l0Wqpjmw5hFvpoFyPLci3ujr+LTZXVKr9ijohPtSMVHhwum8axiVruQ
5x+gyS6oslwa6wWAxAgNYKET69OS+U2UTLXSPu2AO8g3iLFO6ALkupmbWs1rYFzrdn84Xk255Q9I
C33JPiPcDOVK69tGLCsbzYu41veV2K6yz2CNGzoIHnDv3B2FJqyGyU7hUuyQTimxXq6xDgG7I+hN
24tTYbra8ImqNcQZA9XSLE5zBipHp5iovRoZva0OpYx1bRlin7Lm0gxtL+Ht4u90Yskz6h0R0cPe
gyzXgD3kqyh7NXwe/8YYCMSSiwfVqQZMBrEdu6rn/m81fIFDcG3w6cgTZyxdD37QNw+1AF6l48I8
FLqUbWEsYb8mZQcrp4KRdrXefjtSDHMvrMbvbr22EXpOEFbnKqwcaWs0uBMD85alnNkgHSK+kaNb
E9Zh1zmeQojaTJDq7H+5kYbs/P+o18QgOZN1OMFCr46kZPRKk3L2NX0ketA+4Bcy0DOud9nsnPhA
NfpDAE+3pZqgs4bia3ybLnVbujdzaATW2DWnQrOx2oBik/+VVk+aXtb9EuKvYu97BFRc086Ww2kd
tC1nxPlyb34sSVTqqK/pkWC/xPrMk6v/iFqoq9upTpRJYGl/PZLHqL02RDmKGkCMnAPE1ejOxPCS
YoeBVF8UZd+By+uvPZSqhDV4YcbRfEhO1DhJS9hrFR1QIX9ilZuEqya0k6GiaJ5YNwEoc44ioSb3
pia0gXq3MeychIjP+AVUEVpjmDnnzOmVjR4+4X7uuMeJdmti8mzjCep0Oy13Tme28F4mFUNseW2t
H7tmYAYRdtbC+8eRiQBLxvOGJYJzT3O512WPxfb5GjNfSndF+encH2b3RA+CD6mKJUMo3o/iO1O4
8PLG5iFyo4RsBEgHlRE6HBUxzJM82pzEaEiRDS076LRWLZ7CT8peroF3jjUyZCisFPdlJwDkMq5y
s0TzXJjKmodZpWq4tRhf+Ypj449z5kr/49JbeFv0Y2185TO2KYxIeJn/fJan4WhBccaSqf1NFaSR
RaB9WBQT43YBuRhRgR3UIcIUG7sapDb4wlAKL5BYbur46PxsmlyQ9a8BzHBSXTfWCB8PxOnhAwF1
e+Cztm0LnvfwJ0+oJa+36f6XheKAQNLsTytgzoHX5iv/hG12j0WvO+9dbR4GiZGDe10r6HjsSLwr
AIgtCH1usK9Uw2wVZIoXvgD8X7WVI4v7rmCIfpMavlT8dyBG/uddqJYZahPH6pRz5XeXvNGtBiyn
VZGmiV1v+PoDRtasDnDAXzTESoNwV5kM9SmvqJwkux1LzCxuHGKwh5257I4KJjoztHWvzYyelG7L
8Tj3So7AAjvzrTeUlr69lz7cIAbH96vOLemtvlPGRrqqS/NlPw3d5IL1eh9sX237i9tBwP+NKfe5
5DytkEM6WBVhzs/aq5lSBwMv+/2xmegDM38yxznnoBtkWhRbKBL8oWjZYurbOb0Xq4vxm17FXiuh
s6yiDTqnZlFHAFc1Pw+MPVwgT2wJCJ5qo95AEG8Pbi8/emOASjvq7Q31HLST4RUePn9IPm8WE9L+
7bO7QBtG90Fb5msqLOgLr4eO+t/f2zfr4TigtpmfTfahVFxy3uSwfowxmBq0w/cg3F44/jc5HycH
IxcznhmaKzaRi+1SCeDnGqfhg33e5J/zmAUM9kbjNs1TAfgzAK4T/OzjFO5+JeeYJJqaIyqN9n91
qXwaIpv99YuyxnZBtMC8BYkYiV+mTUpSTlsl2zwrH4sfkNVWKFpBlc4YjJzAn4u+/je8/uVmZSd8
sRQCEpEyImwDrOqxS6ysTFlzp3ic2nBRRdqZ9GwXNJPsW6qcy93/VihotZOYhlHVqqe0eMjso0s2
mVvyMR30QjgGBiF8aZUB1etFxtvnwNOjH6hydEsy7gcreChDkoJjvKOARVGwQ0cVbicsRTHqZoO4
3Ca5OWmKtEMvBvusF2Z+TbpfF1XbRwbK8Ti8YwVqFxtU1hZVQ9vwBuSGfdZ3qkvOBD/gdjEa3Puj
+FW1ygJLiI2FUWoYnu/pwyIvTNIYRvRE6N2Awa1sOZWj3wL/HzlDuUnhMbbloDoLMTJyBL1Okvmz
iD2jKRZl9/KaKZX+55kPuOOYbsnESZaOhFpAL8dSvR3oa8SaxMc8JFakLq6fX6B0EdW6nlv54QCx
fR/i+ZkSaFHFpvmLwwYQpxuU4GyugKEZ8kNNJGkI+StUtyhTQpBSVvPOiL36ldaAWOA1v+tVouqN
CGDszak1Gp5PgrcXQZTJzhW+6xoxiTu9wIuHjjFdJLbT/PcnEWdVPP6NVxxmykFkkixtGohd4h3y
svo29N6jz2xxEEV+fTXVfWbvETAXQkxzs4CGvaZi3Bc2S3oDbJ3r6ndxYe+cAF6lDaII8VW5Xuq5
yqLdSEfcVJ61dcXLP+chQfnNhP7sya/1ocfVQEfa08Mv/gMQCIy7+vd8daLFLOsiEyXFLFADl8tF
ZZACW9PFJXqLP4kPocZ/CZprsSYJWIMPzD1HuJaf66id+gAGmbDOCMEuhkQMAJEXP4AfUF/WXqdx
OfP9V7MWk1YAfpQo27/8NHve8jZttkpkIpLy1Gpb9HmyRTqZIOTriEah+snkNzUqeUwFmwoWEVsY
SvdpJOg4JCpSJ4F9y3nenWz8BxeGM0OlS0P1eol3diVgZBNZr38XlZoZOE7J8E1wz8BfOC6phWy1
2TJucD7XkAWIvLFtUMa16vhSDtPFjhpMJowhSOUHPggRDLnrGn2OYCX1WkBl8IsPfq7kvDZPtGr1
6VOuaxv2IntYCucxGnBfgUYN/3FoQDVjw45Jrovsu2K2S3AwyatQ4zsPBSkwnzH14WUriilrvG3A
uhNZs9BNX02kAvy42pMrhu0A4Z/WUl1MAZ5HTpGMMrbGHxpAKx6jdmDKc9HvNGXBn6OVlbeTrqhi
9FdkOgpmrhqY9gqHbPw07WWWJN2InFPiAxe9xrBk0pQu9yVHvIWYKltgWZME8PWV9WIebfW36s9W
YLyflsqU9sp+waj2dE6S8TQgOAQs7Rpz1GHVEowQK4K/PI0ktbtW/EucOj5Tyy1JBUyMhQ/tjb/3
29oz/Gy4rb7n7LWnj0I8Umspsbn8CKuKW9AZLnQmIwOTYkySK4HMgoKu3qCWJA7Qwpsi7GO0G+Aa
WrSLUhHbCN8Fex09xYkHgCqWsXVIyDiYGzg5XGjnozqKNf2HqchKMC66UTCQQvPwX89sfSuWKYu2
5bgAbb1wuOaxgXgRMKOuP70Gpss33eaVh0FYBlszQ4NYOi/tW403yY+Zfg/D8M8K8tZWZfdjgZUp
tv7/CMy15brSdWLTmhSwEpKLrXGcygepOmd9xEmnv6WPcuxg3xpT6r1m/4awIM2vS89IwGvlk16d
REoPH4wUkKlrshNhZs7vsTiVMs4VVwn4+BneQRHfPLIFED5D3brVZq+rS51RukOOKsoq6QJ+wrpc
fJf9XUSe/oZcwJCZKrz3c9TA/7brnFQn3D367qItQauhDtA37hkBrQ/FRlTmzkXripexB/cAJ18k
sXowt8WtgiRlhUR5YYwwiYAz6TKGWhmFdyqtSEOWYJ5UhOaWk6yB4ZNJRRpFp2AMFeqxozV3oW5O
SdJ3JViJ7csEESyTxucL2ISE5OEYn4JltqNH3miHWyF91hczhCbIeFGkOINKofwTq+flU7g8FE7s
xByZ8cFR4/f8MKuTabiQ9uhpGFu1kb4SYuzBAV0E4JG6h1w0Rj32nOIMCUaH49ZMx5vwK3th9FEk
Bvdbr6sUZi/EqFGHzeDVLdSdZ933HkztcWUelTnmPgbBuRC7qTan7e6IL9QUOcL0zkfgR2SihnA8
PMqwFcINA8JollGWA63PvqgD4ZTmp6ZxwiAH3t/os/MwClE1yrH5/vEWqCAsrMvNjxbrejP3MDGp
TSROAjMBNLSWPnAcs/+PXYkbEdHGzZDWIVwzAIfAGYK0ONNLJerrS/C0d50938nJLnGRBRahNa6+
JgaNht/UpVXPxy/J8tXvDS+LTON/ZQ69QWgEatjRYFpCaF+dvkOdv1xTH09wiSq42n1u0EtcO67r
/33rpF2LCTALITYZTWPNoua0RLeismAHBUStheYh11iXyN1GNRNhy2NjOxg+9wFMEZc7fzAYkAnm
RaUOeGD6I0SjEwdN82jsJ4GXyQU/+YXTSPwMg2z1BsURFOjgvmFlrcyw85iG6MSH7Le994tbjuR0
xaV0iTzkMTadfYwIzW+LnHgSj7MQHJHtYoAyIiZ70v+AdDP2DViN3rvNsZpsOzV4ZdrWafa5el2b
1GRd8XGzWhkqbz3LD8Aw2bFz6BcWc384A0L+BXnH1fXV1dA5r9RFFnMnVFFCx24ieS9B5uXHNwSg
Mukp5+9Kns+PbWiezHUqgu5dLDmt2Lst4cK3dZHS26RjemPTxMWbEetsle0fD5qzSlQ+dY7JR74P
ZhG+lyi0i6C2ldzg5mZVy3dYiwmP6E3vJaDLBJ0OzSRVav41EOPW7nF1jS8Ar9REcCpEmRpgvmhO
rfVRMXG4plWaCQm+QF3HXQMHYypsZBst3SCxWP1/ZQuVyAf/mGFXDVWaCWS2qEwGrcSIjeZgDAJ2
9QcJUCzwxcPaKMtD8DgXFvfmKQc0do0pyzOFSL0lTOiW38L6kngktUMdfD9P52kyddaL7G29TPCQ
pLYqFno/gh7sdnhYObeZu446JU2+zPJ9dvFZryZKYON7VFvoEOL1rE9O5i8WYwUWPg9gmSGxblHk
N6FE3oizeM/WtnC05DE+yIa15zrWKv5OaJMa0gFjyUT+6wovCVWL9guj//zQIfKx4bOyvR0AUuns
oMFgCap2Z+xADDYTKbAoaQ8UIOCHuKmGGVFxgSpM6OReQH4zjFMvTgfqYJfl4pdomvBHEZclU8nR
vlejOk6M5TzNY2RwbiIZYav4le0gXEkQy3Y34HkJjsmtA7FCe3F9xJTuwUybeLjnWZx/5UV9jTMV
xlpeb5gOXXPZzJgtH0trCMfdE0ZmEI0c0vt2xJxONwFHuLG9NNFD+6DAZTbpN1UUmB+IBpQwm4MA
ybBEbhgez6g3DxDYc1A5LQIEsIevSurnwDrw1sbURkdUjXFt1XzznvDlf3nTPD3lj06OMdQ5k0ZE
LfBY8VnswBHfkViWY2Qad3f/Zcb8VeqLwdLheWLaXKwylAuACgMBEpufSodrmCg7/7+PWrUi4GOS
bVayas3zfWHTyD8AxRQlAsmu28E6Rrxnc9s6DO4L1rpKiU97k8PBdDNNC1F9VJI8SeQE0VLmqFOf
0DO7sqQU6cAO9y27ipUcN8T+IAjNpgUHC/5McDI67E3EQXCTv3VFgDqfyYSaQaUtyONJCJ1biVgG
H2UxjzeSzWWuSFM1AFxVknPIE5+tmH0AxBweNtZTOQgSMkkThIx7OLFuFrJJmoRSGT1EJBuPuIBu
NCsq1b0dqClk7M6I2J0oqV23BYcInfaFEUve72QalQWjx+ZxTb09y8HRhqGqcMiWhJBJWmPM5NAm
iX0DP1jXU4Z/LKJ+3MVIycAXPd1N4AHzSJj0K6wo6QK1BwALDNK3cP7NL6Fo1owMcX1tIu6jwz9O
goNphbOc6X6JoLUGLQByMYV3bey+5VfzoMt5ppYJH+wZhImrSEeO/gcVocIzZRXckh4oqGMcy1Lv
hm+CFh6tQRhAg//IomWzEEljtAyJhChOjjccq/hldKEiJsX3Hp5cgOBPZI0vjouVkXGWJT5HJjIs
e4Yl0WOXRb7WLBVr71gkPQgPvjc+dGukTsdM82EJybARF8+UUqFmmggOj1rNRWEpPYsAsY08Zl/S
ZNrYGf4dYyINialw4q0hP1ls83RWFZ45x/j90Qe4V8omEAnbH3sdq6BrfX4SZMYr1wY/cmOO9jhE
xDrIwIIi2DYPGk9PhW4CeIhKtzLg90NNQnm0ickhVIef8V238ksXRfKEPC+Tux7lMczweBO0fNeT
hgvfVg9tzLh5H9M3J5+z/gQes2UE9v/IX5pj4YNvcqWDknYPwwQYOGwsm/U5Qk8o5SJHocVBVWZx
r4e7mi6GsKtjd91JQmsPf0Tavd7efb6e3kPV4AEAg96EfPmzBdNF1UIkA5SPREBfPRrkohtbu8MT
CDnUd/DlheCvbrNdDS0zP4u4wcc5RzLUoJAkoQFCQkSx5q6g8T1UEadpI7XjBmsRJOWBdoLBohkb
wI/rRG+RwHxqEBCrZexdra/tUrA7Q3vnnuPx++Wo1N67nKhdwbLCSLLN+PiLRNCAbYadETmK5kV9
6FVR4UsvlBRjAwZcdx3vM9yaK7nTD9T15lNp7XXMbvU9J9zjDtfO4PFzzjyAVWH3dEis9hJZy8o6
l/NN7PUIb6jYjkFniVXLNgIjW8NOQ/KOSzACfDucc6Sn/uWPv9uJagLrE8tlmfpo1VMM0C+79Vgs
/3o+TPtvq5hEpcFKbUZh8lA7hgGs5e5K/rIM8pmRA/GhcJia1pUxpw+MtSCezIzcZSfQBqRk8uyY
LtwVJneSRBK6YNaiEEYLXVunU56TfOgcRrNr7J+le4qkwRLOrlI0nHi89VEOAYuZ0TPoaH3U1bor
XuTgBxxIh3uF+4hiE9msHXc1wdOrWh2TI2639KqOZL1Ti0JnYTUac0+N7fIHmp0LFtk4SGG7uCAG
rdIs4fN6tooXS1wo6L1hASG9U7OfwFx4WxilrKVF+lpPLfMBporhZlyS9iT94gFATfjakKkeN/n5
KtS9A/+gAhO+aGBrEjmZOSumZxpxYnYTbn8SgdkW/tzA3WIXwVqDaQGolaTs5RSbFcQB+S3c1v9M
6vNIQHBucZaN1E94bHUEEGTSqo3sLZ9Ruza6Roj9kssNEqVCgbuVrt+YquBxiSZkFhl5KD4nyu7V
ESJiYCpjgKChVnnCzLdnhlbv03Db1E/n0u05zhMPBC+z5DPB8vtlBeYpEXZ0tzstIaqcUdgktTyK
gGZ5WJDZgiFb5jr8NL3aJ8FtXNXaV/jg6l7sEO4r48C6fU+mK6w1OXsWp4irirxoRix418ZYghtO
OfU4oxPG+yiCDKOXooU6yzSSz76j9bVuovPTW4pvEyRltGQQ84P9VoVexhqYEzmoSDG4MO4DJwRw
q0TmNjVamHQ12xJ0qerH6QizbBGTKgOuLRvagY+SZhA/vIBFiFmBNapfu3hOgb7/t82BWUxl26Xn
+KBnHb1/QDdWk0ZKxXAG571pkWawYYutUJCJw4xoWedCZh1cNNgoS20eJREbhWJkB31hqRN3u2K6
O4prb36Bh7bdsROsp35LbeHahqVAPQJdHU50UF25toLLXVHdwRP2BHAeaCNmAC8YA2VpmnEnMwPb
h+ndq2A8xnVVnvZpM4eYy2o6e3jmvi5crnT1Oi1mxUap91dn/l4LiX9jmWBn59pzoUywpq9A/bvt
1pcyLCIDh+LAtKYllzetGHt7QiUAxFXPe1uloi14RGpg8y0fLLrfRSLB7E8zo2uRhjwINsvhc4zw
BFMAIaMSOD/Qn5JANG9S1qvQHhQiiFSGOHkAlEzFFpQrwvkK04Lluz5sWUdoMwpHuDJHgl3Xdh7y
Bj9Wm57eXoef1WK8X8iqp9WeB4qKCYsdzY5UFrY4nbQb40AIGLha5nWxWOPkU52e9TauvmeEce1i
3JFXNUUORMdpWZAKIIWabmxMx0+DovsxkywJUT1Z49/Adgq59RRP+Dd5G5JSxJS5fI2PQME9clZM
u3hZVCV/deqPFRkAdyX4J9Rx0AOXksljI8hdzpC6sdLoS4Z3sn6Irus1zUTiCL3sr1wPNEwWL26N
vh90+yG0XR7D6Y+R45uTPXLRuIm+GpVRaCW9FGt3/i5cX8OCq3J22PLPbH1oaPwplHqMRDl7RGlL
4L1A2Hn1ud4Rv2cZ9GwrtFT8/3MZ3r25WvC0NJmT6zI8HlKMr+dC7dMEo/HSFKFXhguH8MsGL6sh
aXzCaytWHAzHnxXCrpcVsh2oq5swHSauOrCoDOwgINQFYyMGqno9gjCNRliarOB2fe+k4XVwDbUj
ZxbwrO/VFCDBS9DxD6Emovtyf0ZBW+dSSNU851wAtrmaty0UURR/HSuhPNFJlGXS8VjJdr1KPQJX
myEpTK0N4lnuqrQgx40U+M7D/quYSDB0SO4DbK2yfQMhKbyv1oBSODjsHvD6Zms5aOmLC1149bA7
mkVPenODZBkkE4WXHYtegQt1YXO4RaXR4a/YDwEENKwnP5TF6OxzmcMQxoxeNkbMqpNG3mTp99+p
nmcNE+oZMx9po5sdhRlh6LIJtBCe34jBKdSHy5zKV4GxDAzmZPALnxmNXQzBKxXBvh/6fEqd5w6S
IwH6XwZUL4EBSbFdOVe+TPaGfKWxUHIOSEnZ/Z9TiCDuhNl0+tiCu9q51+jJFISzv54wf+WuJ3BX
zwG7/r/IOoLrvefOAgD3iZAiIBnHQc6cifW3bkorBKgQ8ZCIOL6bQf3aikbSqRxUFk4+LN5G1Xsg
xEaHIsh+0LjjAqoUV2tM7fzj/ZkF8CnQyyMFKPWiFpE/9dd5m4CvStDpLp26xOUfdSkxvSor0nHk
vfND5J19UigAqDM/ubD2ChJcu8YwODxw/FQt23PStWXJkVzUN+p5tfmVNOU2LztAt4xmZeUGzeaJ
LB96Z5+TiO6LxXAwKNMhSyiqbNB8y3ol1Q+RkvxaxXOhpBkSxkUFUcXsZOEo1MylGt0QAwuFIIi5
cxOlrfwADajCaXXh3WhfhqjIk3h8fAr7aWSygXc6OlU1+XzC+h6W+uc10a+EPEXa9edoJ57RiU+G
AfH8QIqS5o2HGmqPjxMxcR318Tsb4eHBUB0ZZaihJwfncvoKXnsYW+If6I7BVituu/YxqJ3Ubco1
3KWMBnr83ggoAjj2+RhrsD4e/2S0NUjoGIVlEi7ZnFmSiUGiHIHi7TGd2K4qcmbOzDUrOSG6q96N
lN9pz/sJig/HIrmnWQN6XHYBfoZGCoRCI+2EULTGRU2cfZD21l0jgpZEG60351OgCF5rgebJhKIJ
6wAAxNG9F1zwgVH8YVq9yvkrRgf5vHQ1BWT4+aReYZgbb9Um/9MvjV6qIAZp1fyhDMydCykCjHPn
u+0QgRnMl1NxL0/cwJ6GbVkFhU0DCpuPGyNphQj/BvLd1+bsr3wG1+nXzMv+MbMaB9oW4+CrqV6e
Ne9g/HrBcOnlhDElIDlJ+OFofOdZuDY2zvYIvtxkUL2hCW1JtaKNAjRIn1IRQIsy3H4JiaTVb9mJ
K6cSc/AICw7+VIEaTeDJiOymeIvNZES7HaCntY9D+deWAQWJyGLCEuE0RWwgl3QRcCnTostjxrMa
5R5BF8rS3gG1W7t+qFCjmeMFyPhr/99HiTwYn1S0MOzwFfQf8vHIdVHvhmvDP+n1NaMi2xSjFJjs
u2Er64iWW4l1Zfy+2z2GeHR916dAh//leC0mJb3OmBEivamvZClW0mXbpTOZkqGFeIMu2Js/tUse
8DcVLFzO91cYxFaWUau6eDFcWCHEbROMyh7JrGuAQDkqcE/DWM7MTbD+1Og38a0Lqx29E1+e3XXx
bFdRb2se26YA/tgvOoscwzaWXFniubdtnpBSaff+gpjHmXdNJKw4lgI5PAWNBJ4TOS6bEBhIUivD
/IOslK7J/FOkg4rQGOzDVDvYNp4iWTMTN4tGpFcuSX6TQXHp7QpDetLaNzj+MsiKasFFwtG056TQ
/zQpqXFgPH08kj5rf4+ICGPglpGLDHWHBYd5HZ7a14+FW1qNIIUn53dW2dySsXwPqBObdHFFEayp
P49DWgRWXuJhjLkm48BT0395XL4wS4s0L/Wgd7wtsiJ1ZH1miTW1LzmVNYm7jt69vOEmxn0J92bd
XaFvmqe47HqYQYx7QvsFra4O0LYJJh2n0m44fwGagcLikqvQ7/HZpfJt4dyHtvkEVsnulKrf54ir
zDmx/H3HLgZa9sRBbCmGnGHx7m4BjVba0egk7HsiW42FctnKbzN9e8IyAQXp4SrTkrcfgD2nWTJY
QOdbSodvnzaE3FemlJI47cDouLso+xsdB3z+mB6OSu+aduOzkIyouXLmBCtzBCesc/BQ6egIp8AI
1HDvhspcuDEb5uy60iDPx7a6bwXyEOUh4ebae5sebWgrXyR+myQD4wT34gdvvlP0Nltxp1w3MO0f
i1crl+VEXEx/eosAYtKtAs8WgzODgv2FqTsRHLN7PiLoxUmzdE1ZK581wt+BpPfN8GQbHVRDVI2+
GrJE0EDnhgpFRH66OgY7PtnAnWGPvVXPe2B/flHclO01L68d2o0mW204TclGXm7Dpgy0XYZ7eV3H
9HwvWfzdvAPWF/2Qr4RPOboIeXu7FWWK52N45rFjN3+ijtOx754o7dtYWyaai+GLmdHTx7+ESJyJ
8Bl9kBZmljjqImog574Cs/JtQzJSAMP2mYJpXLmqka6JVAA13PL584ywH58Cut7GS8dFZ/8V3VIh
RziDLyC/cSHmUr4G1yCFTg5wmv8YcTG77VHwAlQt+HhkkNTmNlv7/CPYATEh0qkUcOzMZUyd44ou
FSU39Ynx8MFz1hBPSrU3WS7QXvxkexKnUDNbgyITTQYtOwVEjSMXmVb7S1GRApxCxrbVJ2mvrIay
TU3iuRwl2mWFjJleWuXEImB8TI68SHomm4oreplCjGh+0i335paFcFNBWrxSqcglwUxeqMCDX6++
VRiG9kDBu2pD1eUY7riE/orWgrqdwd0YEGHR5GuPqakbmP24eBqnyf7KxOziF9WqD7P0/kzkLFK0
RY5hQKOqqGi74p3Bo6tUrYWVNOyXTtfWdYpc4nR+9rBTTf7LnPSyVRBrdwXJwzVtGXS7uknXfRgK
qlQRMPKycxX9NBw0taQQla56KijBzwX/A19MbKo1gvYUBk4ex6hmz9PyhmVqIShHvtR4dshD/dhl
PxrbUpt+TOct9njWtC88DOznWpLEglzqBOuxcT8Z0LIVYC8Y/Jwz90hBnt+IbmP7YaP6Y4wx8m+H
byLQocinN2ct2UV9aZ37N/upxbytn3XNhzwDRWWwK079Sk2Gj0tdEQJtHGGQr6HSebOMXRfsLQGB
mHKR03oRmHewa8egkS3t1hMecNC0OjEU9oK8BxCxDp4Ej7aGwwdmKbtHfo2v5AlJabQSTPrxM7yM
1EfxespOmqLrePx2tF2ZOEVFsQlmjgZDePSbUkNaOLoZfNQBN0a+tvn9q0LJ/UvWXUm46tNpeylX
RMf6CGdpZ2GCOFbDIYTt0U5nAY2F5cqwei+3NnYxpcJZ2U4lfS3nPR2DFDkVnr2fXUo8rivSPP71
KyLyO1Fk4SuTcXJu/Cu6GaAYpPt9UA4zhFeWNBGceZBPLP7JMMITZFyI0p76BDB3DTCA8+480gz8
EubAJrGOVGbOby9whT8mX3U6KDTVW6Wy/5TX2PQhANuANMdKB+LIIRhl5z1hEzjYFKjuJDFJcty5
OUc6yJGFIdcy2u/EhuWD/7/zu4aqUMlH8RZHull3yggP1xnXJ6iefAJ0AyIU5RR2NSqnNId+tRdP
MN8r+z3noJUAt+wd2uMPGzgNSx1BBoVAtnDRmdwp74XSygmRD/eiKOu/mG5OQn8oqvhVTtOGGenU
yitbiPB4J2U+NHPm4HXG19dTGwDpsfR3HE6m7yVzNeoprLmU8/Nm5CzbBAupzBjmY/s2++7uyws+
g7nTSu4JarzfjNFMITKIIVUmOroYuKvzULxN6D3SHzlQtDAKAW/sdlgtlGEGhj7dkqA0j8kWuN9e
Q/yVnw5xBEsSsVn7ggvD8yzLHbBoHFNbZoOeIir3Zv6dYAL+c0Tc1UkGjxACt+osEM0PYrZDeWUz
J/9Fnfen9+AMEt3tXHJiieYg27PmAGYPr94PL/4Fq8Oh/wK47jpqQkNpckT4cuvwFtUO6Ea6XSb8
7+wa90OGRcC0o9S3SBypnf2aQBdziRi5xQy5+YUlMhNozsbI3Lr3HeQsdfTff3XubJsYVTg2sOPw
xGtlTT+MwEhtpTa/22QmWEwhyJlihtwrp7NQsFNxd3bmc2zgTp7vYr+Dhuep0W8uHL74GlozuLkA
cbpuLq0yeN/eLFdxW75PHTlxjucOl2IdjoqvwFYG9tnaKy3zeMMpaaeEcA3bZ0Jmi+GM+boxZRch
pAJ5roV3OzpNZBv/BmTKKzTa/lad51WuIR8EyJyU46iRpNgbiXK0BHVdGozev0M/ZOlRBnWpyRtL
tz2uiujpCOAuk4VE3wpaDEkPLSioihN2a7Wih2AzDxKQTFGlJrRRM0Ol7C5HzqxJDQtKkHtz7hGo
RSbyxojSeyFMItgEHQn80UdXSfDrmLjIXQQOmAFuvlDsdE5z5DrUngiKEg/E9FM6vRNrB0UnVw4c
wbE4SpbKbppQ5zhnbjoV9vb7g1EqQMo7RASRrc/rxijeh0v8Wj6F43NuL+1VF0bIwsIIV6hbBNSA
z4dprLRjcJMFDO9Ly3CQagpxlnp4h9Ocs0XZ/cMGnmYVGViaLVccDiYYqWlJID7dKjPjCewYfRnD
XaozcxCw5MN7UMec+GwWYPNWxX9y6bdrsfWRw+vKIimLib1tRw5iDAODC0dHby+clZr8N9fLdKAg
m4VGk3oMNgks1aZ5mexmMoKxkaiVP32IalOxU9AsPOsFsWDCcy3AVvkOGgBooIj2fHyQ2hNjYCtU
d19OzHI4kje18Jy+nbPCH+TsNtyoJ3cGyxzJAlIuD3QPssVfUpY/k7oOFxf2zI7BTtkWnUpxBXa2
5Eo3DzIH47IS5d1RApXir1D04qRXQI5WhtFCjCT0GSQCwt0MibgBFYmm9ymckQ9zA7Sn+auAJ0y+
P6SrZbvusl98FxXJm+Ck2jLHdaq8TLaRqV9IjQM+vaNJBw997926hcWW5yQ/8QGsfnGZVqADeOoS
WMNrSWPNIu6r0PaQboQMrWe6YuyNLgftMy8c3iPpn9KHQWFHNNWMchmuUZn7zC3Va6659dQU2kNw
T+2sdI2Pf7RUqTgcMNyjtg9hMQTkpZFYy5SzSsrr+dKOGfAK2BGZcOdG8ybFuC7TrssOxJ1DCd/h
X8TbLIisG94UU5HlrP/f6G+DKQDFgZaZXaoZm+zalWG4BXAhtNhW8yZZQZ8fsjY5lrrYI8YqZSQ8
nqg6sEx+beR+zrrIlHuVeS+qN+PbVsXsAo43p8m+Ftmff9sMMKT6/6wrXuCIF2eaHmd1QEfJO3zx
qn97ImX2Yly+jqE0dDNHKOBNq08zIsLfGRAXsVUppXJhGrtQnzDJ/dX6e9py3+1KOT2ZA2VldlJx
FdIvvf1p6aAIz5K/5yniYCerQjun6jEAd9YTyEJWTXbAjXQcd7oXqp/2gdsx7pA5NRdqKgKUOHZ0
A56zcXNceW8Hb1X2hzZGgm4BiJJVly0/Krz8nZptSg27fcSEUSrHDv9IVC9cWh1FOTIvI9pWvaMo
sm2lFXWfJ/6+jXF3ztPoCbCMW/pfxMSdTkLH3X030ApOIW6I5e9gru7dF8o5rQ8YG6DabgHb8P/f
H21UViBAlRlS45zYcO7I0fMdzcYF3TlWtl77bDH927zzw4b+OuRlFR/qOy6qVaRiew9417XRxFfM
m8ZDb7P/j3W58pF4ElHYqCxsNxzSnmOhxqoUxUnR8/nzYSxwdIM+fgDJrjVvEml/+LLeQLIyrJUS
FI2XZXN11bMDboeS34rhLmX2nslkcj8q9JWY5Us94hpnP3MkdvCb7GvGmzDtsNGfojkFEY5Bkt77
N1lIbfxlmgRdtoEsis3gvhwF/LAp2JmhTbD/TSbPytProf0OjmuctCElfJ7IvUL1MfotCOiU9+bF
y5SvbCp57Y3RV3mlYuUuslgn6L6Idcx19h3QqQq+AexF5jbZTGK83ZizlzMQBJjjrv6QCQxA1D2R
+jy70OeKcShVzAvTEuG9nbnvFKb1Y/8cl3ja4rwTFVSKbzrfiH0ML3DE1zi0uyaaBU/PRRkgWvF3
yT6UefNxF1O0JZ6EO8ysG1meB4kO4IM2V9mSDY0P5r0d4mxgF605p35cULfy2lVwSZ0Nfk8dl8y/
T+7jmlt1/nB3TPIDcrLVZCx8BgsREdCj2Ajjw6tRPxx3ybYYGjmV25ePZHHnB6DLleSSFsvUGNUy
NDj05yaKl/sximEFI7d2YaLaHKVZ0QOqYx/IFdfnB4bI1tXrOvAtzyHDOAoDuBfJMlA+/UoDkH7j
DOsrtRvMq+d2FRI/qaLwHxyWRIu3lKzY3aQ6XOTpFuhwsLOK8x/uux/Q+af4H3d8sLG7O+kQmMVE
PFre1jlwgHnGZvpS6TdAktr+j9MXRBWpG2dwPtwlUnVvFeZSM72I0dsqrGOsTG2oGNqJt1vOlJPl
WUbxKYkHbbTRvyfm+5nkqPJsOg+7RtFQGgc0j9pbYnNBA56zSb1eJdz7t9FRM+D6p7ttMLCQFBAe
NAhl69OneX8YkgETkjE0rD5Se3UH1hDeyWNCFFt+NpGQDkicAS56q7eT7XfD++gzHJSnhBwCdxNo
jc59pzfNG5z+qu2I9wGS8hbTVJ5T8DRkLEewJ9RIaU6Mrc6IelOg99FFuMtwNN30noEyfxeffNYX
+TLuf+zZs30lVt51hyBtGAuLKokZjNDQd0JvqiBJXNwdAuQXEK7zprhr+cjyUM9CLDtjNH4+EkR0
rvLt7T5b0h8yocTpEXUHi6i3+cWCDxql1PNuOOXFbO9eTfMMb3jVaJG/zu0b+lKqT/E3hOCpOf6D
slbnpcfNmskf54rzEYrMBKo8arLgBQm3IwW6aF4XHX/M1kosSJa318lfcYDs6LTJzWKHiZAOUr86
mzmK1gCZbf7z9ZtxYDIrLzNidvkFqVm+OEUKVs9Fwu/ai9HxgFiJ7fqP9M3UL2pPQP90xMufCHGn
ILa7GRlbIQW4AckGP8cVv0XlMqRuqWY4Rmpu0Y+3S9eHrlBS16Qxh/xHT0g6/f1Q0NZ2NDstKwQ4
WKqSeQuf3rgNXeIcfkpdVuZD5K0o58CmRT72JEQbjkLIIzje8Yi89pnCH334v/0CEeiPNGZGGOHb
jOhzZpAtL+EQonsuyGG9txXP3sk4/md5zmXQpkFQB5ynEhkDrvufxr0j/DwKq3Xg39NY9Kqx7xAF
KabiR8/38Ni/VngMoXI6zC3jvFwhQalIwqUWAlk+i0eBhXGvKDjhmbTUED3XBIvYq2ulYHjVyXFL
+KJCcjeyYCCns0Me88hBciFQTJ7s/yhNXUm34ae2d2KkIoeLZomJZQWL0hGZAKV3Dme2hNrobx+/
XXi6Xqy0e8EupUAinyO3buQiZEXT2PGdA+NyY2NJ6CUWs/1ZTo/VReOc6zPbRuyfMMNfsLfSmbVd
wX64xtTgQFcUr3Qp18dYIny1dYgWK6asfAnKc0AH8jQNHNENh36Zsno8n03oPbuh22Hx6qsgZuVJ
JdLvpQC6wnitcwlhbDIqNPTakmEWGALZR5qfM4xn5vsaLeSb05fayqZ/UIYApbxBDAflq1SyTEQx
Az+qnSnS86/LaD8lXzrpiLTO4pqDWNAGFZ747WgO46tts5ktAAeDopsE/6tjX7jk9dUJPU+X12/d
iNpxKU0cvEk4pL6I7eNKOqH6e0mRGQc5tmaLxYyEQqb9HqpFvFSekiLSA/LkAzC+8U6acop9j+Kj
nfNiXjGanqrlAntgSjPQvFJHZMjgzr8kGcYkVipowRZB0H4pq3+bKXbJzq2stR9nufGpRuXPgcbk
IGSYqXAKmGlbvGmE1d/0YxGuiOVdVyvjatWqPHdx3ocs3aSYM0xxLcPtH56LoNT916787H1QxOY8
FPFVkeqAIBwPLMVSnorJmpWWAqpRi3VxwpLq/tYPgcirtEiYPqws0/0k8SB4fA1F0UpsD7snkkaG
PPsM5CpUdTSsXXOg3lxcwQoBmipxJZQ8YsWtY15lhB+RJ/Sgwf+4CGUN/dK9jAJozBb7K68NL7C+
QU263j99Hjwdk8rNlkvpYEmQAlnaoBzWZLHHSc/AAVVYBtAVrlzKII1EY2mbtbRSKiCMEAP2IOFL
Xx/CpjLas7scOczJzX+8XIMMGH3ILS/EqnzMS4TDRyhFQpxVeZ5M92AwVeAIvezrfRAKabJbDSOB
xsXIaKSc6SX2H6iKHLMR807PlL5M6f7vXoBDDOEdBZ2psAOeXaIydCwdL92CPpGIlpwwX6V9GdtW
UrQwsIAv+dsHpe8Z3sgWlB4teKIEt3lvV2J9rqpmGPAQyieX7bDdnhwasqjwaku1jMMhiPkomsac
AdGtN8207mGlbRuRhJHuRMVrwdSata7q5hE8WKaHv6xcnO4xo7xj0VUZX0rlVHnU/xDi2OxOLTrD
QMec2tp9LH4A3R85R0vFrwokVVF0ewq/43YoT6ZXBmLOPfExQ+TpoyX/9DkT3yOpGqCYWwTLG3i2
D6D7ZmIgZL/Svt1ltyC3TR/NzrvX0748G7DTlKC851MbV4fyDWEudaVExDjcDO2OIKJGYy5dpLWM
WbpcphCEoMlBtN0A6h8fZtBHKdFsxJgiTrRO9pxSGgUY71Z1+TKJWqQkIoLTUNT5pFwvaYwzt2KO
XubE1Lm/4+aVmW0x49jUJS7DtzH6k4Q/dl27dy9wt0QBmVaudKjb3nOYqsu5EOo4AKTlDeri4c6c
eM60l5v0Td4u/P1LdggmXkIlqjLTiKWWqs5sl99FoOvBtgpqkiC9fKJdUi67SVAAYa+DH7inC+w8
W7IlVHsxy+l3KQGI8hlDLDHjBSDpWw9875s6qoYB2MwHarXBCy8ERf37LuUeGiDWVcl2GGsubiMU
b6C1BOmDHLbB7oaC9GrVEPpTLlSs2hHVnxam5gjnUuS8hWp5LFupvhors5IqY0zE+8/oUr6Wluoz
DUA4F1FBgghew4neOe5J5NAtv64P2iMBySwRbhMzT4lDYY31KZHkruaWyRCZMEh9IMFTCU6//ZWd
glyxnbaHM41oyimSSfuJoy49g7hP1or4hsT77/mIgiI/EnVtbHtyoMFcnp2H4MsLm3Bt23IYzqUP
VYlrTgOb3STySSjyEwiEXRM3jA9guGSKdGty1/RhROLPJdAGcZP92rBXqopzGg8cHbpA3s8q2WY/
/zGRzP7FtDlZzr+3zmVn/IFA6Lka2kKBJ7PjbVNIarH65GsvhV2x84Rhzr1dU/lA1+Y5JncJV1KF
iVLgPuG9xN15cJM+D4CVcxQoWhofiGpIctT7kZi2QXV+9fZ67nCEXM2r1KI6xbaF+pC84QhEZKcf
LBV33Yxz90hJsC75pG5Tr9zZ7RqcQDBmXsh/GEcNNYzSr/qoOttKxQsx+JLbrwkjcJPchh6U5cC3
M3Gk4voKZ6qRN/QKBTnmx7aCx+C8DO/08wgRyDNzise5aTlorAQWrEo4BoDQqGqU0+en1mQYjN/t
8QnH0/nKVlpuewNHDhEJ/EsC/uKI7zNFY746ZjakiYcY3x6riE7x3s6moCTw+hVltxNExmuSOsma
3SjMLQa8k1zZ6ZDeHKcICyOqK+VJ59Pw+2qc0gKqxp36uAfGbic+4/bjZa7JVd/b9NtCMmRxCBV8
f7goxCfCHxPv85fR7XOZt3lqJoAkXPBrM3jv8e+EtvBtkNCNun2xQyCgiyTEnjdoSyHjK322xnZo
KHjG+xu6/YZjtkPr/rMSnV89VsVa280H7KkW2zRMurCB/LEUzYkWir0PkbdBIf7utmxtVNE/r2wO
y+QfrQVPMfQ9doseJqAbbTvXVIRDX0Ckuapsmw9pf2VpaV4TkRI0rhH7H3aqb3Q2rjTsuP7oaYi9
dHSz1KLViZKqkmVPWHDC+iN//pHCS88Zo+ihVLT2VoIZ6/LplGLP11Dyt87EATrnU8tcCjnT+aOa
kOGtvecT05iFANZ5ZtfbM4khIbGi00tBicHpX6G40s5NurfedulAUHNPsq7a1CBdEpkA+yJJKuWR
debRbHhMBw7h5XIxLaaCXgRqfKsGCyv4xBogoVpJmjjUUmwHcM1QNWQEYQ9G98t2eqqFMDGJe9d7
RjMA0Hq55pg6CINugeP6VYH115mfwU0u97f8Q9NzWlLMKvx2E+tDoQnqkT+smMbYhv7/qEkcKO7A
aeF0AXolsUIsvWU82fYAXYNjfA3aMz/wn+E8SllX8KmiEeB/iIcW4RBbVYWxi7S+I82qJ+8eFlvt
ynRWBoApFTjTerXL+catzVUEJMrHd18+J1R0DZsdAYxXB/gyEvO7wKDniywyKVQ+CsYaTmq6++V1
M69BCXJ2HkggtLDgTfMvBYvo9GScX1AZfy275RGj+B9soeKBThfPyAL1JRnTvNbr2vyEPBwccogC
XeoAMzv14Qg4D/cnqowpyvOb/2H4xASE51S1/7NeXo7Wx81VD7ohsGaHqqJemc/DPbqefIjVsfKH
/EUTM0z1zt/6mirKTRZ6cksPwIUN4lykH/OF//4rfTq79lTXyUlrq6pBN9OY+VrQ/TCf7Ie02TgF
wLIax4pMywR4rn8rzIungOFJkyJF7TFvlUtDr4M3Sm0TqnmvVwLeBxzrbrnpthACjGgZevF6swty
gAyc5X8xOkQM9ew2HvIFQD5ULKdWD+6BznIwMvpiZXkQacxx9kNZD0nmZO02LscGm0r/Xdpyk0zB
M+PJg8Bc4YaUrQuCoRdF4W1ogqiaB28FB78AG80s+7OXjVUMvPcaqi+gyRoHabJbqx6XkFM5q5Eq
4z3PDYA6cuKsywh49/8eEpnVeXZCXQLSpp9/A0uHShQJEdmfrtS9DwY0FzmBVvuqt6uK+p4d0EsQ
TdqZcllAP2F6J3+sgm8vaaN7aT9kZ9ETPkFPBBpFhLgoIQAQgkWdBbadr0b6f7SRonRrAOvKerJO
Jd2v21FiPULd2OkZEpWK1rThVwcGEFTGc38i9v3Vf582zYJU4AMuHvW7V7WYlub4Bt7xswOZ5t8X
NKoRSbSesBnHMLm/rQZgiqPUxpin257WtOcfhAjVTZGn+PZChwa9Yc/E7vCVEu/GqBQ0PhSOcJIX
TW2QaWHouuhv6mvxudMhvfvk288+K8Umc0DIvx7CsUgbUpkV7YxEhRUtofq7j4elS/XEGDNeHp9p
NrAzgD53sgiIhKHOdH+0R7qjlYN2MM1aTwzODemZfsPdEYw6xYV1psKZqSpyDrPuT31bPTGhkOcq
BIvKtfWcTF0Gex/JK5qYVOkBDhUhm9qd82hE3ShVirmuNOWOh5aC0TttTQWP/21G8ucIrZyZMOiP
NnvQepyz3UQDNMcqrn707zj+U9cBtcIPScEjXdzo5RjKJojSppocfHctkcu438K9sAGzbOy2t7/J
TeGQDdEfhtQuweHRqCI0OnWiDBc/u4apSrMzxpxGVgk6OZrw/yeoWAfoSneQQ4TCLsnDva9UlRnI
jnfw55/gtYS74aHYVwEazk8NyQ8I3Q8Mk0bdGRWdWDAUc3i+eNX60zQq56UEfBgKxTtYwKC3V+Xm
IFTfIGTpAR3yVY6j/PG2xK00jSUHzV7YFKR2d+zHJ5W6d+sKg/cPAr8xJS43mW7DwBSIOOqcPaud
S9EUDKLndoEGsTM+1yzNwXVKeAcRhSzUjZX1D+fzKBT9Rfg79tQFK2KRGmfn2j6hm0RQG91vX5KK
xig2VLTQKZKE9OcK9wEHE0p6qvHyooGYY6DI3WjHK/IRLNtPpBu+ZMK/xuL0idNJTpHGbmKCq34G
3HORV0Lg018PVNzgqRTGHQh9mD2TJv6M4LBeE0NqJa8rNV3BAYzOA27HHPdklUzB/PLreEuj/JRO
ltjmoYcyiPDoNfW6hGbIGAgwLBOX1k/LzI8Un0tCg4JEk6gpNOmEnJB77GGD0F/yqRLSHehQgBN/
HdMXeDuLZem5OLfKV4dG/y3dFEJP0KqVord7OiUNMcGPu1DPD3tBO0WR6Ah3nU/0YdHJgple7X08
VXtDNvJg5jYCrbMQSiA4AIB/Y22pAtI0b14+NJMQ3haFemZC06e7PRzdp3immwgMJX4VfDIRQS6X
1eRVWeXUHHKoGMpv6aeBfImM2fUHP2oodzb1GeYK+EWkPMdZPJ3RZ8bvT8y9yNI8t+s0ce5th2SY
nvW4cdjJbzx38mNJr31Az29pmvSlJJFTbmJr9D0gJHNVE8jvlBRbYRX4itPg+M9E3QGj2yD0KmqX
4+nOEtIQx5XvZmSLToiUROdtZj//JPfVIS94jAESxPpImfqhlWtN4D4AOzEtK3cKTuGzNkU+eZEe
KuRKrREdMQ3Ud9KygFenkRRUzE9w3sUX5vvBwZJbW5ttDjZJ8iQPtBSVFIuk/6hY58uL/mbpjo2m
Uvdfcq/Sgwi0Ifhj9qBIqp5sO6hb18j1dROW+qg/7CEv7kGgHXNItwd1jMbKbwJY37ORO6Gwnvz+
iux9WY4GSRAR8fLKT2ER8wx76ND2Y/o13H7Ht/wGgqt2por6g7QJyd0Fgjm2j4ieDSYgFIuxcWoS
29d13UvMlM3n4qen0V8Tj3YyRwzg3sDlvnVWMllvSvMm6kmznS1qhU9IEg0mAeq5fF8QPxt02MyK
PPXmsaAFdQw/B8K1S5I/YUsJ9AnSRK7R/eGgjVdcY2nB8bMG2PUjNwvaITMyO7OS6hKrwR8sRssF
mkbnniFrXPvACkDB2RzA24qWx77+nDencU17lOCBNmJ5BoEOgK5szTijwzRY01cDU9Tf+S0CrYfm
jMA8tvlQCIRdBUzQWr+mhnsB7SHGZpf39bODOXXWTY7bOX7PHKcqHfmGUj1T1081qZTJDDo89i1B
yl9sjMrcqgwtR0IY2i1SCBIQ2ApgFmxjaS68IeJ2k+hV6GwQR43jJh6ahpTqnNjJ1Op0biRGk48V
fVhHnwPcTXV9q/avG9F6boRp7mFyMAluBE7YWqedxI34NnCYGeu0YC4Rd6BF7KDbAwnIGoIex01c
ADTgEqAOcWzoyl4DJcVdttzuA/G5mUzmbpEW//QhsqNM04+O5dDpVs59Z+CNkDthBMmw+mjvNQc7
84dOk6XX0NgL1P5AKsOmHZ+WWtnI0ollgNgTuk+No+yHurpH/4SE64wgOpxgMahB4jGrLVaC/fY1
speO3nGuYKqz7GUhcFn3rPBD7K44DMmuWTkZVIQUT81yTkR7VwRAj31Q4juvJYbw2Pak8ltpZmJC
Zl+kDWg5AAyD3Te+qqSoYtkTRsXw26Z+q9UDLpaEDmgsiKhJLP13wAGgZLIH2IuL0XhSxTUtbp9m
qLEG5T/ETG/bdlACMpZX1kjwp8IRAnrZlKfQbrqbtOBA9h8hivdDQni3TNOEomkTFA4gK1vbXNRi
VdecLby7uDCOoMwyL5Jd8tEyzjQvwUNcaZ9OlG8BSsK5BGZdgfScJv9vlo/63ofeATVKYt1LjAO5
AgO5Ot/vvzFBiJLdfDVInJuO6lrUMAQ892vC2BE/NfMr8XCa9PviXTrQ3LUBfQ1+3w0lASvcP3H6
fAPxt/1HXNMsfegiyeJzvCgBCeM2FPLzBAaUUj9uuEmsa0uqxGHt4FonKp6eWDXbM0gwgkW62sQP
9iquT4qUOnIDmrbMGObz2ugDlShC0bfIVFWjEAU4vNB7B8f+zUB+Hw9r8Uk0e1uj2vyK7pl+8vAG
WbIMNwMvTuxWHyAjfku39FKqU3gU/Wle+IKW4sfqJBUy8DSvlaHDeLBx4Z5GhDuq3VwFB+Cng4Ix
2uQ4/1rhgPY2Nk1d/4Ap2Wh7ziWJ8fQPuApSyvvoonMGBjZ5O3dsdMsaj8lgVjfl7K6XIBfsllL+
JJGswiFyl5T/KOVQqxyJx7hNlAolSFsqhhl68qUvHbtL15aO+zEQ/6qYhqY9cxh3NZuXvWH9CCBR
AN0V9LJ0ILlYPDeLrPYSSz7gI43d+19YI359hrigg2Ktw7F9rF2c/WHmrDt3V5KxO8Kr+SVGgmky
VNoywx7BLyWPW+NO8k+a36e8ITV8zA7gpYnhdIJQwsJhzGYlOEiyQNqd9422kkMe+JigAJXSOxJr
n1BKd6pKwaNwVVTzIfkb7XwG/O92Bwec7jPzDAbLKz6Kr99hltQ/WKJpinIXTts/RgOIA58lUYp+
o4ruLuZx30osYwZwS+G6SDHMYqB7FzJrwAKZ/A3DVW2P0sQ6PTdaeA33QVKHF3NcaU3Zeyu/qbin
RJmI85YRlQncOmIK9/JMC45QnFGuY6ySnCgNWlaCoxAr2p55Naue+8FLzojgK3dTkz5QKSaNTL90
3jzrFjyafpBcpA5W1ED6ykUK5LQNIW9gab32EOqrfbGMMrAzSdPu6BMkz9tkVRf01eC8YxdUaE1n
MTi9QTXsjAmMcGVL5WgXrLsLD44zFOVVWoE41AXxRQCoSL7kStJzEAJtEUtUMV+dOztJ9+e5gFqB
wZcR3S3LlQAtB08VpiAFX2m7ZoqRFGJCUPbCmNBpZy7CAj/axEUf0Vr0zHJ4Rxk+mG/bN3/1HnDM
42RL11UKakCItWhAwG7k+3CylmRKcDt4P7cDeDmlG2p9UQ0tfH5fhuhO+R0WQ+/B1i1d71kCRHd2
WDlNCpqWCUoJsVw24SXO7q706lyonIjVntVcPGZn/F/qQqFLxsPdeOWtu/bdpsZqtyCJJSddCXmM
ROEtDFmE2ViTQiLsCnd3j92WxS+mJCNMj3V4V0HwR9JTm5XroM8tUKMNsShgd48DRrPJDauScyUv
TsprCjipfGO1MLz+hcLegLqX4AeOR4QRQDiPKP9uqY2kKUgeU/cS3zAOVyEJnBDZ8gz0RId5Q7BX
7MDDrGgblyPOwNU/DyNvfDkeibENWFon6vNlWNJAtUkq9h7HO16/RPfwAzjVQ7tMwfJ2Gjl4ZY2p
7yxcQqx+9Ybmuz+NpDXosgFDH6exelWf9Uvx1r7/HAdb7WbVaObvUATQgPfqv1jY+Pclyg3vDF1x
ekieHhS7dO+N242uRmQu0Qyor8e3LqArysOsJsWPkX4bB4SLkKAhGQGWQYho5vVAn+tJ/uouoUlm
mArBzMYir9ATY/MhO04PkMi727LgFaS6QSsyE1PH0V0LWKXhnTcMcX3Eykf4UVSsldJ8u4BMRnGS
jML6mugvSSuujtQReEWhsJVjcruVKSN7WxiNelkQk2S7INGfN0zz9aSETRW8AQFFQ7RCzo/FfZGy
J8zlIYgrnnW7MbXMYrvL/FQ+jFo99Myc4BjiDsBvmxXaZq/tDUv4xuUvePs9sqU8At/cwk5IUk5J
IiwL2v22mMuMepbngCZb+a4mgWzkrshWf5cvJxk98lSdDt+w/MOkLii3hzp8PBrZ4WM0RNLMqzYR
04y3Y099o/llJeZcTJ06nCARCkEln8ngf4xF4Lm+5pi7oFKOeHGXZMK823z97+QDMEg1yoXqm4uq
/LPz8BoYxZQ+pnSk3aTt6SK6cqVX6ZXoq5jo5W+CnddNLbA4PhZ9bUKyjeNfvWFHM9d4wdnlXXZD
0BoNy1LwQH9bZNDVwd37fa1O8aQD+VrVLYoH5aztqxDtmjn27GSJYo46aIlRTyZC3RTxGt5hSFcT
6HQCL5sFqZT1zHMMeejZX1WdFF7dSc4pN5TqU4z1d3hUnXyYpufcbw43e2iune7yEg0IVnjiwGL/
uaVCdCsm8HZexeYTIdj9FZJ5LwL/sBg8g1pgwU3HhZxG5UZGR44bFtuoA/ejQybsgJyQ/a55L64o
Zypmy7Xxuk/YdNykK9imxqnJ9eauVL/9dd9StCRKGM/fmTffiuIhZZoM7iEW20H/42vqxJZtF6+X
Lh0H9Sopxv6H1B57Oyt61WtrMQQX7DpfWhg1mKLtDKCjZcK/C/k38x6qXxSERPzvN619ITHb9E5n
yuR7AKzHMGYE6kKoVXGHMcOVnX/i80aY48VflSZIH+Ywlx32OmOU+LB76r0+XMIB0NNaLt6W8o4K
C5nHeS/UNpVb1wPFAmFcfipSOS3LQMWYQ+Nk6vJ9gPPvrtMj5Q/1cquNQtQ2Fvui0FXh2AE83L5G
DKRG+dvMx3PbsPfgVTsHes1qfozYds/Nwy/jhZeMUXoumJZuguOJzort/XpuYZXcCdhaETT9SnJs
gL5uoAcHWNVskIh3uctocgcP/gAhl04lsJFAlRWpjSKjja782nycbDTbYWlVCTkzeNj3eVg6s3Kn
Q+ZroNPuqgvua5o0dB0nPWXqNku6vOnvSr7Smts54DJeSJh+lPPPES8QtQw/qE/oMaAE9h+/Nz8X
6dOmrE/SwC2GNtWUao207kYFrDTi59cDCrCg8pnHZXNbnyRRrG7Zr1n8EaSZM/5xGxl9BZFWOjBT
V24MYKtUa0Ee++ubd1pWkvEwx3h44R7wmDfzvPOEM+0n4RBnbw9pSY6o3ioAtQgIDNSQOPEUUZtq
dxxdZz+74xt/zM5KKQBJwigh9V1XRHfLOJ6C86rGMOGaT5p9qVPpyjGlTi1td2BuGDNaa4x7tayp
kKNm3Jp+khR5KIUItR5rqbu4ytzGjHCy8ui+LWrnFya6QMAOD5nvE1R6zp791nBrY01ZeGTWbPRe
ChNNyJKVjzYcc/s/37isuVCd3jN16wJGVsmvnh2cVWV1fVkyWJGFZTqdtX277bfWxbKc9t8hPTPJ
duXrmAbFYZPVUAL/fnpw1WPrEPU8PaZUOFgz+obPmduUDOMoIOYhrfVHbzH9PUjxRPtkeAGCyRvY
mLJm6vBGmUqLaYENUfnFQ5LyEPbEP47d4C1M0ACjDoorLWjXrrYcBS84SC3wQaand1eozznDA2x0
dkty/hcShQf6dPmMVlVXaAM5j+kB0IdrKzTXg2jFkMGT8ykQT2VqHWk2ASFT/VAaTyj/NYmtLjsZ
xp9iFoie6+4/VK0MvvWN7SBxwpojxuDn25BPdPwEQ5Fo1qQRx5IqqcBB1JZcwpiMwM19yzcs2YTu
pPvOn3/5qmUeiUp+7lpR46kNqRZHvTOnQjcTsEwBWzVxhUYerwnayV/2q6KS0l0ZXmwrhm8wcCDN
8LbIPn99UgSC1d6BNxO/6iXL/CM5nkqRF6dJPON8j68GjSxZ6+MUJHuWCeEaWfx4lhCcurWvK07r
8i5wjEdkkfIArCWGJctrqlbkA+5mtarpWUpABpNpN0Nw3MZwjWntaqO1hKPaR7ossuijNFN+FC65
jkhgU8G2G1FVG6YC0dJ4HoVhJ6rkFNeZse3DABkLoLcl6sL2VZmrpd/gwgujSBPfcdnvmMOWbxIL
bahy+PzViZF39VO8DIgKV9S18wszIQU4O8I8qVmnwxqroWITH4SJf4Gw+EM+TWz6KXzAky4iN3h0
CecgvqWgaqkdL4fvq1AhEopGIPDmSCs+tiVc2DxGCEGtHrEjWprbY+jwpcc7utQrBttJWtyFt95+
Ap9UltG+D7w9e2+pSZjuIhQ+qj+9pn8y7xFI/+8nivQlv840Ioi32mDdAtuQx4/M4skLfs8pvxev
9BfuCLNd7RPqXn1jLOQRZzXEupGoDaqjbzzDjKxBtfy+v2kg2xtdpWNY110miZ4PoKHYDqzD9boK
/TynstU7btYo40dyKHzpfYqdTWbf1bGMY66x6q9NxEBlqaYszghYu3vNvLwFLnFWmcR3xGZa8Mpk
ZJUKvbbQtwkhHW9dTt5Nk72u/AMlkifBF3tJrSm8IhultEyJU0rTgrLZisebHZ5I/fIbb1H9tc2k
pFDbxwNggasrupr9WhVZqNKEyQ14SRvLvchHIpvi+j0d8m0ZRF++xbmsZC8Oek0ojeq+gG44yWJV
Kn+OKxASBhuPiiTtLcE7xM1d4vC5ekD/J/o0u/FBtgzXfOzOP8lkILL9H/cLKi1smztomnxaI3Lv
nwDmcwl0m1a3p0GA0TPKUNTTOAyhwISX8sHX8Za49Dj14+grn60Td9IpA/MM3Qohc0NWlPMkoMYo
rWOt+Aou2YizNUMOZJoEp2wEIEk7oARNxw+KwD7Ir5faJzGwIgVZz78yl6jS90TTR/yI/WNQ//lO
l9557vS+z95zqyKlzlf2B1mveAmTApeZne5e18ywwA6jrWHir5hCePYLUYIu0eMK0lBhl3ELx6zF
vpegtIlvvPhOJ53I3OPuxC3k1lqcpHn1yZARuvtrXv9gpyyAgstquYJJSngbRYocwhnFqcqNIa++
a25/Qji770EJwhb0RIVXVSjw7SfVHP8S9Q4zLWk2mhfzi25miEudpuCG9U7gbsC9cyUcSZ+xB0R6
GgP1iqKZjrRuWalMoGOKAVl5w13kpTWKNzcu6xAhT5dj2nl+7nXOZ/JJNfAB8AsDYM8VB3e7lxk+
ip0wGi05QGO/ADMv4eF7J71ds3TWvNz/Rs/Y0dU33Kf1okC5AuEyLHJwJzSDI7YIH1lLIf5Eh4Qb
Z0jm0VasDM1R6HkEBMQa8WgZhQ1LJ1HqwZ0r2oxpOXlYqSjLHHzaWQ3yg4bm2AB2OSreEtplQTga
RyQNhNOhiSCVd+thsMu40WCm5K+9viS3PhjWxm37+LTVXLTFA3fs/mcW2ChYwn+gAntYAkpIXw/1
reHS7nRSkErDGDgl4jhYfB0Aqwan/vv+Ofprhf3WF13APouypOyDv4pPcL2a4vGxGZwCJL4gyM/B
VxbIMFi3L2AFSGvWqFRw+Z2LhRQyCnDHwSuTJehtYzDsyCYhIE83ZE1boDE3qyM0uJTP5+6se812
JYFHk5/p2DFydn9BN4AcCdkpEoIPJ5kRYSDTWVw3b/mMqeFvms89nBHgE6+e50Dde/96QW0UAt1H
9jIFXYN5/KaMUeVWeUlmo/O8MdVsgQFEN+CAKV/aJ3eNorwfAkoJ7uoKpD4oOA/GD2vLkVPAtcbl
/9rM8u0BP5IIGefhNM6C4CK+uBifl2QQ3KVR2ZwJ6NMkUuVgLxsmbwsRc5sjlAi+q4SOXluKLilQ
lm9zWerH8x11s/LKWXvDrLPnQJY/TmKwpIP+ObL+HlyQlWZ0BUcPIZ1w+ENAak9LJZ4OEe9UgJgt
dReqSENw69wGstJwj3WMriH8+1WT2Djq7qwSfDyjwVYBXefoI58LtXGyF09EvUscJp2cv+dQtgTR
YJlSkvVwaZGs8BBBt2TL38BRhkzA4Q+ykPoBjb+lzEIMCHV11+0K2wi5TAlYPwpe15Eou3dfWz1Y
6iqPy6woXxcFnluarg9tUk12P+HwC2xauxirYGWbmu1HU/jDOV4gwdtva9l12K0wu3ZANXtPdHQV
14iViaWraRHLWpvAfU6qYLMdBgNbA9LdIRBdloe9a+LWGLXumcc5Jjxm6oEQPV7vKcLl19sODbHD
EeZ/lCzRV4IWq/OhhuFz3jMmORhfB+lKIhKUdOOqN4a1jRigUNm4z5HkcIYCDW6lMWIb9bNIN2PC
jgyjG90Qpy8V2Z+ZEXK0tA61xuHhUsdrf5zhGeWEGyR1Dpq84eFIq1yWoQ+eFQcfZBHwOwhuXFup
c/19Y+UwLAyyRIyDftiEfZ0UuV0SqDUTk4EbuHeth7O9iV9EQHEmeKtcg8Fhz/XpclAuddjyJ7qJ
XoElE9yl1XrZqUIWrafpkTtGkeRZi47HUOYCaSAEeSjef1cZtBa5JC2gsPyv1VLcV6KgnByd5Fq/
D2CFp2DbtbEcZNsedDFbgKh9CTyPCwH2r1f233olSmd7jHMBwqSMt5bEFNU1nx7yeQFJVnwi5kMb
qLFwJqRdzrUg6z/QMM5jTX9yIr7c0/Q+UQAKg9kAbJLklMNPZR1y4se60cPrTUh7GFX/gXzEzNNR
SZQ50OfwyAoa37NXWtA0paTvP0S9Ld0fy7h2luDsaTFRzBWPvRYloZFzcc1hr8kj5sk310Ou+r5A
2ewCH0fMLBCB/SbaczEcHYfQrGea2ieEgHK0M8YEHDN4/IBtT0hpp+QR66cRmaz01ZSBnMOFsm9h
3xL60EgyP8F4OJsc2J5QLzwGMl83txvmWKVlRWzrMxPV8/VPeMok6BPElG2Xqe+xnhPpZroZf9pJ
lSmniEMckSwYZeE7jZF6gfTlcYTF1+UKPclueHmRBY4UY+A+3LvY942xhQ85/Iqr1VW8h0T3KRwp
xX8qXqzN8cQf4oUyRcWqYtCoukm6QMBsxsSkcYGcLSVKB9gTMx3ZDqQz7v/sbwK8Vs6jN7lIA4ZA
NFarPWYbXgq4CYkniXC10bGqTPqBLt3yLznVzkdYx347jRA66SmVA1278bPaQ4FwJ32rMnklu4yH
MoP75Ai8SNAO46RxikWSTKrC/wNLQku92Gd5L2euhO2L5DX+ka3UdBhmrJa0DZkc7F6G0dZepgyX
KBs1CfKolKIAP/7BVOxLFvXBuQTz7jJZCFmyJf/RU9TyIvyyQ+bn2NTsV/X2kQ0xYI0Oe+biV6ez
74mqVrKEJcQgAdwDmV7avuMKnhJkEgdo0Apy3xNBR1B9oN4MAb9ExIXvxdWUhFPJp6NpYlAAzCin
lkYFeFDC8hH76710g55vMdM2DqRT8p4R4H/pSHccXa4y20iQw/ToUgydk6SeKhSNYsXw3LTRgYxB
ShA7Hso/nwx34dX3Z7JCggu7UQfZlhsHh30D3Vct14CnWA0jSRO5e6LSmX5CIwH3styvv3A1GoFz
sigc52fJlzawWKNGhGdyW//nhRVZAdI7Th9cJoi3mq3vlF8qzvdpN37xmyX8QxlNIKkcyiG/7XQo
Q7SX4RJOb5L9/1lzVqmocxfG7bGi9Zwj8nRyQzNxgEVEnus4eyt12WaFlequdtKV8oKgqhwTRc0B
rGuDxXDSujBOAfiVAZQePzr9NSwiVvUgz3S98YLbtI+55qlpXPEoxWVoF45VeGbhKm4fE7ONmGQI
eKwNfP6lwUuI/oPCmXOYEEha8KCs+F/JxqkDIGTGnD+qCRjucgngTdrNoc56FTPEjVPHK6MLTCH2
xuf804HnHHhII6js8PBUODZho64rsq6em/Slstn/rM7RMLo7uIqsbtSaQiR9AJKdNrGC2L+78kf4
eFvCt0GaeM3C1f8ZTsfmNj5xDMtl5m0xvv6jBjoU0vGf+5tTCOUKTLfe3PtffQeAg9RmiHc/X00D
pxYlfl1ZH7YD5bHPmCCRDHal1BMx4AF5kbPS+0i08srpihDwJjNMI5W65uWkPKCNXMeWYz08LXi+
W3iR6pYB0xwhz8Tw+bNJV9HGTV/qNqrbrDE9vlmdqx4GajCJyEHDnCYtOij06Oar8a945TbdM2PV
IM3G8Bqc6q/NGCeriVQ3/I69Pau7rdGIMdUZIn04hG045u/4L5xXdaVLB1ss6sFb6N6uxItZCzbI
Pm72l/iJG8nUicDp8RRUx+7KQpkg7laUxgcSzyr+YxvkWwsQo1mGDUZAqA4f+E7x6sXPiz4Q/6rT
J9mWYIs9ynmTaDcrsr8aH7jH9eAv8f8e/HuIHQ+GCpwyBsMwbicuF4KhnrqgBNR3wPu4PK8K0Rsp
t5PRGW6IjPyNKrgG8CbJ7CG9F2JCAu5P4IU8gq5I4iLArCjNFqhToSVRfT6JsnA6uwyl3M+J9SVd
ya9Tc9wUhC5ZO9+nXNtP0a/cAr+czw+yT8AOm9yZDqdk5+oe7N3/RsgGqipgcquEqrJC9ZIzp98y
8uesQZ7WcBxuD/V+DzvKqqoA05DAnCl5Qp+QYWfeiKQhto5xPoUt5H6ecNWbq+Qe3cR4Vzifl7hA
Ff447uBPe2d3F4DTcZVI2cm/nNgtfpkJKembFrR/SKXxPWkUc49z3wCmBvqFUorsRL/q+OOr5iuR
LjjpMAVNI+ZB4YCEG1/Tfj0llzrxIUJCe3x1FRKxV0yxHZcSCAni0kO1ixvqXv6hp3bTvPLz0RDq
3b9i+quGx3l2+CSHODqYPADsT1ChyuBWcVi6FvhoF6WOEznNmGopTZQSpJo0/PUSjTE5foeVX2c/
8Fm5yCynzFOET/N/OqeJTM5t8JZZ353I+is6LFp0w8DQqopmvN2fQnnrgq/jdHdRy6xPeghpABUW
9lT6DkvBJKQZfZhc4q7nqK9WS8hPGZuRwNa/10hi7bDzEWGvzz/lpknWzFQAzYnHiCL6XgMoTSLI
9T7UYB3+5T+RkubwtnXUODFnjpPVQEEks8IrCiPp0bqe1YBcM8iiWg9vMNUJ8IaJCKShteFdPsVZ
XcE07Y3UP30DNYhm0ZdOOzi2F13T1VGhbI45sfxNKJ5ujk0k2KT0m9YOgy9kqGGAGjCg/NaOzc8l
gsB31/IMsPygybk/7gx3PIK3QVLu/igrIpS338iJrSWayJXrHeJPhjVM7P9dGiHXUMrJR58cvo2v
B7jqm8Q5OHx3kKKatBT7uBKXuRwLlw9Z2aW5OVBt/09B2c6gHlwnytC79/3FaSTXoJuYIEFyrNIn
7RBkKaHtCjgpJtpHGLryZKCW5n3PemudLWRE4NXeqSRCyz4/kWbx2x21wDaiPC/PjCRrzyNHySH2
IaVnyAvR7TdCYTiSdbsfszfH4BZYvHGKZNvT9Xrr3HcJs0e9yDsV3W0SOCI7j/0+cgXQByu3H4HM
K5xFJ5xvSq2jLYzx7xTxqkqBuSd3/VBY4Lfm/5X7Q2fNmZUGV5na8NVKpEDQsbpS9ND923/yPFd/
VwV/b4PwtQSoykLcCTZ/fmCzwVsExq4nAP+tl2abcluW+YI0go/1PMe2BwaS7GiPj2Sc4FzuXT7k
IC2i7lSEO7/eVZjpBbXC8juOkZUAJyYiQqhB4dwyBxqMl+xtSiqk1368sjAp53XjulE4TzdEzyFq
kr0XKJR2ac872OzT/8VQU3X8NupYphLfVUYqCZBKNfH+nw+sEzx0XMlzQXq4XnjAptkg8l0vv+EV
tjthpzJugrdtiqxJ/Js4BMWrUhg+OeNi5wU1hu8Tp6zvJk2pui2N+sdbunbB8bgesKkY4MCmOauE
u/zoydnZuUQZvUW779brMqom/ZoYSbp30ziirK8eva0MoVredKZqy65010EgwKHMLBgLcYRcYFFd
AUsQuVWybWZOamhgSGsD3Ld9HDqfRpZJsR9Cvd+vvT2e/G5pJgBz1zvEpPdFmb7R0mpycfGcHsdA
UTzpOVO2H23u1MmtdrT5ThPG17RAwHJYOA0we9w+IDrICJ8RGirx38Rdr72uHSTrFUtFPU+r+jYJ
g0RbWot4z3qPrRqkbUg0Dh7JsBBtzHelobHDNALW59ElUkHaQcH6sDOw7GN2fYu3/TAW1Pb/nwPb
Y8nn/uhcBfSYR/aiwg9hPmXTwCyYRVmZ9yf1dDNySJZupffoN/9A65XS9cZ0+ObFK8THEBGdb7wk
DFYYG6NjqISwZCozIDiyjAmGZWP2i7sUV6Yr7z7sjy64lOKqMT/54dS0cnup7X2pxUlXvQ2GMAGW
3jvlvEKgLPilg1VU1O3ONw7K3AwSW9QQardIQmYJ2v/NVdJ+9D5LQc/9S2GE4sKBMYTTb0VaHKND
HMqMwlx2lMI9lKJ1qizHdc6t73XLKxSUQleKcqUAEgQ1sjoDJ1VNzIROQyNnAemicohxQo00IdkP
zoMhzi7inKUVfSXlV2dTHP9C+zOdxa0MITS7tWC62rA1IdI0cKxj5DsvnEFsSoIBdMb32p3dgtxs
qenpbZotUd1xAKcZtX2x1TmBed2mXCgD/W5DJS7USJKVAGM0J1/KcFMdFWb6gcjBFVvKan+m+THJ
W01U4PUR3ZXQfjBy+F0mJT4ZkKYIiUYtFaJfbkQFzRZWHzlmE3qkQm1hucHKisj+9rbB77x9KRRm
pGeOtXzljed5dAnU1k9CuyPeiX0S2QnzD6S9OEE8aFop4lq3OQGAdzbPS1DP0ts3oBww8yQ782n+
iTvheQ/aK1VqlUIeIxNKlgFE7+N8HioFe69FjmZxoGijiSYjNssnF15eSmcRpdTgPTQ6JzF6BXaE
6sR4919FZOVNIzYFK02MCyVyrXt0kcKoQPwbT4nKgstFwDslmFvlZLeko1YeR92/YrMiy99D3hsI
SZnp/aI0b9zIJGpiNJU2Rqvu4zYpMaO7Ueh29BZ45xd0xUCV/h8aW0n+yptBulw3QM4Xzqv7RiUV
wkqXJpRW8flqimlHMca0N5b6eDzj6H/C95UTdGQNAGIG9iqxBQNciyiabsinK3JJ7C/UsK4ekSMv
uuSPWmMQLZYvQ7v7+zKAqWkLLkSWcB1QfcIXvjDMa39ARxowyT27JioAdjnbqedWCqiMavnqwm2S
oCzPYgLRs4dtY/vIKsc47DKL4jz7ZzWMPj3BFYBdp4shk9VIhs5dpLvVZbq78DFsGtIVRWK4j4H5
onlGeteBn1/UF+Wb2+lmp/b5t/OUjyJUZqOUhmXv/rD2gdcVvUUAFDnLqRVpCnNdh1mVIbLjRfg7
m6cSWckZAKY+FsBxCh1DMyo5skXjnuk73FCd/jvikUptN9MqmlFvpCR8A4qT5hoJz5pesnrdoNpm
Vn+YlxhrYGJihFMaVtCJF+24VzWdS0gxWmQICu5+814RFFhK9ZXd3TT1GFHQD0epqOIjCx0B1hsX
GrZrj2BWocHCKB1j1auaxzGG47GiWk/VNZJgxmqe5H8kpFriaAcvWS441FTcCx58rQ+PyrLGVBRP
DC4fU+wo5pIFONUDGTPu+o8rfCAwc85GATX47wQrl/xCoyZK+3SE+nXW/sNakeDnM7oWNWJLPReL
Gu6us5edn8wbjCFt4Y1jSCSIX1U+YFSAPzg8iQ6T0KZprhpaE7ZNvLKcc1j7AW8aTe5W+20dzypl
8qmaFSZ2kDXGTWdTo9yIOT57+X8N9ezh6S9CVrZCDdoYpnAGgRyDmJ0e3w0mq7oglkdwuVdc2+oS
YFjQXQ/B2n0nyNbEDGPe4GJjPbzqF3QlzbRCkqgSioUsXWbLN64aAh5hBRFmNgiFfhtfOJfpUK6v
WoDx1SBSWid+keCLqLwYhq18ekUmXadyBf6YMXv9kE2UgrxhzOpNX5jCZdLC1I8dno/yA1bdvHJk
bcV4Bdkeph8kJvEVgMSb5QETxgGBdwiaUgTo/nrM9hcC3FHrWDYMUOMf3SgMrC99U10m7g0eQJjg
vRb/nVRnE80i3g8aJLJM/HYa/XLVyF9K0cGoaqaCZHJ413ttNHboD44JJ9W5SEpPHFBbg5pnWZnr
/hPtmIlD6Jb1XwcRgJD/Konua1EdCWr6O1Hp+1IYQxYs4U+fekTMwpx0bSeWJpBQU/cUZuMiS9FO
/BFAtMZi4C9n0ObmsFbEbInUZAY7o1qAp4OxJIg8Esyin/JOHjIjJkRKtZ6aqeFtxtWb1LXqBWv/
yuyijbE9p+pq5d4GT3nZHDjkmdYaK2d+/VOLqTVEy+tYuux3CU6xaAvugi7byyBqLO3xgwva+Nx2
n+mLV1SLBdgLFf4FQtUqHsLW1CjzcSN+2/lyGWvw28/1dPGPAY5Z64f2LbY/Eva0B590dWNa3d0q
cQhX+L8FDYhMBVGrqIQM9SQiaMXbTjdHwrBHe1z/hhiAbIbFF/mU0WGODHLB4mauzmy2uBWcgmpm
OkQhYGQhI0ZNLoOCc77iHzoPZQm1TUdYdRz7YlvFf+v9n7hyjLEGFuY8jCbiB/2QsXsZmM9BxJd+
SCVTi3pr+aRXPmTqZpkWgQuKxH9j6nt3n1w5L6pWNPj5NZi2PWkzyRMc/NaweM42TFPaO3h8ufYx
SLMd0HOyOVrQqqzty6uaF5RvTdfuNSSwmgYTJzAyCBryGYj+6nW3UVjNSWLTxSqhmC34JSA+0F2p
Lv7JBn31ll38ctRpJc6f0JTeImGmeeYwMnaKoWbqEDdMFw9qXTIGMFIl5PVViIYw2DgjpM6wN/Qy
jtVoZAwvxnZelMHNUyIn83YzfKkYpDBbxGIKRuCJx6uCp+ydusSzIng6CUEnEHoGdHyGRSiL6dCV
XRPtU9wDIddAefVMN2HEXd58caCy8OXGGbgCQfvwoy+ZQ1flwkBO7PVzAj+OV6dVC3vVXRdt9q6q
PYMZgO1AfKS+WdK9OreIr0wqtB8VPvJT0sRj6ca+SLeTqzbsta/ICiaDJtJ9GSc2oFM2kKWD2dmP
VjszRbM1wubJC56MU0+bP9baTfCRPa2d3JndsHQPJAzeMRyjay5zAvpT7xHJyRQtMm1tbaN5scH8
a7yQ1MKRtBZ7565XOSPMjZvxVnZ6ICpp9hL03yu7zUdglVrFmWexGXOjU0Emr7FpCp7A+UB+hQMe
Hkeq+DRRdeML3+D8T2fucgKxf5GbktdVrXHofuBmgdwI4oFfdicWvGF4WKX+rX1CnEYrvcSdl+nE
CYYvQPc1V439fekxhU7GhigmxOkd9crmVwq7FOnFFbNsgJ7jLtipIY1LXDlZ8bets6NcSXEOvISF
883a2x2RIIIqYhgCQ21C/zTbu0TeExYRMRi8HkjUA1Jyb8d3tb+3YUHdi58LMDiG9r1iDKffkX+l
cTxGjN1nlC+1VElBLfWUOqc4KzF8HfRHm3Tb9q03amj6D1LkcZpvIOENAYMsInNDfkXzHE0NmVDU
7h8rpEfO3l88adcbCj3COsSG+8wyPbcJwPxbgvGKPR1JWzvAawJ8mb33ulyZfJ9HD2jQiodrn2Bi
hZfWLxxkh0PPnQ2XuzTDw6TOxxzOraIN+Bw0yBh7E1OhKPhWSODUrGXeB0sLdNhdiiHEDNxJWBsH
8Ae0YgG80CC87EufUN8d0MNjLIcU5bJeD8bc21GDItj3VhagKh491KCzJSFsOIFFGKf7bZqcpavI
VoQ9RHzAJlPgfSnixVyOetkW6vw3IIu3tEZpDoSflyoNDgcyaNYAL/MYZ0luT406DyoZCMi17hqT
dlUX5iKXtNVTGfiBs2evpTJWlbCQwQTdYEsMsBwRz7hHG0s6D9Dc7LQkVbtFNAsTTNrKNC0kQrcO
0ggdOPsZu6wOdqhWdcn1zaLnGdQrxL1A3hUyJJ7QZmYdfDcev+ms+7WE9ZWbICzYmiq3NJ3d+wse
2CgPUGfix4svpBobFb8Vdy053/8niEo6N0IWBx/Vy7i62E7li7AMiZmN+Z+9X8HXYXgSo2BGEU4u
Uh92bOovsAwTLUL99EaOs4mDldAQ094OmBTx8gSSrKEswLyrLeP8ThMN7wwzewJOVrv5cZxnOMv7
BzRWE5aQsGMU/gCiCaqnRE6/S8+s377KJ+t6r0UUxtg9DAbyZqxaNu5/7jzJ6Qw+qknnr0432nnB
oQ82i4mhqBSAEcbwPuXxs47uLeg7fBjBter9YQJ7ZNO3SAauZERGtPtrVHowK/zX+6xeN8ARJfTH
YhLb8pMCS5x61c/gXer6dXy5w2n7C6KRYLXc89uftohYHaZe67QzpQpO73FHwG2waELCpoSvelR0
UF/tdAJRFZDzmVIbVRxZ/RViqFYSLqXPnW87k6NVdcizf1mQFY+xeERRhlmMykPMkLTa6aO5y7l2
iGBkaScuvvswqeJXF96wATaezgVfaM++2IsP9rX1LqXWA5cNFyZD/pRocZQELfzZpcKIXaDzsbRn
YuEo01Xg/kfqeRBnXAiQ5mvoqpyMWImUVNXl32vAMzn+cFzitZX/N/yhCGcL6afgS6ccfxX5pwV0
0/fIj++vDSpjcRqYNtEkQvF12FNKNb2JKKoU859Sr3w9U42nPo5XnWdKN9GOjyBzeO6v/loxpItq
xmVZJqhhAMQB0Oz691L2bsh9KP+tpQdJLuaMdhiAWRSGYu3PTjyPJOe1ExjuZYAAFTtCjjeeJ2yR
nsch5Onp74TTQNQ9+JZ8roDE6tzMjiQ8kVgem1QllKW9ui0gI8zh0PDHGHn2D1GJdJ4a9qjB/QRH
y/O6npv8O2xBB2phKtvY0+3vWkJlQZMPgkxXw1jpR+5OELhcqhKlJQk37wQSDQL1jTYNN6+WwSCh
JiC945iE8GSLZjeA59oJWw4gx275FvJBon9vytxLuG66iNbeQh9CXDWf+v/UxtmLoe4AG7spEin5
4bFDSxdvajyIE3y3EKauSeyVcrazq5esBV/duO+McfVxAuYxfkoQ5bBrLn5jEf4iwCqR067uDNo2
SGTDjzchVIkjSYfG0otDEcnBqmWb4UAWbbWmVdIuK82AL2U4qzMQ75Fro60XlJAIhA/1+oKGhtJV
qEj97OYk6bFeqva0u2o2wZkATIX37olcpSwsmvv7jGPj/wIvLkkYC4RYIbu7SOMs8cvSzSTxp5JQ
WgfIfqVHBaTnZMyWAXMf0GG0/a5/gHjVLwHVqqH9Z9uDF4Yz6VNDjXo5NhjFlc4PhAOBXRza+4sP
DCq1h3Sv+tVbZ9/o/fhkbYMX/J7ituf3cDZFeKIMdgiB7o1AjXNB7f+MynugJ3z/72qNZUpdLuut
1/eVqWGYYpVjmWmlOO9AQ2GvCIqqenIHMKGMROmNR3e93bIgTCWHmlVJtCibPDpQRVV1RLp6g5Dj
WxQgLGO91pNIQiaDbWSAmKJ3Gj/P4MPoLpBm9ZhiCM1Wbp5HPoHkDRmo0eRtdmNjJSoLK99888e2
jOFwoNsXBxrxxqTnC5lvM3NUJzWG4+CzBnGsTvfbJM+2OW0zidNAItPylm5mmISnu3/JHy29PcU6
2tandzjffxdEvA3YSD3xaIQToAM65JArEakvsEz6yIfWy3WncZDKblQRuBCg0KImxMbfF6oMGtRh
kyJjwQ+4TCY5BGecAiwJ2TiwgaH0s0Y3QXvw6M67IBGGyrf6y/Ov4uKJQy29jchQmjZC/u7pLpuA
QLvkT+8ClrX2e0jl1fJbVMt8zapuGxx6QVY77y37AMyAxFLylxsBLYrSSkqtj1gKUvkZO+HtdDVT
nJ7e+H43FbCCxomtJdwE8A3yGAfI+OB5Nr6Aca5HIDfsM54Pctz3gKLC2bLfU9RctRqVDif08xjA
1O9ZhLDiRuuc7EW5SEnTnP0zDpTSW2bCxp+isnj2Fuf4TE9wZQTnIxZ/ppygeQPLjWd+8FuskZxN
rOYuQJ1Pp266pilwfyvUSgjGIP4q6Sm2uNzhTltyfUWdvGvKQPGsDe7DxzzyBIwszlwwNkBAVcGY
St4m2gv8p09xNsKdbrosyjHhoOcbjVgz6NQDef9tI+raVJOw0y9yLe7RG28lhjOyxViQiooY6An/
fNWI5fba0HRYEHerxChpqLboq5ekOexQbqAZOFT91OR3EOec8kyqw29eaUqIjfTioov3Ajrkflaj
y6rOe4NgoQOa/fbiMjvmqPVsiobb3NgSBX0pHq8Z3gpuD8keOtS1xAOsfmeRL/m/4S7TWdbogyz7
e+7E2vvY706+jPf/hrJOTgCi5v3XXwUG199SsQmNLdmrxhtA9uwpvzgGJsI5IncIAoXXB5KUKq/G
Vm/jJpiFjdDneFbo/qTU6QTG7NK7fay+4CXWrI9lene9PZSmqi/jyorpwx2/NMynKEBrOC+TS51S
KM9aLHr1ClcChDpvVahe7L3KhwhDGZ8smgpRH+WbL3hb1tqHV6KTMTBwNd0SZbij6BOWbQ1oQlPR
WZ78qrwH/Dl/xGd9KimhH0O1bn9ugA2OdFtMgEzSvqKhIdV3Mv2pXVnUkmhwVEWPgJZgFRBhn+gR
1T970L8wYMBoA/vj3w6jEX4Ib4/dit4hu4C1NNTs+LdosNXNbVj9WGHcMNDC5S4YKAPcK8nVY029
Lyl5ejQBl0vUH4qKuLB25SM21YGHxeSMZUMTCRBrTTEkLRsxpGuUeb3YfU3raSm4lregrNblb1pN
e+0jusF0sxcjeSVHic6n0gOQVee2BPqaxf8vRH2KR3bTKqtvqjyqW3pXDzBEGbF6KC1Me9v/L3EJ
F1UUDwI6EiBgPVDHniR4FMzXclCjcSF7pbzgvqOf8kZjRxq6ALholYKtAUCWMuCk8vwZ6Ji3re6m
nXhgzrW9+tzqmzH51/96ZS8fQS6Nx6eLj0HdimEcW2MAdxC7Si3Ms/ulVkKEvFK9naVF7JEBM95n
Ok31rDIKTaDQhDgpwKHfviNI66dgRKM/LB72mLE1NwmKls3LBx5aqIRiYP3o2FvnhnWBmIwyTLru
IxLqOTxuop97JbkmP+lu5mhkF+U7FtEvQm+stgtF0VuqqE8FMXBm6nY524AhQarlD78FeBaCK/Uh
lOOsy8mWeE1NZdHsG+NdoreEaTUiqdsmTPvMlnW3++LCpkCbV9YdR3+QjBYqGBtbL5D2wwWba9le
CBewhH5L5NM3ocAblvcVLIoxERJhvfNnzBw5tlXh/p4kRzQq9ILo0K7ylU5CkmFW9iTqig9TSx/+
lX6ZEt1QMshSUWaIO0PSMcTUPnt45hsnZzpJQ5UJxmt/ZWYhFGL3pamXl1K2MUuiMGFHR1u8D32D
Wa5orcirKTKaZtEb8p7zBrdo84yCnHkl+H+GRuft4pFyLJ7Mm+uG/vY1wv8dSBUri9JMimNnYAR3
7WQHxUevE0vIiJhAzZvNsoaaFd4h3DCOjtrbm4q0WSitTQsOkeaUmOYEGnsWJ8SBTNYB53mRjiHt
3N/csuSJ5EFlqmFDl06DM8KeV61stNWDn92TLo44t1t2nMM2AeRalnktnZ/ibxTaRea3FwqhyzN2
irUcZia1jCgXxh5/IoZlJaNg7SeBMYgtQ/9fC+VFVxh/GtHlW1Grv6m3KP/20TP9uMbRgC50KPgT
EouSm/wigpgfkMEta7hxRdVtPsvYYLO/pKteoY20H24l2KdlInLnoUIVlUZjjZW1sRTL3OHJlW+d
5rc1+yOOg1nSaV7YC3xbf6smtF88ougTB1+Idxh7fFM106rDg5rKjPyma/K6l1V/JknpR82cxeWO
mLV70qZj2QtGAbIngKveKd0FHc2Hb6myxia6+9XCI8xPHsQTfWsf2W0kyNhJ2+VX1+Dfi2fSFDHi
nPJqikmWkvbMqxIfP3ZE95h0EpSOj8fWistBTg1qEMvd9lX+Dm77YejnQwOikWSYrnaSyl1YlF1T
Z2pAGm83LNkOwFPBow3GZQ6gDuYFEfsHojOE/xYaU/vmumndfF7VjDwpH9rXlXbBwdWA3VcRvmXe
x2symneqYN+ynuqMh+xtDv7iTudLOhwvHpL2w1tGl70OrYVz+oqHjen3o1lv1uJP8W9bNc/PeZcV
XET3u7QAxp5u5e94kIt4uS71wTTGn+nQ9mSf5ZRndd1sPZjFnKoAmTy5FEA1TFrT4i7EpdUNRsti
q37pE8SeLjqbP87qEuksYV5fGRzmZYN3ETspH6Wvw4EKnHEWhr3EhLltRv2D9+bn8aPTPEMy8E9a
aBWGDwYofVRlPfUfomgvot0qNkl6q3TDNkGmP4TM4Odqc35l/+IFeVof2OfPnWFouVjPFYm2CXva
Eqle7z1g8AwDtwqdnad9EZgUSA8nBG0z8SaogrBC/Ql94bllkSisGDJz3/dQ4Q4l6O6CwEKXezx2
/xVHCPGBt28Xj2l3gdtF+A1ZcZ8oSlE7bq+SHZsB58P2VZj+VP16eI1K19N0LF7K2gTS86nSTo5N
4L+53PgCilkFv75XCg4O8kDth2u6N7ITYHl+DNKAR2m071nKpiranNAKRYpP9ADExgQkYfO7C/vt
sfOfeGkYhyDwjSIqO6ugFZ5ulzyPB+QcheaWOlVlIrYh6ZzJG75LmfuzG5DuTDY6JYQAvwQobUct
f1A8WqdCwku5M2gCCCcVkhfAXQRQ5R4ygwFQj0FaD3WTbU6daprE5zV404u/RHxGdA7jw0kXpt0H
cCbTGZrvmO6ueJhAXVV9wzvQMmeJMIBRcwP/EpD6hLrW39QOoQmFmsDW1DttAr4Z8wF3d+GpFyf+
RdW9X1cHEo69DWqbkm4+8lMuSd/Ms8dSTyY3obFvegAm0kfLu2Fr00GpK82Pi4tXeGqkGvcSE5xo
BiL/CrtEvlCRyNJRv3/bLN3kemcKdodU1NiMwkpA2y6jNhBWR843Ew5kB1NlqhHFvISAsFVHtHQ2
m4GcLAuZ9DNISv+awAz4gcf9oSJFdfufPKrcoYwEcUsfu3oVWMmqRGjXq4+HwV//M5bPc7ybpiej
orQj4w/r+tkF1cjHXq3imkxeujGeZ2q7HXvyPAFkzv5RFKDtb7gh6G9ffs1gwSmlKmupGcC0xYUA
PYH6Dbo2h86XEe4pV417LAsFgAM6GSH6xqKpb8puhZ7hksiMzksqGR6+/vZcIkxLBOpWOVYpnc2I
2T7PK/zYwS7nuCEJMdc8gRUIciWJQdN32f80A04GFj2V5t+d+VfC80CJbeg2hIzHWgekDKCk5QpB
VFsuu5ThYXkMU+vUT1NcoJ5m4OLGkuY/7NyH49d390sOWufweygOJWMCI104/yj/WaC99F9101K7
to8qBc+lcxztFaltAMpKzkZswLcyN+oVeOusu0eE27tKQrM9EknzW3jPmLe9uPXP5HtzDHFMsjwd
yOki3E/rnvQjKQ5HW/Rl87th8t0057ddthe4VskhO9vdgJ4YLmoxGgotNk2uLMNG8e+JsCkaL0/D
W/tCfUp4VDsJcoRLFF7NljB+iyJ0wy23xGE+gS00lKs9AFs/CGq6oSO6lSxe+v0jrLA7quCO7vao
0fBJ/iVpLhzoZERfsrsX/A9krZpbqrqiE0SZbfAjCaIDKqAD9N1uEMTMjuKTbaTZ32w+92Qy2xux
3lsWbgXgapvU51IhRo1ZNqy32OscCebleNlYmTFPMgzJZwAoCs9hJ0a4cFsI393tZ2x9pVi2TpC3
vv2ZgERcIejU2yLXc7zcBVKuBozWNOozidKZghzFjTLa0PiJPmF7u7CxOOpaUZAp5ueQ51gKMxuo
M9nY5BmUqf7nXhAw812YTitsbCJsIfAfj+U15mDaRX7mkCWcfN6YMlUwPKmLrX2Kx/FPhcJavuym
Zfs9Iunnmp5OdmRZoITF42OCeBYpHm5flG/oJkzzHQZcj9WSBDxcRNXAQAupi5AwYKtREL0j+LJu
cyL+E56h3rxozqn2I66yZoDrl3JLjaOLyUZDKNBY9hks8kC/0JwglpisDFQzrenyfH8hk2orc4Dd
1wXJ86uWXR0ECInpxsK01X+b6WOSwMKdTN9PPcelaF2EsJ57CMSZq8x8S8iUKQ9zG5aOlubkPB5g
rEDEmKp2ofQusEJleUYrkykjau8iD1v9n+ZW5ec4v17l171eBFfMES7QUYmYBavQXovnWTR0k+Kw
uV1X6aJpX2Bc4lPUn1RdU69NIjgKG1gj1KYf3O3SP13GD1VJ1RYWbjCTNCjn7zAgBo19O618EFxE
85vxx6KZC4jMIcWYqBZ5h3xNza8XETRB7LfXpWUr8ACY7W4pAzUs5wy+AcAn4YwiVhOLMULkjcTw
oHXwEWKeVLddzM/4/wcgMSIfSuOaMcdxiIEQooMZwiSK4pbosZZkmBTmFnTUKC7RTH3+S7NzFQB5
gp7W0hKjkyzY1x4/s6iKDXK6OnmFBQoFkw3jb3UDNAx35NFmd3i2PQamcvcE2PhDTxb/cANiE3mr
M3yJZ+q7GZFgjXu89R/hgVMLW5jeJOKiW+fMoZ4zfLhL3OHovXhHoX06ek1p9992kL7F04pJlcuc
rKvW28EfagN758k2rapetGIMceuc/iHe/2oRiIKOhVvnAwNwq4JJNz3Doe4Y2Xi+iFAKEjXLj7lj
T4FJVf+aShhWEO89+8aQ5EqggjJN4OdnF3wUcTNqlk4c9zyVzBfFAW3fwT5HYwxW912ZjN8c7GVy
Go0gyRS8DR1O5IccNCkhYGF9qNONU7s1moH7jBlXFVqEPCL0cmwVSmaQQzaCgJ9h59VF2pmuoMv4
IM3wMq6CmZajAee7c2Lo+1992S/K5eoxF4/R2JIgQX6bmu+0hRA6wmLxzdlAV8bqzTOvVO41VNt3
hk4R7aB78RWe76SofHY9vGH8RE0i4TFwW1oM6czit+Jav3mHGYKrCn/iSX+FXIDw42wguWxURAny
yxW0cyxlxySCQzmlub5AvlkKmNoLYwzP2xZcGBsL1AC0mG8lrF2W/ti/fuBrG5UX46FAXGUzhM87
hmQj9DJX5BrQ1KHEaLbMGTMn9xea51pitY0fAaGBJXiOMKgzvwOGGVAC2XjM7oEXm3KnV8WdvUpY
C6yoxrC1wE6pQT3UUmg8VNKmZONFJo4wLHla3VRTufaOARtphm80C5bCTy8Ilyiu90PnHDdgulCK
pZYlwUY4ykJG8mZTGmfLeXdhbaxH0m/ujvJUbX+f6yHBbmbZhOMtSXchpJsc0Q1xlXRkDxRiESE7
qsZ9MDGfijaE9jJJqP4G1xoEEY/+qBMqUfee5tMUynTIW7IJLTLF8NasgYtCoRZUXX8M7gkgEq3o
qm/zt/mUbIELrLwDhKzWkJBwXI5hCJ3H+mqPhubWiYQ0dVMMconGpSf94Bm9b9DFAEMgNU5h3bjZ
POLs2aNUnNRHnX11W6896V/K6IRRCdzVfwC0TS7Siep7b/NrySOKLn+4oEyb36puU73BDm7LHvRH
4qFp161RSaPE2bYSMlksjV1ALIdhK8MyAgZmdw623wYqtC0TIbAQsokmc/+wiJQPkuzEwiW/XIhE
hqxV+aXeCdR0aWhBSzXhPOleCE1yigM79TVQxFjWNkPuJbGkQZqbKdlU13IDMs0Kz9FSLdud9Lu3
BnMWlYgYFvUYKZw98PdwfAEGPets+ljsJzLYuWdPRyIL4kSZGMzBm5o4k6CfFd5C1FnDC6LHqhCf
OD4MGISL9wuvlpx6vL+0E7YuoLMsgoT7EWFKUcUyu0G11f+agCCxtOaz5tHvJUYwxZqjX3zbbVmJ
vZdFm6niyYKDVgwAXo+ceDEBOBJpxZNCVyQSgB5+8Hc5h7Lgep41TkHNHWe54g+gstPr7Un5OfTW
GOrRtDnCPA+QcNZLLXwIw7YLDm5WGvlnVoqAGaecq5ejb1fiuLvVAAkkqKxtDhBl/c27wnYelYXa
QxMRQelxBbeQ4aq4/MLngjxK9WtqJWiG76856zq7WKHo+BUeWXxOYJarq7iG40+lHmWOXwWbHEBa
sJ8c+7B1clwehHZ8HMfvV1bVg2+S6CjqJT/bjILj99438yl2Z9SICg0FSV0PJO6ZASE5gQmmQ0b/
uSYwyuO9Ab65kz9jtRPN/+tG/gmZg6zIEBvIwCNakz5d9xYPgaDOtsYW2Uuj80GmgVjyPPin3a/4
MB1rDIsIQzJxyGGyQO3zKyVaSJVcge0017roBZ2qUu9b8v0IRA1ryNhWzBB19ZpEVLQXvSCshJS8
V+P+Thd8OjQid+kLcoEZh0P7tsIGXgL7bI4DXhZa0WH3xJx/WNleIOaVaJRoexc31QF1Hkmk/2v+
qptyF+2ZOCG7+8zaZ+PnA4gcnj/9sI73HpGnefjF0yYzt3PY3O43tnb34V3IKep7ln/E2MKUpiJd
qZGNb/82Oe597zhK7ibJ9RsWVHcxK6cNFUxhvTMPLdcZ5TNPFy/u7Co+vpMhGC/Qpe5t2Zt34Pgz
yYKowEE51QYNybSyhib/OsRVuX+vpVIrNDoZL0MDDkIeav+txgXpkRjeL1IrSyjBQJSZ828pViVI
ua2sk2Zt5Cd6JsLv4SX691OlNuJbXaCaAxr9l35rQCc7UGjLfnjngisknMPqBv6GVAbFFz3ha5fD
dn8KUBOnayQlzLjp3/HVS603139EHSVmEJeU+BcKMkyg9cXIcD65qngHamStFADm0/bwiGzNM2Dh
/KRupPafN7F760ZX/04lQGJpvyl5t1q99x8CjP/MdiFbZUD0iLcRpUPW7aBmRyLamWrRniQIHRqk
FSLlAf6QXUGHJ7DP+UTc8CH809gqKlarCLHQ2Bc0b6N67yHn37NN/WR7DV6qkRThCmKXd47mV3CF
b0tkIpZW19grz0t6pv2WsBXqz57SBPCp6n3UAnbclDYfxq2d0E+fEofiu+WWLs2b48jbKaI9OYf1
uf43sEyO/mOs/oBBASGUFvp2GgjH2FY0E4ZS24LMFUpfgf4osTc38MIAm8iEByWWXiXtKPQSyUhs
cTYg1doUEFtBW7uM4r7c7tWbQrm2tmJfmyOZFFJEQxr9VLAtdLbZDbVok6RJymTrxx9BNX+BXCaV
gBhF8vM09mjJAsZdQdmclV9dWUhewwk8UarcEvCCX2c7bVw8jTqiwvsWh3iqRd1mHvellDDccwHs
xkuo1ULzyJwGuv8ft916yDPZq/V7avwcjFdycG95DgOBZrqEfDGPU7ZcALk3FYfln1UTRdWLfrpW
jvFfWFZcpZZGFLxai8wyM3wOGjgzkIH9EhVn90KyoOP61yfZVQdQFDCnYWxB/QVhbmr50XDGFHFO
5dGeu+l7v/gzoF2lhWMnakR8p6/MSxeIQje0xwJMe50HFwHANts+vx8Aaq0GKqda22MsefPSa0QA
NnxZIE33dA+wjT8LTISOYbf4c+Y7YMNKxISq0toSbIJ+BVz9rfr13BYTapQY2yHm8NXAKdFJabii
2xn2PX/s8H38+M/B47Ab/MclA5uJZax4qRRqWyU4FZs0DBVkqszIs6k+q+jNc760RlUTS4owbvlN
2Yy+N49lDS6AclVuQ4D+nBxDOHeen3qDJcBNR0xLV2Myaq3/1KHoOtNDWRwGOZT8E+/+Zg6czk/o
BS94/iK8EovCmit3yegs4s7RiMYNN9YeglrQGkVuH+/Ge3VVzFI20toaFuyH0rZ8PHjXmB+FeNjz
CnYQ94jFI5SsxjCVCKhMDQo8e051EFfsA5yVTwkE8HTZ7mklLDynLaeJYtw1mKCSRwf31BJPxjco
0bPXrVbq5/YN57Mlsj4JpoOFYpNcH9bbxZKaI5LXN9QK+/4HyR1FveGeENorcOnPMKy9Ku2c4MI3
dJW6uWeY0cXvxfF2eiE8h0n/Bjw7tm5t3Fu7q/hDbLT/anFITcp21jlMnVOpUFxodap8NIOHWKFu
P/MOfx3vb50hYu8bqueP8a9oPspfVug5KA7LMRljsibNwBE/kWFXdXH8Z9npnxpRUSo3ecLbWOrx
j7zCSerOFWsg5HK8eDmbUuM8qzFD/kdPTaFvH5nOw257BFmaluiEFdBz+C7vwhpbTLE0147NhHNl
PY0WCnoLZZtaqchWYjVP0R2+/b2UaVrsXbtYyxq4itssFst5+/cECdEsxXlBUbQVBKOzRT684UBj
U5eq8L8LutwT6gm3U34+e7WoF2R1HyhIF4+7pjgnpwKhzaLoeMtWxHpPiWtZW70HK1/h0oK/OyEk
I7k5AOMywKDt6pGvJKdlv3zhwuYkHaKBrd8MM2rWhgXQg6u2ni79sYXGBe9mHCOagaSpmG3RZRx0
qY2Hy+HXNvD8fRIMv2RYy4JJnPmrAAwpHx68cNUYaB1G5J27BiywZu7gw46uZTsU261xl6Dq2E7l
U23eFtVd4EjAvrPeqIrp/oczGSVRWYrNSEtThReX8/1KkM3v1TueGk8wK8S3f5ZimwzWgZpHRLXl
Zln41Ga8GS788Sapfl0LSHYGvHbkGlH8mtwCu4MMCongFRzlc/dCwS4wB+pPvrfudjgaIfUTR2qS
GTJsyH+lp3T7I9U62SpnQULksVsjn2UcFn137L8lfVBEfnk8zgO7qcW9Srx6LXoSLdi4kYTfIjz1
a8mmaloihP3+u5T3wKqIfKDsdBTEemwG/uMZ5bkOmaY7BbWZDH/9FFB0ESoWbuBBl2rtuoPp1mP9
ZHFnanfLOKI5q93H9jv8ctXedbzw9KKqW5kDEb/p/LUOB0ENEpRas4epZc0ThRhkcJSSe3sozn7i
w7IriM0mA3Dj2CU3qwyUXwvqSJHpXE/e9mrD6ub5pd83RguHVBvrThMpBBjX8ySs3+qQshayqKLh
g5PB9eNzc7wvJOusoeI4txgEWzvVj83oIPhgfzPqYIMMpti3KpW3If1xNDThKQHQtpAiQcK/d5bp
kgF0IFuhWSmIUpP4gXX9BLjVKn5qv0r+4YlB9kaHBML8y3NI+tNwiysDndXdHVMlHZyVodfHyc/g
4Eztei3NDB5niRssVV7K1yTLkwMZm33esVPhG8tceLITmyqbwfYb0zuPVICzIsnR34UqHxGREn+E
ChMr4TaqCSsFvYGdu+5LcaiK6slP4itG+ah/sA8oQzuiKhC0+NlbFxxBPWFX7y6gDLy4TBS7d+iB
lDVuhelvEP4QG/ki3H87y22FYHJYMf8ymPR+njTk4R/6h0++qRWMJM2FKUMTzhqvIMdv/4vv1CS2
KZZyJ1h1hekhrwlBRB4LCz+lTBnz2hHTgC+drqPA5nlx42XfsR+CB53J1z5/PWNe0BXqlJGUmV3K
Ms6mfLuMr3pH8YBFmlUirDb+uF3HrBltO4mizC+sZgHAU0u1Pol4oo9BPpcjgkR4BRVloC6jy4DK
jZ6cSjGh/WiCMqkGrLvt9cOOwlwfDYefIF9k0GRlRe7lVgvhXt7JddUiVIg7xfcE3/Emus5p1Crb
QosJubR8zkbSgKtoyR/F/3v3ne9dh78esVtJXpk0Y6et694sD23gXtoKxCWw+z9YgSlA8h1d8Jmf
LeJsTUSv0EGWK+Pssz2H64iKKdQYFJFdXbHIytv6LEpscj2wtfvwU6Y3xa58QuCePeDhSeIAkhfT
cKvcrCCwtDOqKM7A5jU9yoPov+3oF0eNkTw6zFLWoAFBIUFtJVYY/ZXoIP+Jd13YhzwTs+dNttUA
WaWuzr7W6CMF5hOGOvAHBvI1FO8srQikneHiq6naRaYcQ5STz0ycl2K+ed34unrp8bSCgSDvaB9y
8w9r+beuTPO9/zqnJTxPjGD7hd13PYKg//ubQty9NvTx4YPUPfx6a0TauRxyaL+L0qzydq0oTbaU
VD6/iYJTlQ/93SG0EYZ3DhQJzsQPiAzTGo706n7jctdk8m4nol4hWoGzlfrHRzUqG+Nv9UAudNg7
7vcoJxoffHeZcoY+unV8TRjb+XMODYFvlDlOjS1yhUTFeVmt8yWn0m2zmDNRiOWs1T0hhcZhncqq
DlSpn1sTFZvkxE2AOGBY1tiFGs3tJWDprO1J43ehG/lhsWpdoBlqc0pDV84g2pKBCBlnPHvDSO6S
dRcPl1fD0uWxUOvLgts0HLqjl2omSAsA+fpEHp4xtxabW182smV6PNAS6RPwBW+zQChZkskcOnSp
pCUp7nxIa1wlB4iwqSS+haKlWo0HXKgjLl9HpgZi6r5E3MOBPIPSer7KF54NfOgW+3Is28vDSSoc
QfwvhFPfqeZ5GBhLD6eVIYLKy//+iuAtD549qNiZJsC2HRyUGy0p4f+NCwW70HO7EBByU8DSfPd2
+t2IJi0zDYj4n1G8Ewvdgib3WF43RkS6guHowD1XkbLhTxy6BAFAhndozlTI1mEbryIepEe5nyfk
OWTkXLH9ZOAlGXzZbBCd/ZMd0ngBMzbXQLzVF5dNTHwMnx9ppkYlNum3ljszEqOsCfklJvF5JXiz
gWz25+zNdAFY7m2nzpvwnk5e9kUfYe0WRNIUZ4/wci9LFyV5/fOFUt2PYRq3fuZncjeyvLDmOmWf
5/ja4AN8nn7kx4xK141Ii5HVyJfR7wozhxL37mBONHk3L6/6PbDkwM93wzRWDU6W/oqnmQpOZ8TG
Zuc0LB4ToBAtFs/lqUVnlfwHZKQxJMUP2lirrnGOg++ul2dj0iWX35/GHy616waXJe5bvMqKLoa+
feBDwKVeLncUMLhjySMEW3hSSewGzLgOhEPYD+7UW3sqVQ5ETAkxjlJro8ptbv/RMl8G48NTMFlZ
6keTBxS3pVyfmxKkt4sVlfRCmDhJ+r9Gwi6qz3PZg7Ol5tJU116wc9l0zbtDVLJp1XyDhmGXD0YQ
qPRcse6gFodF4QyzxnlBtOtAg5o2bAe1RjZyF6QfJj1YOTPAyiFqSvlDR5Ewg09h/KDvS99tH6So
qQLYbGmpi4K4oLhsFb1H4LLPC3i2wZCy7qGD+pNv6Wseaw+mdgEoXAnjjazlLK5Wco/A4sbEK7VR
594Pn0voONL+CHyfqu/mhQviTjlxUvTJu58H+N2H7nY6Vj8W581XZ10ouiTnsw/o40IAN0vsJCKF
P1lnmff1xGiGkQa+MbEMAzo/VJ49yIkKT+ac0wDcuR5A2mo1MyBvZ2VALZJMtak7Sp+krMSjK4gF
FPILm7Q5f5ajwuV7jW7eEu0ta5uwzdXHlY13x9jVRZJR4bfDyUc5vBX7E9WVPRXYaXjZxbO+g8Gg
6WsxoBtMhxTKHUUqkR2ydB4RBfBb3NsIt5Z0IaMD9XZtFMGw7BhfwLRiOq6ADNyPxRTjEZzZA1TD
fMUK3WUOjFjyUvg9HcL8LWrWgpkFQL9fho2RWKFQe51gNW3+nNzrEaWSZoVbb/e0AW9aKrc3kNQb
6ofJI3ifT06buq8mU3UksME2AsT2sDnsJWGvyvrY92cl62GQM/0nR5CXDGwq3hSDX+E7WFYMxRz3
NFvsyLDClzQM0kyLDxpJFzShGfjz3Uy5q7QxZenaXwNplLtsfAYPW1xqZSjK/tt+kysZ0c4tGZLI
MrtdAaQT+K8vSRFKd9TCkokTh2XYUpQmhJHurl2+7gbjggeywTGJMiQXRxDxFuyFhSHN5vXvIEhG
Jll5SBGbMRWNBvRMovt7pqa+OwFpEgX7cjmr2sMVkcJ0SaqWYCJ1JpHs+R06hXjQ+CXjs0sMH+Ty
ojxHdSUa8tHBjs2wVRh41WfM2+NxOGJI2Vbrx5i6L/nBenqLEfYX7hYBT8G9YxBdEpAiWGxitI51
3fpgHq+YrNoM3N+dZar0IwJUCTKuw6DloD62Gf8WsjBh7s52tN27PqdeW4wWImRUaD7VsNeAfyWZ
VY6dZVlb/EvGggfJtK9y6sbWZ231U9Pomg/c/1oCgrG4eYCM457dMgnkqjbZSF/mXNOh0iDwFTDc
eXyivka0TdGt4XiDcZ2QmQnJYtVHWdVaL3/jsXouGBFVYJVw8y+Jl7o58OdBkLkLcU7OhiIH6GHb
eTbSlNdaIepf2sMfKDgHiCBWaSBKMrltsWeNH9toJR2z7J/Mkrj/jncxUE7TsDz3GylqDI2SGZmM
z55/uI06n90aMnNSt8RRYXMI9rixoKjgt+SiPUWsK65i6k0XMPClwRlxSNtxSyzT9cx4+Z03wD8Y
GXKyEjOVdRyHprmLuh4/g78BCJO2XptlCU608SKaZTYSFsFK69DPXzAH3NGQ031tEwttImqCJSXt
FnWonQLilCAPGNWToXA5+xnVfajqKZ0fzv7O9b0+DoHavuEDObycJ7DFPr6zcSgwng7OJMVkhmAk
5KfE5hhdQhmIKyEKa52lDry3qJSQMMH0bu2vqQXN58ta37Z6XapMe0UYmyjIk6Kcwiz9bO17qgPK
fV/iX29e93FL4kJbBrBm3bLHb5Rq5tzsyRMYiaEpHs81o0DCj7HkvDNemrjykbu85UEc6oBEGZks
loU7127cM7ufJSgZfW+agwrN053leT9XlkkGzBqLY6C4R46iUvg5iUuAG42O2KD2SWh8nusNT1f0
9WTpcvcle8NdxAggDaQNNYZIVT2zLDs9qPr5IbLRcNPZgTCSv5Ly+DCdhkUiBrqWzWETohHm65qy
3xHsYUWcGcHxaRCO6+GOFB4/LYvST9Zghnm/Q/0DuukfO85C13Y8eU0xNF+tmlyWdB1BQtSYq/pd
AQ20HbVpoZYQK9XC8W69b3/v6GI/9ZE45c6cmWd2/GW2Me9sjGzdPxIqUBqHk5/rAMIH7NG4zGR0
Z2v8xp6IWeCspqvcsir/wfKk4vDrP7lt7nMrXGhut+ioRbQq6WtBhRBtoe5AZk0GqSb452ehtF6P
2tkF2ZpOFvZ9sSe8SMg2CTaZgJQIhFRpXTgAy3xAZ5fYXcuG2t1D6cndZSsHooBoMBPkrnrbp0GE
f8PtecwprXqnckts2Zwor3rW5OFtp/nK1U43NEejby8KOgFjfJnuhC0dawPvShdR11L8x5Qn+g8d
a4fGxsQ9UkptVfCqhn2DQM8s6vccfHZohr0J0YGP+IsYpyoZfMLogJSU0W72fewPPwJDbAQXcruL
n/WWmhrvhzZ7BIOTaMEm3KsTG93vwBUcWoPTMzmdQ5sj17hleyPhOoVvyD0IH2kU3DsxFECTImha
Qmy8N8mBEQKxHtGd37vuGgnYiYmbZrdSlkbaa28rYSEqU44wqQr+R/J3AAcZvQX66BNd5OGfUd1P
E/w2PyoVQrIUDsNT9+TtsS4dAXoApw62jP4ANsDqDh40f+phY4/R7CsCcmRhcpVypcywlNiISOoS
k8lGOwpyDdgvE5nCAgxpSpP6taQWm+6cUzQDJEPB+Oo94HdXnhphnRNEeEu/oPVHjonxV4Aw1FKu
ZIa5793KnQcMG8KMwI+hqmdsQvMIc/jZI3iJz4Gd8XQAZW2WtjtIiCL661s3e2tIP0cQBJWL1hPW
o3KCvSPiVo8Viv9yevStqYXSdiwMQuixRy6L3WgPMa2MtsTKhcTTjkUFGvYzWy9hi3SCVGNNZ+Ru
dpN3K6WBhJUU4+6jN+IaJUwhYP/MTRSk/gweJ45lXMW42IafquPtc+b/WAsdB2Hbjb+pBXekAikC
n1BpABlxrlYsnCiS/dnNC9S4o32/k3nrdCxghY0FyPCmxpKRSu/pXsDPcch2kdaNq1JwMdkOebgy
H1lyaTJ6hluQIYTOZDdjSqx934w+QmvKyP/zntNaZGSNQcnuvyVks9/Cg5LpZSuFqUgwizHy2yX5
8Afwoijx8XUFrHeEapHLSSg6VHFwcOqjmogVmHwrPUQ3KTUsqjSloopUf2nio7iRPUrhttrFrEXK
yY47t88FfBUaLm23nDfLxM+6uWMXjzmcrBoL9G6KoBcuiPMTo/5CUyU+o63vjNCg1+Q7Bms9BmhK
+LRGZHmvGcxScHyhCXdgEqeDLHe5SitDeMORwwKtIioiI5BSwLe3g9KR3DY+pfQHRi5SzJh+NBAT
62GhsV5MubeBm90ueLkbuPadZy7RLpexWvCytcnUKWWU82CE4BYgB5VYstooy30y/CkVNRKwN8IM
VoDteoT9BdBnwaOTHaaBFCDMpK/qS68GmHTRpbsYXfkA4j+RMWrua4Rrzbjon+bolDluE5xzq7f3
MYArQ0ctTcDGmDNQXn4QBTU6Y1AQkQCSyKVezoEXLvsyfRSLrS8YzshTfUrCrWJ+IEENhSXfa7+U
/UvGFxXZgK4qbBVwrm5gsz2TkxWYnn3MhUqBAi8jcyP3faRvyoBZE06DzK6o1uLnOUnWVcDFJ+MC
Ua30wLXJuBbIvZuigyYpVhHNGvSwjEp5bcrc7bSlBpIZShWNTGEW1pw9N6W1NAEPXYEUZI5X73eV
LnSpJbIl1FTt1ze+bmLXMwAGyB763Oji80PbCvWAy7D2uaXRUXhn8N9wwmrackxAUwxxXRoapzOy
8hm7yu9wagQLK3y52vre2lrX1GKVgsxoGHu9imq+paZv3/R+euJHPmXNiOUooCvGI8FA2hbHOSQF
QVDg9qHSbZrQHbhfqwFcMmTUHyxjQ/p8WgvnhoOvEKyq5r87xOllGkoVP+zpT/HnPZ4ny0OiL+0D
+glPYCya8TiPj2jqAECnmBjNuiuEekDq0UoK203IktnRUFOdAmJzqsHkhVW1u0RFFnVG5gpsWMFv
K8i6G/U1kjYDk0OdUrF6p39CtBJBzNMi/z2VB9RF9OqZq+hRxlEGjxxg0dzgOl9CJzpO6RSg2nFj
NFnUJpBA2HclmU3GAJX/IZTrj1QpKIr5g56vgQwdgijvJRAWiCUypZcxGwh0ztd2jtYrOQlIT6KV
REtrrul06Sm6apE3QicAYmfhOVpru6R7hTMWPnZBu3b3Vb7dVOLyMI2SaJU/oPBNIWBNiTWz0nrR
UsDd4f7B8855PFB1JFQ0YLgGQsBbg7yZYoKWBxxcMTF9a+tflSKGm13qoGCIp138omwEr1Ft+s9y
M//rIv/yf1reF/4enqav5cb+OsWhYlTnXdlXyZD4jVIXOz9XDbcRk2PteUQHWwmMstiKktxnUzFW
23sa1OpXFuEJZN475R1fb/5hT6Nn0tGGIQ4unR396uk1Qc5lL1vXNaU2oOvBp9MMZaZblTngyBxz
MVSYucyWOH3ViOiTw/AT3gV6EX6pbJ46uofBfv3J8/C4GyLFMhyDKIWqoYtAn4Bb8OaOxzwoDPMu
aVGXcrIgZ/IfEaEP7wqtfh6FfxSB6IDQBa1DGauIZOlQIIuUOTc1HzOdJy+OWVgyeTlvsSErfzJr
bKf4d9tI00Y3AKczWTMdvsAMSyBBIoYsQvZc3vb6DZXpuN4+ghGWz0xIFOMst4lRY1BmZhJD2oVR
kRzquN1MWPGZdXwqLjnv38sIStMsibQGChd6ArtcujPC5bZEEOyMB88oBkQQULlQ+1c7HvkyK2yZ
Krg71+uUeXrBNTufJr4E9tadiWOfN9dYPKcov8GphlXSlnNMKqlCkATFtp1ZPVyRECMbfkj/W5j2
qoj1H44GWk7EO0iNzWWy9XQ25MCx4l4XyaCq3KPX0lXE/GLZW+geCjvQR3bb8fkKQecXKxSnvYcB
xVuru+nb6N9m7sfwq1YJfBQCGrstlwK6vdbEfB5uMLxfC8pA5+q8RHXeqCd6Wuh2VUXuBjTFwgTu
vh4+5Sdjw9o702vaOX0d3DFG8E9XblLQZh4iMN7Vh8djAinW0AqucaEK+UFpU8tfOEpSVL9vMc2g
/ApPKQohx5YCNWBSUm39Fn2zn0kIgYUGaXtfQKITK1GuNUpWYsXg8Cn3Y0PPIAsVMa2HI3jMySCk
DdGALx4KCziZrthQmDmOaYobA0tznjoblIvRW4jsvnCTS3j1CHO9MY1U72kSPMw3ZQn49C0MZvxy
TfC6myTsn60i+GprhRx/3XHl37FaRf6VbG9ekgC1QZNCc7uOtwJtH62lA2988o0gljNnSPCqjS8G
X/OGVQpRCbnd5nVxe2U7lM3qubpccjwHSUcn2+KBTxcxETIICZ+vMOlAjEoxsKhO3sHoKl6nMaS8
bWGTBYVbX4Gk7yUe/CkvGozYCJ6CFZpGp55SpQtl1WnMfO1TOrVKsfiogqM2Ay9QmgrKqnopLjOU
oolTumZYEPy/+QAODJDwatAPl7KhZaSpcTWVk/FokgzBrkr87JboMrV5KMFHoXm2Ep+S+lG5NlIk
ItBFgcwfI3kvmRBZ1EmbrEvE1jyF2Cu1PToWVQyMOM0tYLRnQ3lGSd+9kOaBc8455dqx3LpesLfV
Mw+voOegXzVDU8cKyNK5H3E/sLzEHpPJGbD6d4G7yVQG4lM4wQhfAPA9jVM1JeWFWiT7BS8JB0PS
pMSAw2lLDYQRFQFXK7x9T1mLxPGit7MSeKkn0ZcWLjCnpn1exMyK8qsVmKQZtsu6/Wv1bztf82pZ
AikyhLzQH6KVw3n57EY/X3dSEi4IEKQS2xxU5XtxEU8J/cL9hEHdO/OvUwfsIVKXuNhpF6Qchwe+
W+q+Lq2Jwtr2aZ50wPibU5WmC7T8bxh5J7Vx1Nd0q4YNHqaoCRrbg9mdF6kGY9zthbubou+jgTOB
AmSg5AJoPff3SqoYtXbGF/G2DlGiEc51U/a9ZfLj0/Dh83pSS+FBhhFXvx7a7mvpksKQUR/sS4Ef
bBshv27q99Y932/xJ3x/Jyj9eJFnfVrhu0trt6MGX6HPzfLv9m5iBP0tkjbQzySghIOnAePwS5Pd
W9gy/QOeWWKrPCTXp3OAYLF+0nLyeeJdQ1WKIWZjlt6PwzarvCazpOV2QGQQ88F6dw7ekHXv95Jt
sbuURCAZYr3BxYOK4ei7pbjf5sw9UbNTxh3j+sSQvmln82qSeP3w3LygnynVutFZE14FIuDcKAMc
9WPzU96/kY41JP6BRDBQh8vr2r4yXThRa552JZbxqRy1L9Hu5q/uMSugmfo5rizl/+mftki+PuZG
TvEKgWpkQiMymq9lDHnMg8KoT5k2DpTza3MbF9d1XyTxf6gNgcrQSvFuqk4f4NsJyONYX47lZ3vf
B3D+QzsSurRzyutNLnqOpwCcsFOnyskwPN8gj/q4Sx6+anYbAyKHzPxSzY9v96VJ4tPI5RO19mIz
6ukWaPd6EETdXTOZSDlidHb9zjRMbub58XMD54zLxqKivU0KZecKO9HCNOV73qu/W+tmuuNl8OsJ
4KigtvhFUylZBUh+/0aJqdeQgVSfajFKZX7lDUHFIZS0PrE+l1UqlxxAU52tbQmOrGuITnJwNkIl
UfHLQF64GW+4O6qKJ8imhHRtn1tvE04Wzhom8GNMsTyQdiWLu3nqZqfF1VwQuEzrFNLf3ZnGTR5a
w5xyOA1HnFJnFn9BsD6oY4DzE2hZ1y0by0G4GqZJG9l9Y3Ly4khxDu088qsEmXVITAa2g1n/OZcS
JgcwUGpb2XMTjFFo+v84/MXfWuawyGBTDGyrO1NVxV0l1oGXd5ILE0ZJQLfDeBgT3pGJWMNEj5Il
KmaOkXVNq1jC3JCtDKwCm8rL4zZYOWCeacd4V+Si5qsd/3M0YJt96c1vZ3FKB2AySdj/8EZh8mqo
PF+ctq9cSSrpwL5K4CxHJRofQ9ZJJMA2djLGepDImjNREhcPwlrYaLJSX6laI7XJgvfmn6nNDThN
AHqb+VyxgQ3W3eoy+WlFTevCj15QIW5TAtJ6/R1hIapiqVh9ncCEUzKtaQE8CH8MWenz/QUbZN0u
NuJUpO11a86JLjsAdM8fx8phqy6hqlXpo0LerxnbBMV1zHzdcxR6SbTjqPk9Z2ttlamaff0lagwD
4TW0S1PywsyXqHRPmu5VzgeeVeCMoGnGAf17LV90xVfe93zzxoqrF38fVPptkfprBh4KQ/Ojmdsw
Ng7mjtJPCFprXkowHK4EE4qzmdA8QQLLl87ozDCFtsmcdBenI71PaMIbVevXlPsIzEJZOe/kTVJ0
S/JV2WiJKpgRUsjVlBNgRM4xcZuO43w/SGRiytD6kezLXYrqgnzuCJo+WvDkq49I8g6AA5EiyXtI
4Ctr5NZnT9ViZ5jhhGuvynBnNqoLU+rZtS6P14FDCBa3NzKUDrHk0azg/x9XNz1gO36rIAsjKpIS
iZEb2IXfhrnwtwH1pYt6UqnCCdrsnIYz50+zllrfzPkqGZhBAmXGZqLYWwNX1ttQwMfYmIbP/Zh2
g4NKdEhjFOn6cf/wCUF2xsyh647lMipBgJjng5iAonVWwwja118Y4CF0kECGnKx+TIjPDESzAVAL
LlQ/ATECvsWpq8aZjYLsX3ouvWNE4VCtHZfBro9atzHfQ8AGi6gZP6k22l4q0rnsMTao2v0U82nG
CrtyObrRDuCT7T55FiP5urJBEKFm2w96qS+5g1RrXpPvJJ8pU8iJE4gEBqQKxQ0UGU+DzfTIlPcl
alr7A5ZQq2pfrPkAB0/BiJVrFFYQqjcxwPY6v8TCoXRRK2MQqLapHvlV+sQUFt8rSVAY0CZHTMPd
KmOA5AsjT6Md14Dn9dp7Tsfowtv3dU71u9UVmK1au3e+lFym8vV8dGeAX4apGBjeL0eOMxLCKRJu
9GBKFaMq6RbFC9hzK60y1vn4enNtfQi0YOlDjhmEneemI/bX40JUZuIN2OeBkRW/u0hSNTI7hhJu
Rh9OhWV5Lh1bKWZtGu6kZ0ZgMYlzo36DZU5YucbB+sMP64CcSmtiykH0RlunD0F73IOPPPlhqQmW
v3C1WWAmgXoHiy0iPyrqKRw88HsqdnrteLONyWhklSlUbThJrvRtXsQW0qFp5MoZi1ju4N9armJT
uJPEjVw7muftfT46NmuifakBcTEvx10YgZQsAp+Vu76sKvslZeCNZ7aeTmrknAbJSizk7DZC5V74
0Iqv6KJt3lqZvtjl55mQZnGuoE06dGrDFI+OcAkhsqUmvvvkEtZcEaBrdv65+9qavp4G7pS3H9gD
Hs36WruYROB4PlUfsOX2g6jQL9j1N9nSdC/DP11GpijUEzsve2uX00U7PFnbMm4huRYZykkertV6
rHBmP3LvvlEo+Irz0BM/vtxs1z+c/iT6CpD8EYnOlQ8z+0MB3nlOCyJSrZm304ouU7LN6tG7yb6I
ohy4j1gSb/7Xp4pA0C8KDVLLLV7K8p7Zfj99xcHTY61Qyjul53Ik0vbtW+LvKfIx9d3YVWL2No7J
groy5IxvSfzRugO73w2dZMGrNwTvK8jinJSo8AmP/l49yHM8FXLR0qzXtEu587bedqHAqOHnn3w3
wOBz9ToRkukbdGqLcReKSBXErC3jt7V1ntGbEO8/7a/3cpfRSfw7ghfadBMqJ2IN9XC7GvpsxB4O
zQVRQAtlLFujvSOMWDM65I0D9ujcRPWnMcG6zrmtmqvyjg9EYRdhlqGRZmL96jhyl46OBz34zi21
3HnbMRug1SsZKqSFgP4/+EJmRa6GdNbEsWEu5nJb3t1oPrfXHSNXGOpcIYU5Fsg8aDrn+REQ5b8G
TJFp2tC+7YnzbN59fKGCnky6CAfBEbiH6WJ4gizpKOg2iB6ufKbPomYewpASfTXGHZjUdrYsQQYf
EBce8HGN2I9ZXb8sUOuFxKtJVtTxumg0zXAg4gK1uFesC7oj/FgzS6a9HOcJBDTcfqI1Bibzz7vH
Clij8IQzFHLiJHchN5oE5nBFVhahEQFpwyQE/SdvIxjBa+tFb2MRoOBVtFM0DOopFclI9ppCaCLP
gjr9aqrM0PdQserxEPzXP7G7ScLDi70Cf2PbajeQ3VonxpMsE4ZVMmORXb5hcp/c+bRUDK1v/MUj
hRqSjteFIkbpEuXzFUebK1of7kqmW/7aN03//wzBkcfxFJDZbBAiSdMPJZ0P0d3/s1wYltCSHkY/
4iaIdFfVKT9gj1gph4ZSpHmjG3/tAr1wvcupI2ZETmsO+nRR6fbueS44pdmfj88Kbt7pZTiUmK8V
vN2sajiFhKIHVJipC3EVcNzbcTtb1A3gftIvoy5vlmrg87/g7pnWCH7Ie44Bu2zIESqXlIrlODuM
tmuQWC5of4Y0QEhKTzSu4MLbmNlMcbY9R/IETvBZo872QGmMujq6C/+VhK+cSZvDNND39bpyYxv8
6Fn+IRfSAyQCTxKJn/3n+xwJ/oyf2rT7kZCkYtt8C9R/W+LpXBSwEIiRmCEGj8SJwStiEQQKhDhP
hYe1MbhAMHkXLyCvS0hgxn619GaXeq26AaCwe0kbJ2j1FtQCu1m7DX+7lU9RYUP8+wwDswyeUjpu
0lXoHAzQ1c1lY3A3A5XPEefg58bfXT3CcqMjNyhssAWjABVSkmPoA6KJnZsTZTCKBL35K6cpwUPK
XfHfHbfD0TmNdOxdLYNTTlAdIk6gf/NAExJOWBmVwy++Lo7qnfo4xuyRJPZH4oGKiv8xx7r1SSkr
86TVpo3uuSObI7vcjHNWz6X9YDG8FH0pIRFv9gIusLJNByHzxP5JSRLPSX+TaauWXNOK0BMCzm+Z
OQRrdqjkbTFgV4r5g8cM14o3D2WsCJai2mFvwe/UDQTWdGn3Z3DL8AOh5r8Me4nKVes4Je0E5qQr
pth7xxEGQ/BUSDgZcQ0rQMSevI55RXsbynJykpJmqvAPNBss9wIBhZJtJrYDQscZsIDklEMDfUgz
3QEDA5rKxmkIg8ghIorM0rjwUUNiSZFOtrcveGMDXpraMN6p22mMaGmU+3wiPSbFXeA2892KRUIx
FxXh41m1zhcr8AC0RlkWQ0bAw8jG1j5/yN3QhH0q0k0QJ6NGOhtPSG4TK62oE5CWx+wWcGdPzE53
caqdR66l4bnU7BaCZZqnCVQPUHwspzWdUlmlsiiihpo9JOB3MAZDpvzTGFXpz1Iep9mmRiViQb2P
NzEL4Gkju5eKUt7TZ6pUi66tWcDTtXXH2Ct/yS+G/1oa4eXHoeyAwVbFshF8uVTIgIcm6zssqLf+
7VaE0EOQnlbwfTgXZMuA8i3b5tefsVLnwYaMZ1yyFlO6IwNz4+1UPtR/1ELvfdecCEffUJdN/dcg
oO/kBo3zwWuNGzS0cS2CNj3rJ7f8BLLtoUkiJVtvOG+skLMFzFxeg7QKRtGmBQL3ilZys0rFRiOa
2Dt7Ti1GkIzKn2Ogb7cVxXPBrzqHxUfR8s8WETMidTW+Uuith6OiZALj40P5qW1EwRKzAj8+BZzl
BxK2nq5xkES2rz/JfdaaRaTC/hoG+QDZopXWfKuvi+z/FXXSfxCpI7XNh+OYLFcXObYhGLsglm7Z
+lQa2B51Zcik8lchu6qHH8Iw968qll2Au4Xmz54LK0+J2BA9B2fy9P8Z1eI5Sf3Mc3Cdvtillgk9
gImGYnwbBIehN9cgU9wqez1ZYqQ2d6S83nBklLxqLe09D8+r/T6AwFHAM9n7QC0Y2P2BGVM7VvQF
9MJOqLUmosDQ7JKz+qCZvPLH00ma8afLOpcgFhzs60PfbhJubvD/+PJRcmwtQzNBRCyr3k4sYZyd
mNC2BzFMhUKL8H8H+hYJ2iapAanuea3Z1GHHvVBe60cq45w1IiuPxfQZUgIGQBxdUGv18Pse6SXH
Fvbw+slj0SfEMnS7t8jb8rvf4sg0TvtyRIlCt4dtrVuem3A18w8QX0OSQifMRMhzlRpw3sL9HoCX
l4O48O+X2O50cD3c/WRvm1UvuTzgEdt1Qy7WHFyc4EQyp9+5v/jszPFNE8e9jgTPfO9M7oWevasM
T8V7pwufo/u5dAA+OmyKa/X37sHTSjqT3UJQovgJaaEN2IH2ERiP8eqvVX8Rk0kndx0xr5I37upA
/ds/hM1hcbRf6NM2Pd5kcRzJOxBeFNmD/UCLZORodyNYUZviZlejqTVMeSLzktcgbdL4uTj31bk6
uWK7RiBgWAAEnNK4muzSN77EurtqVxhwASGxmIZ3UJSq1r/4Qy3Ls+N4lZzlDrtdo6rvug4p3OCX
fnbkcM7e0MNB9+EKb7W7QA8WRRHmq6+9g+HvULhgHwhgBGttHAORZpV5qoK8GTnu3kCs+kJhDF01
yIKd2qN4EuMWDnR7JD5DhrMFMWi19cfdCKdk9+81vHF3TV5eCrTdraJ3miI3XMG+Q86+ib5uCVPm
Ov2XPEZ1SEpvb71PUG0z6i9qfgWXjakLL4Y03/a+2vrbWgLtDBknGBxKOuIPBbmD82WvSey01hsc
ZCqLFPqnJ9QymVvZgt10tftoim4HZzDg3Og+7BtBJDi/cevo9RgbxmzvChcWAlL7wUfaTNpznjYS
6L3F4SpuWURTXLE7hRsifuUBOS31AOrazJRT9YM25jXdPy/LtpLKLnHVxj9ruiyEfBB7p8b2tl+E
cZ0akTBQrnD+dkSc94ZdK080gMZR8tuNHroVrUmg7AZu+h+LoH9b0kOuNPwHcbrk67DOEQkinWu4
RjjOR11h8xZq6hdfhA6lTtUhExwljnMYq5ktbwY63WN1Wcg7/zVjnggCfXxFgr3VBBvVYdpgWUv+
1Xlrs4xguAeEFcOv8CvbfSQk4qrTZYhB57f9MvaCmDvNT4BWciRae+sTifXPV31b40jmOOyPGzxg
/+Y+yl1w91zU1Z9om8ReRB189F17XHCb8FpkeGmfjPADYnHaDi+UD4ozdT8r45oNpcUTeN/FZIEp
tMuTImMGpaQ+o80RaPYkqpoxL9SAOe7fCAcxVsX0eWMwBoFWPoxvPc9mTRnZ46H4GmbaZBCOjwa3
tZlqBRfJwIdVsjy/WmZYBNssJ/W28nJHrBxNHSswSuXXtDpwyQelkUosxiXqzCs1FjYqcpZ2s9a4
EfkqlG6DsmCSN/EImTgtHwXXNwhhuEXOgv95TfwX2Wqc8norGDwrqYeKSSfblaP0ESY9FF9bdMN3
qiXmbA5LJkn6PxGmK2sF1QzGCTWA/cFinxm9XbuznFJ1DfPnwyA2TV6Abs7sBJpjILP6d1I3SD5U
U+/R5VBPIk4uOspBWFGBYEDtZ6PH9a562jf3ZKDgUDe4G4yB5JiaIXTXWqV0vpw4Fbp8HpMQQFjQ
ExsDLrPoTD3+MgcxM/vZXvdXy1E26XTscjqYtOh8Ns3qqxuwCgENCoaTrSb0WCLshFt1vd5tKGwa
+RljgupIwrc7a7f1orsMSrvnktaXDl+DhEFzJ58zrq6yl/QxfYy4UrwSt8RkSXdsatlNRp0M2nd6
0kiYt8mTu/YoJkK+y1hxLQw6azh+XtJBhkABdnpy1aXdSy7TVG8mwr6WSUmDWwTy0LY8sR1l4qHx
4r1qUr36dKcC6NIWQYbQaZkLNlf43cuBYZoJNTZQoxm9CnnJOBxSXDAAdH7pJ50WKB9gVBP3Ud+O
/BEmqKMUpjOnr0ySARpm5jDsZetcuGJOCAg5Dr5Jpi/E01/7d0HrCBlfo17QRuLsNvhuGjQ5UVuX
nn/JkNeLPlVaLhFwXT7Qirx/ufs+qEhtXyO3h2BmNQBssEoHjXQMAQzBl7awol2pa4qf8o/p3qEc
gm8dxrC47x5IBKo60r4qotUJEbqQeGpcs+kuitVGQjNp6VtN2wJAC53PpSYJ4VwZ9GvVvb4tAIk6
f+hlTjlm8qxths6TiHxSSk4DzL8qGpICbIkRgAHisuh8+s5/LkYs4nZ8q8yJQODHduD2fjL8J96/
Hw+cTOunvxvjTZB9oX+RtTtQZOt1qXsarMHjF8byiOVMphIFnAQ8nleIyV41/qGcmyjOT9NnEaAV
P563+I2bM3SX9PXP4WbL2obIuyNjTQEyaoXTDFHSva6p9dZ6X86a3Zaeq+8UvAIjvZXvYQX4VrnN
XLNfVGAtq6p/VlWmgq/9tJlarTKe3gJ2vqYdt+3k/diKifpl3RxGuPUmWrGzgsTbaU2bkh3vmrHw
MBDn8DjJQql399u/mRegKpSLgBxqup6yZ9/mXlIvULt0rBVmra7MeRy5jVPmQvFCO8zAi5IwIBMR
sIfPCUEXK2/cFLSdHv3Tqr5bckDukeJsB3kClTVvJj/TBBKnpw17mLMNBj+senNV+A6mcxpcmukw
OkRaeKlFb5aM3RDGHlo/OdkirijWzTJgy4UNkvcg/S//y0lv1X7QiO8GS8tU1UuhmZNSJkiZBlHV
EH2Vo9zDKt630g95FYAO3fwZrEelIDSPhcZYYL9T7JrvuMNMzuJ81WuaKdBfYjrvgcW4DulLxtpn
PDtQA3CuXjyqgSgZppKwolD14CDrYKM4zWUzfgtY7mHLzikVml4u5Iu2Msb8cmsUcj5mmQbfK0l9
snJ1xiI/DHN+DkRU02NmWq/AsJKloquhM0h8Y6+cI3MQryAjufHqzZNrjwZJqWmdlI6SNXM4xRzV
i91Aq4Sk3z26ZZU1Uc7CmorSll4++9SIycQu28PXIJcUXZXb26PpaC3EiBI+9HU5qcTcvEQMzYOj
5Mqymep+Ae9U/fZEe6Xnv8472bAHxwpQDkqtJ1WPBoaraEkrXIXoDZGNLdL6uSYW8b0RKyOXw62S
FUys68Y0Ddt2TiZ3d7UOlbs4Zk+o4bBHRLeK3COd7dM8v9FZCArVyzkhgizNKuSclDGmQOVE0XTG
sAUKa39iURWo+Ez+zqBaUnUrNuKxVZex34g/uBbOL5wVbGHC9hb4d0SYJfDy+whLaNgr3ER7mNNv
LrOTl9YvE3t85EywiuBZ4dtjjqrA+f10qaBvB+kSOt9Rn/oRIP2lSiSOS5ZuxEEa8r4bqGwVFBli
9npqx1O4Q0GJWUjf1xmb2YBqvYDMF7DCPXrkP2a3GQbCzgrbmnHiFE/5+Aa40xRdJW8sd8fMkal5
3Vv5WyYGAJG5IvHhTgoc1j5Miyu9C0BeoBrkVm2AjzOOLVGr5peAS3NdaCro5Lt5Ln6bVmz6sBIR
u+ZB8+X1Dt5KF0hK79oH9OwcH20oe24PFefV/5l3xdDqzE6JyFtiwO7o1RaeneN0u72IEZ6oNraG
xO3pMUnG0wchtOg1q2RTpond2KDbcKpsE6TPqjE4/1UQAgqKNk+y6aQQ0gj17mbSrkJCG8DeRFGh
B1wcTtwjRwGEDvWhNUCveI0s4n6dvsfjUgbA5E5C1Inz32ry815rpQWLTTPu2Zdd/BkJ6V8Qg5BI
yzBKHlaIomESxdhaVcdn3wOs9fZfTlh/YUSXockMR6OmrapAEOTCTT/ZPVKrIuv9hHPXIc8rMDsY
sbEV4oXKAFUdEV2xHSALDSP9mjv7joNy2U2UJ7GMengKnir04Tkf59Z8iOKZJRQ83bboUPXzaEYG
NWNWGEwa3QUPVA1jLYRtFoAuK08Y06yXfYCNEJp8+sfBvN6+eT7HO0IZk8NlIMK8O+PO5QSUOjUa
PwfM5ABMW9bL+v2e23LHhlh8cyZMd06g0etGFumWv/p5of06qhyZTSxEEkBrtD0kR/KHCugd2dJO
ALMVQaQZXDq+4p+9DqSDsyVILaopoEannJjQaKrE1j7oedDn7QiKNwwNZPTmTAbyPDjSJ2oSlm+w
Xng+aGUewi6XpTEZvwkXFMFGWxaAaCbeKjrU9iDKvZY77n9Lo3Wtq5uOSWeAqoJxgvFoECJO8EaU
JaqbwtRTF4Kcy7IbnCa8ekrVuFbeadyrWg+I+ihoPbKARDLXpO3XJHeGH/xIyw1g0OzGAH1jQtlg
roXYjqzaoL5uPgTx79g32qAJqsR8T1+/8qQgvcxGmOPeHJePpwilqWilJC2LL9eyYaD3NGfy5l/x
21+th4wzwNQdf7asgtlzVGHUDZX5SRpIyQd7knnXoIPtwFq8PdjxlFxBE4xhM/w+PYk1W9eMQ+9I
KonqtKyH9c/+SrvrK3pK5Vwj6sDFScqXh5oRxiRuO1vblEkwWKmrXU1SirBXs6w7hISWfKUFfpuy
Hzec7WnBqTk0q/xIhi6Q9lSqTXfiKRhIsEwrm9d/YThtKAf8k86J9H3XR4veY8jYwdXNzfsQZlTN
/lfCghDwEkwQEGyhbRGFY3Ypki34InCZ1WFVENKYqZEGwzYFi74mCdQE9O8lJhgT9N9ii7sV/iGx
Varm6niXLcTwLpk+Ov2DZMS86U/RQVtqVuQmuz/liKuzL501r/bG5mN2wkruuT/FJlzn258ofhZ/
b1BuUVtUAXn4dvScSKnONOGEtDomYmbXxRabJIKnP0+jyrUFy26LUAIUtZGNmCu76DBIxSsSkCny
b50TUna03AmdEtB153w7Q1orT+vLqv/GAni+vecsKaryiHAfhG6Rx73nsxmPGwwLy+rqwr04ZRjN
QP6tb8bohJ2cZcixSS1me7ACpmkwXXGPBCs9STK08K2GSVXYHfap/p/v/ON1Zy6SNpNFsgdg9+/2
h/Ur8q3wu4vq5Z41GTV0gqJaL0QUICyZOpOlLKtGihKlgKEl9Ecx6G5EMhFtHurhjaxqsHVijKuI
GlrzKzoFh3ohMNPPsoB4XfdJI3NXJ9CoaETl4VCjbO7B5ZbFm/RVkyPe2ja9Miwp7YHYz8VYD2xM
4wJr1NnnUsAyGLoNZZ+5jRX9VqPXMwmNbVoOgxcSb3NYiFZVctdOL1e/fKOZoiA/eVfA7jS+9ixu
R2BFOE8dKNHiApydliG8flnveSxx3dBpybU2gfpVFsRiNQSPr5isPz1A81sDiYQlaTwU0bAMEo7q
acFIFaP8S8/RBG7n35mfKRuU/ThpU9LjvDygwEqFsD87o2noiyqdVpR+1jhHYbr2eNJ8pyBnCu6/
e5TZe7p84oEaXpU4T9zo4uLklG59jveCrJLErM4GowoSov3Ni26X4CN/p0TSoaIUlQBOjcz5jP2z
Zxbm14ttCpaH2rhTqJ1jIYF8Zg34hLiAZ8t4cscmX+SNDvNUEUQyvwAelkLJqR7sjeu5q26Zcujz
94Qk0Pycub4W6rKvT2IXW2YiwzhrSDTH5ubIwSm9SK+aa0uEZq93oU5KcRT3c7V9A+eNz0Dt0wlt
MKgOCI17RrrzeiF+8txNKDO3QFz8u8TFPBxo3vcCQcqUBdRx3l9EhKpYQ9UxBuNVOzegCxXlu720
SrHrCogxVSzPePitjo+e9kVCIV2nkqbfrHpgLGv5xlAQbrf/bZG1mBkDiL7BXM6tvqdl0UWkC5s6
T6Uwhwlddgy9Upu4Oaqs3INxsw7/47Iucfz1Iwx1FwRgLAhQ5z3A+8cfmFf+GNz+QcZ/zzI4N/j/
MMOnbv8y7+JntNN2mUBZn3YSZbeozezY2WGBwJKIw0/Mq6KDQCPfR0IRb5HNWeR6X2523Y9oiE0D
f2LrW5mhT28yQKAJdmuM8bHPXCAwhProFvxvo9q8bxXWFat9JF0VhVGabxJinJXALlzpXz99Pe+9
pe1+ESQpO1SPh6p0DADQ3gGi79qPD31zFHx5SUEk1wMZAf2wghNJ2Kqeo8NrbAsjYDEiTmW4Zu42
y9PoJhYWsGqTwUAFr7x1kpAb6ZoheXmdx7fb1bNabh3gkO/AzQC8c/0Vo1h8BMVUYwgsW1FpGnnt
rMyiwM0FtFMQtKOx3W5Lliefevr7wP17kl0o2Wg8KVJRO05jtRPS1PYjt3PiawDSgQXn2rIGqTJr
UD5JSgIwORcH6FWMb5mLdX9wXVlZR6WCbE+Xf/4TjFwkuM3PM1aoZXmVYaIZhpppIO0g2DfsUPMZ
j3sWIjWHsn7vZETKx/y2rMxBUFICDimStAM7dy52vMy3FBoXeW20kC3ygb4wGWTlC2J1ffdp2xFc
1Ie7b79Qo9tAaG/DaRS11FtV6dH4VmNTl/irPp3Ugl8yRydVK1oChQoJ9UXP2J4p8bgzuJPqI/Gi
lJ83aMEVO/8dWOVV/1dfGHWN6pKX7ctZqcWeZQ8QvUzkUP1woZ+kGg4eEtWrCRguTxF8EZDcD9gh
QSeSVcff1d0R5zDpxztLpbqCj4fHcdtsQZjRgkEDFTQkmVC8CPlsz5ZcxYAGm2EWhVQRruHrfXZV
GJrBymO8pvtsxTI3cUi6+fUkhkBpMSj0ogVNs8a7Ala3SyV00c7kffYUSbjwP6g+kg0fV4kZ9Khr
tWEx45ccX+HmxnmkgRJ5CCtcOv0RapqlyGUj3xgEveN6SDcwipDlY43XtmDL6KV2D3oa1qLgqWCT
tFvo/nYrfjQDO8ZAeCRPDhTZwTb2RF80W03RoyMxiLknT6D47tDlCeBkPzfEXCDDJT4hsmJEYMMH
Yn3Z5D+jC2rHMLovbjC3rpWGs8XPR7a+YH7u81qdOUpQTmsXkPPzXJPDgKwTZFiqbsraPBDEvuoA
O9QtHsrqs3h3MP2+EhHRzJEs+SWq/VOTCSuehAWZLrhT2oFQA3ddVInCaguygfiunuBYg2YhLKtC
1dSGhbln9PjXqPnZAV4JILJAEE9buTdHYLorkE1gs/w0Zy6qrntlEA/0T2qey1dX4K136G4Fg7Mx
86mLnfXE1wVm72XthR5zOK60lORZKMKZQc92eOZ2FK7UkxyMrdBcdA1l/x/QZatXl2MkMZ6UYwfG
co8L+AECIdXezb1/GisGTCiOZzqG9lR7cPtjgFyDTBKN3eCZB26ueJPgdCEG7IDvjciibnvKBLn9
LxMhFiJWAHZqrhg9wdIddWkrbO9XAUsEF4c2J24to+KhK6xNDCV+U2+fSOi4K5Wyh7S85ZGSqUYQ
Jvn/Y+MQlkHPY6d+ey/PXFBdTu4pI4h0TJYRZcU5VrRq4blXOGrzdL9bAQ/5Oy4+iUJszeG1kwiL
5KfXBNBALhk7+eqgAabd29c4M5cZlKIWGzguw+BNhsBktpI6x6uL52mfTlqb4bsyuGmaZgCt7EAG
nmfq61KvNfwBDK/dUD7TXged73i0cgPxQdkuzMECLYSFGJCX0+A8OoVDKf8FY/mW8sOkHt3Ix+9w
yBijvb1Nd2usKuw0kX8wZWLI5ZAVp617WQKHl74j04TM4dGKuYC/bO7ll+0QXLG98OYb4Bbg02Hf
xg8AlJIaImze6SlU/1H/aj26vsMYoULuQwOJjaO6uIjYWc26Mr+1Np+gG2z8a3syVnxKTev3br2l
ZwjVBZP/U+YJYCYdyZEaA1PQOEtlHjM1JaYI59Xe71JPJGmWXzwaMg6qtN38I1I/2cC7qWiThMVP
RLIxQZkg7bA6sT9mLgwEg3JnVDdrsgXsQYU0o/oeVA5JD+Aiw4RUyQm9t806b/UXoEJJF6a7NC/Y
dGsPOSXeFBrdogC3/hxo95YWVY/WWTXIqTByGpE3xHCYrVfFodrp24fvlYCDSGQkL4erKMT/jzoz
M0F8SSsZ1DVQ/EiZbFfhTL//AKzHgz5ivEcevjmt3bu8etdoMhgNloJyu9m+t/qMNOSX0B68+6f/
CryxhLuGHuPzii5g7SvoqUGlWb+o84cRaUmR4QTX81ti1iTYzqyWZzqygj4vKf6Knd1x24NuFkcP
jcAJNszabYWdNGVJMUHZ+d2jajCIX/OW5E1VqJ+8tp9kl6GOpFWTEENEUfW75/KJPsu2zeYdW9DU
kP3qnJ4mfdiGeSzqT07OpDFhFQCiOxh46M2Nsx/vlxqL1tEAaRTOj4bCrm1AlHE2IMvE7hbOfhit
uUsi7hKrtcox6EOtaPJtIhpvMzEvVw3FHq7lCzZVMY9ThiP/Lj/FZPp5UYkY6UPuor8vyXhTKHMD
+ts7jLIylbmKU6KSQhWrVvMHys3ob40EfuP+7njDRqdnUidcD6SWpX8pWp9yBAXEerTLdfb2W20r
S9nvwiOyt1JMhNGAkhQyEf7FetmOdS+N2m98+aOTHhMFBvqFJnF0JB1aA8QmdHg6sFlcUSzAIOgV
9Q/RbA7/GdNFg6UEzeyj6O85HTGf5OIfzGdutmWRW1v8XVB+MlAVlBL5igkZB8ujq09KpCCl1xvA
soJseJaIsimJ2VIaHysMuZ8fqLAGz9lLW0BmxvIqXcb/dOgzhNPZt2d3+PmM3yDYcG37WtVpzZCV
iyvR85va9AbJglAocijnYdabLBg6qLql2RGN8TXiiyHBFqYSVIdSICEWea+U8jOq2lMHtoa7iRv2
+fWDpjE0ZrgBRHdVo6xaWXHuG4u9TlHz65v+yG17qibnXEXTkYie8lBf2N4+IYPEddDZUtcxJ1E1
Aznx8+zb8UtGA4HKL0PnsSPTKsuaNCFU2RotTf9XuF5y7jYDRBcjbhQZdcSVEVrKmKVMoYwpp0Oj
IO5tu15SLK08yC7sUXvIAXmYKkUYPI6GtVsrHA4vvnQw5EXQc/p3EtqatjUAA6ZYOLH2haPS+jZh
VzDrHv28NoHxKj6xulZgVOxgrPSBbrvpvJAOOdvhvMCbejS0Uzg1Hh12HAvmV472XU2K8np1211A
CxHtDf/had2yGN1/Ueioo6lVEW3VTfEMfWfxZtVfiXbhpTlyRQ7s559vf0Hcf2phvCIWkikEla3o
EYz9HYKm/dBQPB52eaFQ17/6M0WmFMbHVhc291EceBeb/am6j1wTpqT72xqabGsdVSWiSvEaH0dD
8lEoxbKO6iPeR2mCVrcXnT+lkWObFAtx3Fq2muX/ldrIc6dGpoSJIQSpzrMgKS+OG+2WcS5XrPTW
KCtDC1iDePorArlzSWMd0wG1dQDZdyvJ1Uk9sBGu/HN81iT3XFYfrygDmx/wbcW98HzXDw9b6cnL
hRA1k5t8lYcJGp+B2ideVueJdadTxf3uc4zRD0cy4UmCz9/1N7H82P/ch9cxBWG9Nxus1uxMYKyi
n7Q6lLGeVAFom7nwbFvboaIACmHLBJAVnDrtLBoYr+ZIfBF21prKa+Q/39wuGP0nxrEfFkGQnCmy
dkhAFEV7Xu1F57Ug9Dqjo3ZOffhFV/+mo3+oOLacYj1ZXuAfv0krhCZUql/SLj8rg8KNsMNm1TKZ
0zmObGPlxAteVCXRH6VXa7GzuApUEePMRFxsSksBjSCbfHKacgRdESSKEEupQu5yCH/n6AmYCfBb
xofOJX1Pk/k50MOw7hpVuqaws/qklzRCvRDMHPzfrnjKOsjPwrlmN4zp8GeaVOyRts8DhcUCDFy5
fUDOGl9ujQnn/U1JFaYHNi2ZFpmEFEBut0cbaLawacnabhnV4VKqsbxcSJ503FLDogia3atyiK3h
e/Jutt/lfcEkrjsIaqjNK34q0ughH5/N3JdwNKYCy/uviv0tdt14MM2PzacFsPlfEtlfXMRY+VUz
VUddh+HaGqpgeRXC6/VLk0wUQpxUIyTwROzuWt9lrTnwB6YinsjJiyUf8X5EnxAVpvyfrsE7r9hv
NK1l5EYpWXLSroFQl8XE2NWp+6ZpIgovmmtueb0UGaRfkQjtsoStTSXZLwDjn0eJrAMcp9yEl6Oq
IN/P2Rg1j5Q2m1t6DnMmx3iZiZ1ANA5ctWJGfDg6qVroVPe2EL7+Xwy0hnxJctS7X2tYEmzZ3dbB
r8SRUbZ7HKEUnTteH3uLEK/t0yV1iDIdFi7AvNkt4P7Zyg/TP6EHV5U6d2KNt78XzqowR6pkkXkO
WBP92TtDURWN45BY5FjpH1ov8QUqkkXK/jCZA4uzfZeHS7zr8Z10i19i1GhlbE+JeSp7+3+tATsz
lNG5NFLGeXarM2h/bri7WWcyQlqUneAGZo0GTQU3dNKydiQwaOHtxJ4VQNxpXodzqCnxDplOcv6A
XInKC8BIph8mtS1IXtRG7c2bLenPetf8BmS/7dwPnko3KVdv8kkE2754y4iIoHAJ12hbX3WBTVRG
nabaDIadOHcEPNyf/Qtr/0r0qTR4C2ck2vVPHdnxdga+SJgTYwEOCKx0G1jzM9ZFAnXIqOkiAkuB
Hw1Lw/ssCuaAPphLJ77XT24VREgGhUsiJ7YKsm5qbgcwhGSFch9vfQZbJ80FXbAgrgtWisocBHrN
H3Uqu8czLLZhkygzX4rZWFQsbHoLqGi7h7/tugsyQgoEI4EnBfv8MT40X0DssM1+sEsvT2g27lKM
5ZUzBIma/XLqt6pvwmWJNLyDvPdDemMVR7PEf+QSmcuEQUgvQy+NxhOxO6YtBUbTsnJFLecf8H7u
grqsLUsNDs9MInC48R4Uziw/Q3KB/1uDgG5iuZ/euBBHOM2LCk1ZVWb3FCaJ0sDrDM2xT5PqDkwU
5JpOisMLevNgb5a4w7Wq4ZRhT6PWRabqrS6OqSFdT3GSG8975lQMmNlvCOofxli84NuZkaUMlBMw
UemB+7ScMH+pvbrPfnuEL5o0QjiKADOO641IUVYA0FEaM06jzIok1TsDrPZEJe5tDCmj4Mbs0bvw
VChlEick6Teg4BXY0TS2I0hg5n689rWsx6YvFizSdJqpTd7la0gn7q3to5vStclJ5nfdOI0PP8Mo
xXN9Gydy4ps4J3jAVmCZVm++NsoDbIawCP+mb1tbMmwpey5iUDZSWY/zik7VJ9Dok5nTXw6BM7Wq
us1b9gN2pGVpq8SEXw2uJ8EOLvij8SJ3LSflkPnKAAwvhcSns2jV6x+7/IN5QxAtKlFcrNIFPdMu
8E4hCbcstyYVtopEHVKg9vQHdT5dT89TaG3mIX+zjodH6JJ9Ibo60whXOq4T9fpbE7YYstyoRx+h
yI27FUm9hIIrW1i7K0GXCkF8B+J96H/Bm5W+5kNKcF7PMcoPGj6YpehNay8SX9Vm+mLupNdu9S3E
OImWOh/Ms4slc2DLHLfWGS1u3IoyW/0KHarwjGhGM6r8Mi6z5Y3DX/KbQttC6TOpNF7WubjvMcne
ybl2iEHqR6FifniG/Ov22Z0+7DSvOQFc+zbxLnWgbVoJL6tTbV9LXbSHCyVXLKUV2BbgkWAWZfVV
wp8FNHqBZsTu7b4S8jZR1NSjiuRw8fLy4URX5oP1KHfygsfGsUQtEis+DfiHvRsv2lF0qQA9MJnv
2vmUU9KUbDJnRTsLsqVr3cr/uWIxSzfFIsBy/SyglEMQLy45fIp9nVSVgon/q82WqW8RxPtpdMj4
/B9XwQ53QAbdMS9I0lJLm6LDNHyAdekFvVlbtBNIK72avUE12S3DhNrj2tK8GdYVaopxsU0ZgFfK
b5mXcyrkWRLB9YPLXj+wOaKtOD9xu/GT7EuDC9EydGDX2guUeuJa2QqpWD84LMrkREmedWy+yNMK
o1i2LhAfrO3kV3AmmWcOQfP0mYXi9av6L64GvUw/W4pzbEdv37e9ML/mNQ9JOqc6WfJC3kTIfBuJ
//BGld+9UjB37dptZnCz/I9QbXHSssSu+I/yS1ijwGNlLIMvhO8TShCOtt/2vcasbkDprsUER++s
r6N64RrYfkEbSwhM2c09r5ZTmtiujSS2Kx9eVQoIb6IORXfnFkL5kWtung9aWeChndsHi95JhBT/
AY7NFJeLyzPbB5D1c6yxHglVpfMw6MXlnLBK7nV2eqqbZA3XdAjNyxD0p10ehNp4D3BM+13Hv67D
IHFpOXuWYhgK1BSd8uYYFn/vhtaGO3UfqL+BTK+HiiaCVpuYaOynvmUCe9Qi6NO6nBTOfV3l7i5X
IYl2raMISXN4NGCnsH0tBppz7B3a/gB0yjAheuLTb0opHn6+h2et2inO8pOFhO9Ewh1/qR0nPF4k
s9IyAo/9lqWPvRMeIFGQQssj9O/QcAxCdBA8ix879c9zu0oib+F0glwsxHN9k9yD+5eWqJVAPE0q
BhIa2/xLrB3EkhFFzLEgWl4xG1TAQGQDgoqxnoUSbhIZ/VepsrmELRUhYc1vPlXJerg9qmW4k21b
xXTIZMiMkMjBXHcHLrka6P2qBAfUYegre5+ZsEzxOLWD8O0mCfirhfYbNUkGl7YjobizxXK+Lqx5
Q8OP2CI02E2fJVTqvBiiHj0ar1rczHymEn1AiZvOp2DiZlRuQ4u9/tLMBzCUf6so6+zBttYkjEC8
ZtN/JQoqiALWqcZcGEAq7AJk2cYaUHLcJxGNZggFiizC/ocMMl4n6Z9rsD+xnrA8Z85XyB8QZz6s
tnAoZR3bJxosaNgumXkdk1XOcZH8m+6FZhKX06rafxyKdLbfp2d06UOgtkBO/QtMjJPx6zgo24nl
0zy8G4/wvFvdczhU8uS8ctmu3vp+s9h9UFH9HxB8E424PlWDA3bk+qv7j3CEMMg3fPSTwYmqB77j
p1uYqUu/9caRMPBNkk/nS3wfv5pfn9hiwyzBSEOSaFOaLCpu4rXQ+n2WM7EacME2FPlb7Ypldzgd
eJBj3feugFCrmKAm6hV4m94uYxOFvoS0E/ErWbhaaOgZDmMfVu6f3nJE4MWjur8qGhzKbcluzcac
kkq2KGIVYVonyNpCq41kpuNGT7S0Qbp5E8pVv/PI8A/vWbYgPSIqRqDp1YTULE7IIu6lfEpO53X+
fc54MrI1RFQ2aUT053ydNDxbEWU/P0+14OJV9ZoHAeAwKWvYvFZen48ASSogQgBHZPpehR/ogsnl
/ms/29YA9fm9zuzXonNSQJ4h8SPyDcvBqDZsfwQH1lg3EovjU5ZLGGKzbMtxYsAmXHSQfeCLmUai
lDytTx5QYAd3iQn97iR+mhY+dMfcLPv6dulvQOBFLeVE/9ooU304zhrNeQSvGjjOs5UBu3IhWgL7
nz/zdqWXD62f3m6/HJ0Zsoh6LMo8yXBl++OADf2geV7ePLuDOSpF5V5js2mXGOSKyZPG4rnnDVzZ
MOlXjCw6MYROxWyNRO4+wT9nmTl/5vktEHTVoLvHF4nj883s1i751hHoQADecpJ1DEXDXKhcCz/C
XXeZ2cEeLVcZQnGXpEnt71NL/5Zli5ET+OP4sHOkqzS5J70lIcNo7W6Z7Iqx6JYYGR310XOMDFww
/uWFWrH4DVMeod9+SqK41zjlbCop64dTpZO3aDGGnJ6A7Rg/CjeXihIcACEGaII2uzMcDxvTVW3o
EjkN1qiP/OqNE5wBXKyVf0xwjOQ0k0aRwv9DTUsfHuVvS82cTuvT2co6BssMRJv5Wbqtuw8uFIq1
Cg+xNSTY6thqDfBh+ONhDdGMJgTc3mP6vt3QAbgelpoEC+e34wYzFmw7LUaCkIsEdfaYEBhYFGYF
NdyCiQccBkmbVUTWrLsn/9k2qmKFD9ZDZxr2QXuD7le9GV9PkMSkGzjpWp2JSziRDTCtOlwQAROX
K7PDtThfrQzw1E+LvCaiR+S5wdUak0q9wz67Jwv1jgHpI24fnswvi95sj9VCS5ka14+/SnEYnlNb
gA3BjhvLvcNGPjnbb7KhyRVo0jnesDrefv2tLIgt4wpLuH4aJvcLpjBk3pCzHuUXPafImSukmqeR
fpZywIlvhNUsnOtcYRuPpSVNmn/uvKoOf70xb/PQMAWFtp6ZhbTDihql+C0xkv36aRNHjyT0ZJ9v
aiNoiQXPl9aXK+Z4W+Hc5rQ6H1bY0qr+xCkcdDEDtpIco/Oba9qzZ5jX9N5EkkbqjiRSTKAXOv17
QavE0xN+j0bAlJOV8IACYJuWMr37yuOr5V2TZ+qcLzv/CIkMTmG2vzJi1a5q6Rdl888UaEMvJiSz
gQfm4Ay8orOKKT1l5TMv5DynNvacSBmKqwijGi72sdmtFivGYp0ObF6wsSGRfAMsROK2P0lceywF
l9V3oKyQVXmKzCKJQgJW6DriA7r2eFVlq9cE3tsI5L4FhByyyBkF2DpHinC6P/YCL+uyhKgi0gfG
1ohuow/KgqsRqek4qHuZQj1RQl3uAyfXuxA96EXPhIROy7Cooni30AYTkoTmMwaQVQ2k4oRkPkv9
KfBnzrDfNs36Aob0nfF54alLmQ0bn91YlyJdjEj7Ey4MUUejYIjyK3mZTyjf8sKIPjFFUXEYaqmy
ot9CbcFGqap1IDMbT0bj54R5T6EdTg88GTRz7jY0pfUDVF61hS0fQKmehN451xUNQvP1hK/IgQoT
WkvzVIu3dfNQJTty2UFbJozHyxJ8iP3fLZwn70wkpwyjjJKySrGCQKN6Lvxr2bnrpON3/EmiHZ/x
0pzFG2fc2/G1FiGWY+uFV6iPqj8VBJonU+xe0olxxScC0XnxOtpx+DzWbTMPVWNGN9TMOFbtnDQ/
xV2zth4YCFAhxaAWW5UOV5sO1R7LtUmjXr6LOxQciAVgme3eoZvKONcCF+qP28v88Ktc1gobQ/G0
cZB+mNQiaZR9hgEudW1yfx+Ddn7eKxebVRDVB7SuIqiDuw7rrvVeA7vXY/WM8P29ah8iieRHH/uw
AxIXb2a513XyV1Js46xgExz912nKWzjRdVLPJUcwRchK/1XbPZQnagQssB5u2GX2EPIrr5g7fBtD
HoAZxEBFWKFsWWyMwPerfmbZ9nG1WtzvFPJ9sYFyw1lx4K7YxGNg5rtZ0to5t2ZOfS7vGtwjxfXL
VxdOlAKdlDZnO4wIhJj+pF7eu2RH8+sZx4yPW5WUC3DwZn5n9D8QopS+flRQsp5EQF0XVn3rvRqo
XmXRjXseC+2FOj4l/huhyPOvpJ7y6GD+SSJtdu1/aiuxuyc4ktQ9BYy5uGr15tCinFHgfM/YfOd8
q0aFrx3Pfb05jhOoQqi54mBG6wYXnZGOwc0EY4wzOQ1CW86xaL7MzP0tbQIKtosJp72Tz+K439sm
u+qAXyRgblv9MBVYnak1kGTQQQUIVvAHVdzAI6OOEPHPmyhzfhSaQlo1YdowwZhsGLcUUqApuPIW
w6N2S8zKmCPh0qvvgJBhXiHux19DBLjKJYtUXRcbxYUNg1gxSXIbQV7DECWpqt0YPkDHHm7JEmbw
ZXuF8r0xKCRF0H6raGnORS+zqzkRkKR1UTWHVVCv3kT0GIyfeCiu+5hMj6VY/tsE6OAMUGIZhdpC
vlvISMCf6W1wJWV0nXVEhv5PWScQ8brfKdId9Ud/Ozau90C0ChxK+hEKdGHIFSFMed7q9J/2H4f+
K8FNvfP6AO8ZNKnw990dU66k4SISCzB3SOEGnrndANv1yiazpDUMqbLQeq+Arb6Ei2OrNUoGU3af
8ukDTCCMZBlHTojAw8XbpMOfwBxOpXGWksxBU/xlVaB5ZD10v0fTGfD1XLTKw0xaretDyaoi8OOB
RoOKDFIDcNwtRVRxPfL8d/IT4yT7vKd1V92uPpY+RMoL0+5V6ScxfVf90XYpoirjhu4ROuoeCV7B
01uu0q91IbZ06QQX2JStvw1FLuV5XWrjxXIXqjNMHO+QJ+N/UF4M7Y1lMQ5hZ1+ma+hRcTDxRXE6
5sPKRDsYLWLk2KAKyTAGQlXrSchuwNq8NfhAN4urRr7sgXBWDR0XhWPv6Js1JF7qd+CTBJYvBg1H
MduzyVi6gkn8jSHJAbuLvvp/tjugXyqAVa9Ce/npcrbW4CZkWAr+4tliunAmrGedO/rV5fDe23oX
v70d3cJtcZCnGbs5u/O3F2LQjL90JqHomiw6cH64GeO8VL2HbFYrxwF5N45cxg0gtuQuwhylGCM0
QcVEP7raeam2dKZnWlvVgt3V/kBaAqZrxiNBbV27CCnyFJ9Hy55AFCuMRw50r9EQmuTho9aWW9sW
mVaKyEs29CKELMrKTECHkyFU0j5tXIrJJZzk31EFvGzRl6Q+nANcz1t8ih7/Xe/QXa19WA2MeVrd
mllu9Yr+qJ5ZzNSFnJLBkbue3wB4Ea6VmEr8ghQ60lrmnoDLpRpjl1I6CsmZqrR4gJKylsfgnGDU
MT9DY21XYxVf4OPRDJBwLO+ZjMREoWTLkB0B3BgsOF/Hx4mhC1kM8qKouMrprHyYG+BP5BxO6HtU
l0fk078F7ytOgmFbJuaO11QNGgJIcUrLSYRolNICtgVOUpHaFYrm3xEX2L/RcduJ3jUxdujNFG3n
pVl/A4DO0yebaenF3gilukTU11eKALy9oqP3F0J2qIyFBjdlF3tdgirMyHGqyLrKcIDoZg70xVyg
EY0E2em0T9157VmFYNSGGV3WA7wVyu+RfSvBhqBngO6ovEb4VgmkIINu/RNuvu7vSlmPfxfkSi5q
j1kba950qBIXx42LulhslOnFaiD0NRrROnnBPAPPsO2TeVICu8uFL4r8CgWvG2qI3O3mbKIyVQa3
tTeprDWe9EzO9WkqZDSNXlc24iW435UfdzxxaI2DOYj4S/IgT4UduJbBCYLpTVkLKJwraajphCMM
6D/HlHJhPzX2O+/0wQL2vWiHOIJ/uWXlx15KrovPGs4Bvoz25OZnJj0N3ANv3x0zLEu8AwdDL6kt
pf2Sezv0LZE2x4vg5Ganzx5zpakYd29WIDQFNNfNR3ZtxFN1PtXwhxDQFZFQCvLHskNPEH/LU9bA
tx9mPo3aE16EZmPDOTjs9tIK7mNPwBu7CxLsoPM2kxld5zJ8mUcmU6mWcCxIJgbqe/X1RjjtQe41
xVwvQJ6fhtwGulW/mW23ZgbuupG/gZfQx0TG6N4SYmpcZNPgET+zNojohof0UbhEwds7w+VH0RA/
blYlIDX+mn9DlOmXNGNVaR/NUywe7EXutCaLopKKT3jvC6e3rQTpEho7xZJmU809zhaTHHUfEaG3
8Xd5ds0XI+g9v4Xc2Q/9DrDWBQ3JGURmHqJ4eYTenG3r7IFdFUIWoxa9PlmUmZyRM8zUHAYvI6K9
60/1sNpLXUukSzX8N+wusraTiCL+1xOAykse+U9Y4zyhzn5tHyan0KMQVG1iBoPZQd9/ogVaE9XQ
fDXyq0rdcuZDKRhzHpiqZsQAK3M+UfNS4c1rUCQaMwshBjhzRRz4DzMV2nnC3530JwlIv9f0ppbm
L6ORbHxGM/UkQK56jYfjfH4+/OddkTt2Gh+C7DgO8PCkekXq5Nn9WFhLXIw0TRw+7yVw5y+uti4U
PnO/E5I+RS6TSQ64xfz+T+b6zYzadyym8YoOaB+rMPQdq/2HCI8RIzieJ0vd7MCCjiPFazYcQ5M8
PjNUrP0ME+lk9HBHCb3OnJGf9Dg3qKWuhI8OLyRt8vpWr60YEjlQdcFkxbyZylSyg7Tjn3AaF42b
2xYq11FBnaACNdO+vTpwCGx01zMz4dFIN2pO7LNDAftHDAEAJaM4kO4FQdoKkTR54UgkJUCmEhbE
hr+obcVIm9j2Zeh0khIWSjv4wlFJunbCDaw4ajIThuAiAmqHPK8XLMAT8io4UZRDNH6Ktw8XAtmA
ojVFn157Hr/zFEPJLKEctGBXaEaRGh+6RvtjICu47TIGr/SYpcIR5gI24/6eDjS3pGaHlUm4Oqq1
Og0uNUZaK+jxd+MeS96PzBl5YCacA9pv0jIGxDgXtubDhjx5H6Bl4+79VX2Y6dKP+buhJaT+aF2H
wWCCR19rJn4OsxrKrDINGljBjsZb7hP306UKkh+hyfhOzZ85BJ+/n0ZY24IqVp15Hf8JKI+4yzfT
e6oixf5Lmhk8bGKcHlYMk+icPhc03PH6lLElAMvdPJeZhS/sBqvNtkjD4TuhF6lj/SjKkGeAa8HT
9cKFU6ZnxYv56G/Ma+LGw+C30rH41AHicfuxs3M8Ec0x6bdtM2AZoBKnBTEp5ZoAnLAhfqEeyJvf
nN3vGek1tYxqejGU3Kd6hHlS72aaAAJwzlyn7nz1LzNFWQuueuyQ76njqdGFq2GQiQ6jW5FFsw/e
wpbd2NRFBPkJ+CUI9fo2nvRe4RHYjb70m+faYOduu0Bl1MP+cUAIybmMP5ii6HIUf8GL6AtuuEt+
ktLrS/CgZaxUwV4Ow0MnkxvjD9ntclxleQ5H0Aq8+5o5zjtNGACV+CLRhvcmCrRdJvP7x97uUUQO
5kFlVa6BX3UBimM6XfqM29m/UEiOcQi2D8rmIFn99EerbA3VvdWOrvRyay5vVdOex6sca0hqzNuE
TV5D2/WAtdglGcqxekvRwF4pYcWtpiX0LztRqHBByi33GJf4h9cP1Ah/YoYXrmRGoEK5Kc6Pojq+
KHXVpNDi8QvLZq3t1GSepasys3LzngPHlFrKMtU0KqVvAx+eYzC50ABe1Gze3BDkP6nHq4dumsAt
JzjDri8CKakra/OyawAKszmwN9LyT8ZfOXDv5cjKK0IOqRc8ZEIXuHSKPBgiGmQnqK2zIL2SAJLd
Xfev0OLUdhO83uTOARWSp3UFuWTQzzcR1RegOeez+PtU0iezoD7/wbY9TocarK2yP0x+6ijgg/85
V9CgdCbmnpa8DOmQZwqCN7Xg8VW80+Xz87ZuGIHZ6e9vZUJGHgNsx81LTtizEC39InJTL9pOIojA
i8SqsM1ZN69pbucyQRALQbCF8eikD2BThts5kimuWJ9u4501w//GPtCojuhcRCdzrgHhPs+aWHoO
IDxKSlfYQ5A0I1VqupicQT8u76TheK+h7V3DqeLPtf2xfqAzO1O3qazK6duecC5djyvPt2PyRN+h
3QsSl1xcF3RE+rltyvD4YByv0KJ01L9BfRe3cx06rdudIRLBUZ38bTem6SHMSz9LwwPkpRXddQy6
q6ZUQYxCiY/A31R8UMNY+i+iqNUL/zr/LdIDGr4IlBjfWn6SjPkm7HhBR9dEKaBcDtR2T2mHA6l/
9fry40RiKoFsVkwHmC4bRkxi9WOMIsW5gXcecYLGQJKZtKM0jEkAtwei59Y6Q+bgw7Wf2nULrizq
Hi+OB9zT3362otkWGqEfGvq2LpuuPPjfEOzAHBBfHYuYlTJekxaCLOr/6vG+eHv7BpXPRZ8686DK
7v4TTkpEVLXMzOccspOc6cA5J4R5nj+oh5ennZyLZX8ExsHF61Rf9lXxDo4ShntkQ4ZjdySMg8de
3iVgGFCqMtA+Dhqssdc7/GCMFZNNEXjIk+F5v2MZWBJ4LIWawGRPGrLOs8ZuN3GQLeSYDq/MJQHn
kq0p8evtqaCqh5NbMgivRGUmQufOaBx6xTLy0rouQIEvq3HVUPTtgtMphT2waOJUYIF4QRERC7tK
1XK8IKkLC4elOlE10zu9Zvqw99X4TgGkxTNh1AhC6wFMa3tRaohySVHMfYCBvpMpQaGz9AcbZGnR
gzdYaEUTKdt1FhyYMF++uGHFCHAtR4gQory6YwaKoY1ePpkF2uHCR0V4eifbfXaTaeI6RCczCQJQ
hJIHK88Hm0m0zG+oaFC1PyPLNp1FHV4KdGCj/myIeyjf1veopdW/xHs3yC0lSbdNba7VEuQudUEr
8tVIE6P1gE8f6xkxtQducV9lifpErnOEQ0mgsQ2hnE5BLH//G/GMzO/hRelHoQrQ8WBqCSTjicpB
30AOBiCNCwPjQRu0rxlKBaBLLOjTfXLepMaCzdRmF4RmuddgxGVsnelqEQU3Yg+YcKvqfc7XP8eK
A9Gj5Ga+Uo3jpLPQOxtM72m/j7ei34b1PTAyhJxFmaSg17kd9v4rEIwwB9CE49Pfi80dRtLFxcFz
BX1C80Gc9GqrI/8J+GwB4FawGPhclwSuh/iyAhkpGLth39jPzVYd2s8FrWVP17j/R57hn5QDoFmc
+RUeAamhVg3D6Zgu3pcjDDnQOXF1Ayy2yHGLGH8RF5MOoQlkqO7S7PUobmulGE+aPe+H8saFmiNl
9MGnQ0NmXZHTHHEQ7cdiy0XI0EqolpC64Q8U2UoKoZM7kllcwiPEHQG6u5Sh+1/LN6nAYw3rJxT7
G2BbApvvcz4l31+mQWMmdRht9Mj4jirnYMxSSCryPvt4yhbfGrEuspkkmekkA8F34BbUv97LwirK
yVFAZB73MJYLEo8KBGcr02TPxS13xtNfAvPwLlRfCbLmQ6ef51MB2jU9OxT2Si2qanUB5swqp6Fy
SDRdqgBZU0liIaK0AylQmFB8xEsJ5BvJuzk+h5EbnSnRCKYZAbVjgiH6FrdzYeyiSewPgHYQLR8O
cpUt0yXYM0N3JBh9HFhuE/7LbmiadPORMbO6deMIwVmVBGwjw1w6NqukFqhzApKCcRea1GqYM5bV
cc/k/+csAp6Sl7sU6T7VaMx2Y23MUY9LZ10x3gPYP+8kDYOklijZbpX4HIlGm3hVjo7DieUe602v
IZ3xHPJydPCS0ugr8bopKc1gPJ5HmMqW/zP1I5EvaxIQ+YqOy3rBR974Oty0k3ix0ZbsMztu33lO
936AvMZY8Rq+O0yClVwr5Ct6As1KEEj8T/QSCWI+FOryLO2axrFXGJIUnVpty3ynEyEtyxk/jymG
eMZnCcDJO9UG3M+P1SdBv0RL2u/K59yOkk+GCFHceeGWjKshqaKHUJHNQcpPELY4K9fBfrmuirSn
9v5HvG1C17AB9gpj04EJpS4gbXidhI0pFPYgEX27XZvJoiTiV5RZZ5HyU/8TakXfkpNUOW80VSGJ
zO6zqHHyVCtmzkEij2kf/oYpKComlHVrgfvWnBR7G/dO2zT2WuFX89NbVo/rGuuDzMjfmAfc+3Ta
oGBcZ7g+5eEO5JhY6v8VKnjLd8cl1V/W/J/tl9YnddACKgZJgRrucHtVsBf7lBnx8q0E4qy4EbDp
U2y11S11hujCGRAVgzPSDi6uNaq+/YFEO7Nodr1Wav8IK5bvMzhLPoS+fz7i3zY9/Z+lVlSllyzr
rKJeg61uaA/2Ts7mftlw0qx1k6yw5dpT70JxiQWp3BzlZvGQPYIjjoEfZDuAqsET2E6UOfyH4T/+
RCyeHSl+eCBZ/CsEMIOjfRZ0pFGtvJEUUuScPw36RiDjtLNB9SClOHAxj5SkGwFPDTol8E4EZOyD
1HNDwx/CUViHc+bu1u90K6woNFA+1sBHRaCuxwI3CH59Ms/dxO8u3hT2m3pHG5+pbjHQtTAhieoQ
YoxhYxcmEjPYmmm0PU7KIgVfheASXo7ruNTItniuDJSz/mtxeh+oCOTGWozm8vzLYLoyhMsEoxb5
398mRw05GUcmAv07Wg8KF/Sk1aVUNC0Uh7CXRVal7K5S/+5d8n3UkHOSNebnPWu7J/d+I/OmYaBM
ICh+fOtP2NLql+848NPCrz5f3fEU2WVamUwVrVA/13X/3bSlj6fNh+eiKcE+OPwR7+w3B79HyyuW
ptgfT42qTf1NbJRh82vmC2zLDMxWowlewFK8gb9imtwi63FQ4Z1PSSfqGEXx3cr+3Y5sICrqmKcn
BzpJ9AXNiatWkoJ2HjEN0dCySXoHHaiDCgnG1NjmvzWiIG8ls/F01378MjOWQ/Ju0r+wSl4iPJVq
6n9VhiDIEtQbc+BgySk1AXUwx10bovPaQAulgib9n+tKssqnjBD1XcCYiNTtqi0KkoT4QybtPzBN
2SAiMbAL8Bt+IHV97pfnXBD3Uop9hrQYOO9ZKuoRtWMGaRkgvCBPArm4L6/qwR0tvRO8+0EoBofq
53fT39iCaeVcvJJ8SSE2NTPpunPCfgaQXAe3lupYsqzrtMHDI4C/4lNzvF9zmmffYHZOmtOK7p5H
eg3Fl1i/DMZUoTyk6HwgYGWPvhzq7UMkXnT79UsjU2o8cDIyGEhPRqzM+aumcpcuEu/gNrZq60Cf
MYXqg7mIODaIYaBt18Pra2AkyitWkzaII6jdhQCq+ERXH1+bOIh7K6PEOeGQyx4iUtlDphMYOs4W
VVVgEoeaCzP0U6OKyUkzG4cUiReuq2oE66xioGSnVG+br2CUBXtqIad0TnM0zorF8tM4oEzufJY3
Jx0ihPNIXS6WdssczrIjRLkvz5MnlWpKDkgmV0sVyFD8P4DvrygaREsHCyx677rSTgUthiWk2GoW
FbaFVRiMH/ErctY0ybWhGY4gXNLg2gRMTB9NNIc/ItMkLKuBQvQ8qGNuOF9tycddXYY0dLJn9QrA
11BAUG2gBRRAoG0EIK5QuCJEsxddaG34tXcwOBvjEdXf4B7/KMqtRH/YwXQu2sFCdB2Zmqb/wrVS
Vqq0j7Oy8BqLIqqzDpwGwSc3S9rMoo1RkvoVm3wjCbXwPEAG2jvDZaumIcx5+cdC5sUoQkSe8Snq
Frx2wjdbumpu//lCBPqPLcoMpFsGScFDEnINAJQUzTin7lSPYF6n2AKbGHeoToO0URRRVyiHMG0z
6WKpouQZ/xuX2Jij1p/uLQyduRm1OwuBlHtagg4JmMybb+7IHwvqfSqJ5bhTionjmxo9WMbANAe+
rlPPHkKyoS/UlWQU8Vhj3n6KHGWo3r/ylRNrt4varZRZF1IInFu4IZwrW7QLrtnojzQWV+jGsOtP
L91JalVU2zZZRQSCSfwz3qqrCFc38qpjw4zdDUq0vinuqyMhosonXUA/t8pmPURNHeKhpHS0edtq
coxcg0yAxFOSAVHzGg04ZQcsAfSXtLMTrBuqc3ZRPZ/KKN9JfdrdDXJBRBBJMd0Cl0xDi48rLJtz
D725i/PGjYThyxLyDKnzJRcRqNJtgDUAUz0RlhlKH/Gens8Yfz6WJrIm5rYXFqFGcLSQVS3va/R3
LuYcouNNFfHQI5AjuZlaDHcX05miwcAwtGfl0+QcaaJJwu74c9sXD+QmwMhNE0uZ09Wf9IrdWQ76
QDL/bTj62LWv/vHjj4Gzn4ox0K1ig/k1L4CUWG2zL6EDpMGaL6NDoHFVNGPMxsqahepaJ6eCL05Z
sCnY1DrWoRLTO0fbAiZMpGUUVvOm2tm2dSboPkTfWhuzzeEtiYxZ4K6CEQasDjzisZb3YI4wHhoO
st6DfQzwuY39t0fkYGBSZumWVvIO5gZf/sE3uSQkyFMh0OEtASk/HjhiKQyG928M+knaOs++hL8e
541wrTcRg0ABJPTn0g7Ektx2Ym5CYsyfX9/j5j2zvI505HMtZcFGNiYwML9qimtfsy13gBk2ITwV
dxGd+5wLE344z4TU7SEqU9jiZWPkCSZxmuGwVxOq1CS1naGx0BV1HE0WByU8RgyJEir7Sc9dxRJ5
80bLBZxOvmqM6IM04Pu1lBAcb2jYikVRTXt6ATS6XP18t67wqYZeHjPAz5/BeEOqYUK43vPwCL4c
7iLdaBpH9C+meUWcgBF7Rjc2G9QcLW+ZkffSuRiOWPqWSeYLNoiLYt2krAVz5JTnZIVgF0NtMnGf
17Rh1ai47nQaSj75tvywW+cGT0upVFKAtN7AMtPNMYRr5dmr6emiPrrqKX8Tt6qW05eJderQBkVD
MFiK807iF73msN3hGlPC7Je/Hlzt8Pofd1xMS6RtuXMSXr/8nlYl3qmjuZCNuFoufywSfknjjdW9
B7KcMMD4xA4HnnS09s9iUGzocnD2ZgMGA3mz8LjplgQ3ZMVl1MLag8hKr7A58+ItuoRBWhvwWQqP
8d4A+XsU9Ld1iy8jrNU/KAJeruwwtPHu0xGjQg5BKOHXQ3rve60MGypVa6UBpI1cJROv6qrHMo4O
s6PQZ6eBDs4I0lv+W1HwNQDPtJMZq6nOK4TefmZEJbGj3JWUjOcd0quDSmZrqMSiXCIQtJUTcljt
OZKWZsPi4YRds3ZKElFQsnph3Zhdd2LCxHljwm4P7JCBMu51u+IgzUBwjXsznY3XTgNAeeN3hHdY
GpngQwty21l7i70P7fR6fsx0+n4yAWBVWGMXyzjpgFQIEWBfkUIdXWn76Y18AWYYybl2FfI9qIRA
ZbvHqLIDnty4zcFINwvgt4B74Ow8b4f/hRdhJRBgqC02iGNkMvzdaZ7t1Cd6mo2XVw0po5j9WnDC
E8dn4w70M8bHx3BncnNalosrzYfwmjy8pBsDoSRBXaj88i2XriAb5MZoyCMMud1QtJpzjU/AJzrW
rE49iNUMaCXqG4eM5aBfMRIKwS40juDkg/wOBYQ+cU4HPFrgP10oafE2F0dLoRkOlbd8dI+cmWSO
3c0TEscEnPfPeUqnVf6yGATOQNpcVR88m2xOWeMNZn3QGsfBxT/d3fLhh8f/tsunywk+qDLbDvNr
YVBS0/U8GtbSGRXspnpOsGPRXfYSzjUPxnh52J7+FRLsj1HaBvV6NdI6Tj+CtNeW08KbYLIuE5AE
535pwbEOgT77JcugcIqpwX3Es3CmzOmyDYaTSz5h2Z4dXeXOD3HeFSQtevJk5TwlndvFrx+JeFHK
6e92IsgwxUfbDx665LQLDB36UIV2xkUDb4K9cGQro4+ioExlE6qyzZx/3seGDgm4kFxMNvXwwenh
PoTm2/j/4PTPFG6SGGaJNLkyu6bBqix4dVoas8B/yWOwb7KVOA+4RCknAQBMq2IHn25AR8Co9hIi
8TiXPOOhpJ8C58fVwM+C6cKp0FzAho82orELYjopQGcotMLFzM+7Z+dkgR9t8Jnxiiyrz6hqAYIh
zeP3MGH8oC8u0wPb5AmW05Z/A0+BJTAN7wc6iFZvaFFT4KUsaIcv8JNJOhkWqkT/dyqcVFBcelJu
wB9ZkNe8j0AUA1IFtsNPNZPdCS/wR0oqNf39EOD1NGQgnLcqR3hOUiLA7ta/gD5oRSWoQODC4nXP
R8AweIhV1AFKeGzZ3y445vfy5Gl9yaGnZpEb/oEHbClklGayR1tdXQvSTQ6nMhgdsMgcH+pvtCI+
DLkF7u7NCLCiHrT4hYmxJNZPeRF9EIoCZ1R64fFYqFsJNULNl6XEGAigH3u176M+IBtkrVXoKYOs
HZoDKE40WgbVgzWPQN2bAJya0ZQVbCrspKook6cMOzL8q8j6RBsaZoZJrTmL+i+dTvPpcb5G6INJ
PjaWgrebtQ+ZWRF2rst4iBSom+2mg3adlWa5Ica63OQQRC12JcMj/3WOXp+t76rQbGocLSPL6wYf
khsPH7xZ/s7p3CvxDnbnfXzMLVeCpccoCjJGnzwLnKnq6WskEAXS2DSaaAn3dEt73OGGuQ5ByST0
pPzdkGh3pA29V6PhuaXOE3X1aifkZsm/oDzPobUbpUU7Wl+gGng8///Kr/QT4lOTBJtFlMwKyUPx
bGk6BB0MKDmUnZjSc0PH8vC6BzNp2WXwm9/64V2zcOS/ZxemKowookJK6xSAnTjgTQR2PMp9uSHj
Nby9ZD5VHLV5gm4DVPUexqQr1vyFTkwf+aYtBF3Anft7oe2USPC0Xehl5bCAwzWtHyRDwuHOQarp
xthbD8xPh7+ic1AZ8gRltj4VAUcOLL3b2WRQex9k1/RalUgwR4mqKPa7rZyHVW6vRy2P8MEzc45S
ZDL3J3vI4APjAljXEmWEeCPaCuM0eW32ABMwFidyA3TQmrOPBExYjpig8E8e5ctNikIUgynLZ6Ls
nzyXz0MtbaINrXbezl2lSPSwWoskZCwEjPMtAUiiYMlKBToLGhevG8Lu+/vDGEkMGcDsdYRvM1CL
tv+HWI/AuCpXOAYJdC6EeV6Zp4c64pqhNlazEhE9t+mWSwQ53wQu+cj+G7awueb++9jGk+43Qnq8
4rEsmouLXTo03TxcpM6rLYh19A+wngETmEK01eps8VfwQjJk6q9dJoJTnGIlSDTbHJ/28UWPchJX
xzWKMwd5eJ7B6MchTZJxN77jWREC3vRGCOtmoCn6pxhFZa32/JefL0kL2vWJG7sx0enW7eec4bPH
1Mpp6oj/f9NAZ3mVZuADE6zL/4UiYPHy7tIN3WiX4QpXZrYfiZTFe32ZoipEbZVrKFL6A5Gl3KDi
iU7yyuDD875vvTn5xek+qGuTVqYJML98XnCKN+GMFjDAKxvnO/MeDO2bhswxoa84R97iLqLRNvjV
Io+h4iKzXi+OFnXgXHRTTE/Xjtl5Uqtlrcs1ZQPRU/haNyDmtTGo3OLQasVFP9QdBgAymuTuJ1kE
jIHBCPN+KZrgCedgObn0Fc2njyfwC1e7WlBNcudtOSybUxZEJ35lW1Jjq19tVHS0vrJKz0kbaqfp
F1LM0P5xmESryiZp/HnVWVo2mZ+2I7VHZW+XlcPY/vr+RFsuA6x+C2rvI+vZc1GjFod1qhUHR4sk
PG33h2rR91ZxpGXSPx7AHS9UzjtPinUbZNmFpM9jfLWNvLu9iqfa3p5bLgLVzAaoPMLbcS+hSLGu
DHIK1lodi5XzFYsghmGHKLSiMXhxoINgnVqKqAMsI0kIXPaWqzMxf2ZmWaX7yqb6t2jjQaIkuJEB
rDTPp/ZtC4irrbB0na+BWmCCakCv7VgM6HR5CbbVUBANSCGCLi1tsjwag0JwaLJR83QKE2Qmcjjo
8CdxneHopl9I4GfyAw2IN7zWINOgtR9LYjmzZfROpvBhhNVyxX9dXJdKoUyGgSBooe7sG1SCcVFb
wD6TFhu2EZxmcdiTVE28RM1m0cnxYiG1lmnbKwjgU84nwmhZqV6Lfq1A0rRl5LZq2LfeqBO3UkB/
XWBm7qrbygYkNYpwiiesXDtR+N25g13Vy4/XphRPhSgaSKAsNcTQ4nnKezkgpwxQkyyZRlHc4BMH
l+E9NShstx8+sOOINB8ph4vg9sTCQc1+E8n0vfvXK+5feBaq+e6dHuv6av5oNzCbhL5NqZSh1fkO
ioP7pOVuPhWUhrKsnsUJt9Ba9krIvXDVkZhQUn3jVb4pUiiy5fGXvkL5ydTyFU2R8poyhSqY4i/B
+Wmm+RctH++NesNOPvSB4+vSeuPPLidjTWMOPmW27OYvsETs7/C9ggg9qu3H98aDu9A8sN7P3csn
2ksGmxxNghTyKatU/Eern6j/jWWvFl7cPGiLak+ub3sOYNs/ZgQtl4GRoJRvcmbqMX53hwh2eZeU
J0K7qvouCAemXOG8ZK3A05JKaYdhkp/iwncsfNLMBjWMRrdyaAw9chIWN1csK24KbtosuXtVtys2
BLLAuXzbghdVlOt0CaQG+u5zrtd1ZGeJ48R/8TGL4mRSMFBr46EU/OxI2N4AmIkIR8R1XH0oQZei
spaYCB+8N/11uK59xNAVWvzECIkrunzMglycjIsTGppG0RvgQMX/onkPLcS+33XTe0ie/epMmj6u
cVxsxSoIO3nOPh5dBECt53eqIIXlziRRZ4f0VO7fEZNxuPyfSXNyU/NeyaocA1i7ZROqxGoAhIn1
k0+W17ZFOkqjC2Y0Y2D+wh7Q2iCNz90NFWpuUXEjSJuNEnvWT00WM5h0Kh3kn7REh+tytn18wiCS
Rj3uIVhyLyPDfX6GOQSfX3vAJVuhmUzWIaWF+6PLwZn7/3yT0J8XxjyNyherBF1ebVrtZP0wJ71/
3/IAgMMETOczxZJ3gvgZLybKZvHIQF9JXURtskp5K/oLJsDRZfTpwFvHci/tiUQSM3sTRB/3Hrcy
/ZyHkuPIy1WrwVcqJ44iMzNj3WYymoa8qdtGUMiMkTGVpWw8Jg8kCRAoQq9HpPss6F1vAHfBnWsd
Qg41W7kxbNlJXZKbP/QtrZPndASLY+iVzAKY0elurCpXzoERuRe9H+EhWkL72HxgzuZkwoOuK0Ig
Dv4ey5fale/iDJ+6InFK/L5V6cxjz+YVjH2M0XYIHG2JSjjITkdRT2yclfb4oeAN5f8xNvathL8w
rHHv+AFoygm65Q7S9zrf7u1XAvIUc9qt1lDGaQo2HBYTvE4VVt0ulNHeUNk0e+/Nqh7A8pM30o7E
yRnvdR9e6yY2/p3zAXpRhPSESgAnGwiT6T7zDWxsSdXvZPwDIRaeuslqoi7zvbo7DmcUjWgobqZz
KcwHw8DgTYifnlgRnp6Fs4d1dDu2CghxMUODR/22WynE1CRqBT6AqaR6w7pPNJSH+LU/w58jQGvP
EZ0FBiyQvGAwT81hpGNH9gX2xWeQHJSulUWlrwN1O2JZ9uZ6Qa0PsWaXy/93eOy3ZIkJ8vmexLN7
89fuVPEAk+7xjZEGOcmTYr/SGJZxZFat/1G5+7ptKQWn8MhRofLQdVwI9SmIEBQB6037ZEn8IzXg
ZYiWT0Y/pRaYhKdlabZzD5Lpcpb2paN/E58UYz8aThAE96198UwApYE2cQKPKd6X2q5w2jywaRsP
WDJoFZ7psKRT7yp7jBg4to22bQTNbspza5XoosHzTtgB2IDloQ7iM2MapO0yt2ienku6pKzm8IPG
mc/TKuWkgyU0Y0Yo9G8od/nNYBBH356hk0Yghjpaz0a2OPLeO7VFuyePMJAmOLxfoNbbWfD7KomG
YDyTQXFqhTrFkPlRqlmH632aTYRSee/ai5ma07O+IqqjzrBTDfnxfkUS7LPOY5OaPgz8uAataW2i
VgSxEIle4IlySQi4g9N7+Ub7gp2Cy9sz58iJc1qMKcR/hFviTto2OjEjxZX3i9HSy2kjt92swwo+
ZVnuF4NVpQ6ahg9otSbIx9nWIKrlpeAzHhrZStyngCWnZnLcX9/jVEtsxdN4tVZGU6PMiOAdo33i
7SWPkJ7FRboRjod1BSZgD9SOoEbSY34F7ijVathZFh7BxepssxcALSw3XKBbqMHeCeT3mdVlagYm
yfyis8VeiW5sibpTPrQGFv8EqRI0Q3sRUvN54myFMZR6LUEAzXAi3JLC9w5rt45vO7uVOX+P0+Lk
j/fKH2fbHEEPmChz2sOzBMe6WMkyCPb43GOFcTwSMfNbfjOpyEI/dJcOrCJ5Ul4XsE/u24rT6s0h
zjvcm563ESVx3zRf89SozR3ceMzLr5UO6gVAbBOoAJy0G4dfSsQvwxV+Rr96yv17rGE+OoZaRZGu
mJKS3anFT+Sqyl4ra4edh5BFwRRIQVC1toXSYPwP5H+mdQdQ7CrrEt7A7lT/VyTVXxcbQQ+H2wQy
K/3dUqp10GrtmiA2lZz+HwkdYpdG6fYApTNbHrZb5J+Bpi/cRsYU5Aw/8JA9bYs9ucHNTRLytZq/
SRxQxli8EAlvV/ED8jH9O3Inud5CAo6cXMj0CT22WJdyWYBnW3KWIlNTXsb9+OyF3U7GwuS95NEN
c52LiUJSvStmhCqqZSQt4+oS96CZ+R3MkJ4olzlSR/MwsWSkdYjvaflLKEC9HEbOnxWVZd9+PBvd
mtOf9dpEBL3WdPyphdjk/VntZXW+bOga6PT0Fu7E2OBUr60assxRLQ0zbnqhTu1munLkzxtDWlfq
uDQxviFk3BT2Iz2oynBrN+rYTe10m1WIH3qrUQQ2KcIgRBfu7ib/oBIbHqxpFx+G29bu04DAmSp3
pInjHp5P72UDIZ5nxBrJZa0clD39u0jym0J39E4udjaUgeTFzrRppKOElGwagm5HfVflxp0a4ZdM
eX+aQmpKQLITEnc6+yYrisw8Ng1hr+xEUNNIYXXAMcaKt/7ySmOl8ybMzU8bvKhn4F2f2pytiOXN
htYVHHfn/UtZBTOwXPjOduMGrcF74db5lwu7x2dhit9yUFwFDoQaZGxNgSgA+OsE5dvcnL2zFkmv
EUU6dC0JEaXEqmJUdizf43BAlny+/HHxsx+vQei/rV0HMSyiVHTEil3QIt6G8DeaRl1LX+NUGZlD
leHMw6GL4EXADGF/+jlOrPIFLFMs/XeSwPB4yCPjqmtJCxdP3jl6lQX51fv0Bx/xwhQx2R2ZJ42J
OIEXsZ3wMydZAZsSYgeI/eGkjTQjJifc6+3TtvWOM6jXOFz/tJEaBsIfU1mkylJc5fuGzUujUhEQ
PSSerFGY/boeSKM+iFQkXoPKLgCrYR27wjLjYedgn9zthb1P933bvyIrmkczSU+SmrbiV7ScBSVk
hhp+li3LmRQwRPrAULzsVjh4t1sTyMxcT+5TYB9R7zUTgwcR87EHuzqlYT0vn13ZnGkPCwpjADqD
aG5UA/Msa98Kvb6xjMA65oNTgR3ZZr514KCRGO/8kIx5hrKterMZVA4+JLFdQ3D3GjuhKjLJ2gZC
Q7PZ3kmHZxEoFGKiQwP7T4nSa702tT+hfBLplVBXpwFgrqPEkWJAKxgXeP6+iMvVmr7+i3luoy6Q
COdfeOrbomnP1OeflHQ03NCfny6hTkk6KPELz2WqbE3PGVF4GSR5CurQdY+5a2Tgvn1pHAn9Nebf
4LZU66fW/1mmKCNA9rPQjyAbG7xNKOcMnNCo68/kuRYpBYq5fKSElaXsp3xTXSM9k9glGkAadp/m
W8Ckv8VAen8ErSkOxjjn58rhNacdbB4XI3QxvbJ/LnVQizb3p3ocgVv6D4Oe9vwio1LG2F6qs8dw
Tw0jGNF+/eIM4Wqqk/Ze/AjkxELbfWqAsgWFhLDk8t9t1n7nyNj9c7zhlrWIes/t63bfkJtvPLKU
5vzHrzRXOXwjouSP04i2CYCMmR1yOC/xsUaHj1J+e5Xg9pfdIXnj0Q1Zym+Ugxv+DuGpR6UFvqWr
adstSDLdR0ZaOX/f0zhxncdMd/QkyohOvTLK3IBoIVe9dIKKus8+hfXglvR1jR21DygDhpqOuo0I
l2hutUGJFCkAkJm8XZ81jGDR5cOpd/szDYBx7AfdJJvuLxbLX9TA2458hXE+6E1TcTS9TLIpY8S/
NhE5vOFKyWm+sNQ0vq2HoBNBoTFJ2rlCHcFy1NaEEzUoYKAKfC7uIBOjBbtrZ17TfXRH2NxAwmD4
cSadG/MjqjC/jGS6zBWswpdJW/8Py39gq5Qg5gJG9ZiF8Kik09xg6n1Ddjo8xdpH8tMK7tdjWmnw
h+zaZAK8DL0YQwuRYfBxqA/VPvRt9ZH2+xY3mivrh3rTzj0giiYzM3OYAk/QlFUaR8xn9VVjbB/o
HJQWQoSCLfm/y8trSrQJZO+1hJPqfiYVZNiCx0RraFJCG0mBv+MomBDBTbBSmB8+0VlDeYxPktBh
9j4BAYgqVoyHkELrzCXQgsgyujTfHXKLgiofNn8Mg3dKQ5rqpSLcRDvH5j4/xV/4v0ysBW/foyHH
ENPm07WxkoRJq9+ic90uEN2JRa8h1RNneoNXh7UPfJ1h/XoLCQph8dwUh9GSr0fyke9mKxrpuHH+
qwzpmbcoe1nn817EXYx7G9+toJopfjRPR4dgF+Kt85IUF40+vF4Z5Z6+NfQU6jwk6oQsJFaXmtsJ
Qgn/K8OLivGPgzQvdotweA1NYg4BKWNi9ViM0595+vN89D6CQlQUCFuKNomIYCEdmr9pTy6Ki4C1
wo0n5X8JsDIPysRpRDN5ts1XsIJ4Z2Yo8gdgxvVtzOSj1UM12kl39awQJ83Q/wIzBTbtFYqBvJFi
NCUfbnQ4gu9vF24rVatvnVBHtwzisehwjBjostYapWPkpjulDh3mRALVTnI/nqVlvpRxw3ZZlPhd
3srFB7NhYUQ4IylYYio1yszK6uESsV8VM8N0XWQjNoqAM692819ul85zy6UnZ+XOO7xMNOqC//bl
McpsE1n8ZmtVxgI/mpzNvu3csEmU2Nb1J0CSffBAPi8mVIUFBMzkgBWH7e1U+BJcfcY1hGhR1YtF
mrY4lpAKWspGhN1DU6r7PtHjTpq2klC/H0bae6XUQY4WQLKxJwGffwo1FaPutlV8LhEKVmIEQ353
HqPeINhLNZSbLNbnCcdLL9OyMEfM7NYducI0nHKP//O6hb8MtBUPOGxC3Q78Wk1EEEcsAvkjf+c0
QNh/5NnRwhjc7q90rkC+iNEuWZKeLP2l2c74DdRvvB9luRWZkb0gsIXRsXk3oTSuSeNNw+uFXyQ0
GY0bk/ieXIf9OedjdoPmG90eAc84UHtMZps2so/dinUT1nZ6nL39ZckmRY0YC9b8YJqDa/CCn8qH
AcRSySAyckXhAYufCAzubz7Tx4pjNAmScvTuJOHxueG01bl1b/yfv5wAfoRB/WINzU1T30UMl7UZ
BFcpW0bx7uocd6zJwnaX4ojl/+rAdiHRhtlK4m/WH1BrFN3+mcbIjKR/JBo8FrCcBGS9JowOC5Og
LkAn7t3SRwq6InJAeskHSc75xhtP3reVo5Bx7730pVVLDZeTs2+EcIpQ1XST8fGAEduOYlRrpRez
Ylisy8XiFVB1OWHg/CetWDNTjW+si76ZhlYgV/QTRqNm/Eqg15obZXTqZ5P3TQaM6EIWvPE1Y02d
atWW9vjcdc0YiUxhWI/JHpyMgNKetKfh8IbvTxH83QocZt4mrU0BHjSesbaQ/SV64TfTMVpknGRl
sBi4I0PIR13zMqP7hdajdgZP9NBSzEaEuxD9Tlnir7ZX0J34PsQLnAYnqy1arLawpH1abL3xZEph
qFSFGa7Z1+2dKXMDCfOI6kHVceaWPr6GAapeed2CyQw8rgZsoXQ4DhWTArJnC3o+IpQAxDu7j3eQ
raokM0BtTrlnTn332swYcnHi+t+4CiBqQ3zuQaYkMbYHxV3Yrq36FGGKERnpBiQY5/iFXdZWWiZV
R1dqk+zIhajNlz0+SBoLaDcd0m/VwobTBuzjKmAINIRcJySHMTJQJS7yVOShHglJjo05Nqy4gzIo
j3YEwK0sUJM9VimMTvRGgHgbRZJ2glanL3nBSMQVVwYbpGf5CAefQRLd7xzeiV7TYo3L4/lX4Eon
6w+7SUDwbwK8vulDJnTgW8WJ6fd4c78PyqiIgzJdCN33Ho/EDUfd3Jo5I3lTNRmAVWBl/Hwa0Iqm
XBdYkCD3zW7jSpy0CDDOfV4j/eM/vPcHz2IF/5ry3y1uurq0fkfwNx8m5QDfqJoa0wNxHk/Yyklc
/sy2NKwdnxuKUiHEdzNV+O0vK97/rzDEoi99sViZ/QjNxKyjXWkZuP2nZ5fAOtVncVWuG+6l8WHh
Z2bVyBcOKsfCDRjxOKodMb0JoqXZf0ABG/+j3C+3Tc725NomXs2MrxANejVYyOZ/0wwAOj7Nij75
A6IL50GZDL5X1BrVR64hZN/uzaNVDQ+209iPvtCjQB0SnO991oRj1OX41TSmGM8NpDjaiIkkY3DB
4gH7i/EuBSvtFHypuzqEQ0JD+hK8Xgy/0yb0VRfXbFZjjs2keG8X1FL+uM0g97aKhFt+J1wkXxNx
n8q2PKpMl/qh1pmN4tqZpbRxD8G324b0nYe4Wvvymdvrs6xFCt9QH+401nLsNm+6DZeXl9VZ2MIb
b7Pd/7y5881qBWaXAQarMpGCElgpiof6LbgmW6DWLF/FGeAq5I2+EsWW4C7kFwIgfvyi6Ky2rQXD
zcidTUc2lukrg+Ttq85aoR6+rqiryu4W/JaERvYa+Pi0h9nLsPYzO6EE5FR5FdIC2Ez/BacEsyOt
rMhY9QhRzTY3U7cvEp89fgUftOalhg5i+YKsPqoxKI89dRNfHui3p4hAeMqICtw+z1zqXxJtFv8M
TovmWbneq2uOqlTQ6sOgdY7kM/k59e5vsaA9TclAx6wLpM1iTz7J4Cxz8FIYGP1kFc4NSZopaWIE
6SpWXNw1iTb+D80f4xQCPA+QGrspgOTWDJsJxjf2SWJAd5EoRerUoXRwVJ97CI+krF8g1GyQT11T
m9rz923EMMYfy0Za0DeiIJdB7B8+YP8BUCy+1fKfF6YvQhmEQqk1zFgjmX0HHvFR7/Whxjuqua9V
N1GoAGwGcFlpjQ8ly3Wlqb6t7HSsEgHfi1EGybWATzLzLo3eliSIgozYbupjUm0nCW9pM29vXHbi
aN9AKotLMRp/XF8UQ+FSDDZW+RbRM2Wp07oLG61X3EaQzMytT2cYOJrjKKWbQzDLK8JdNcbC3eua
EOOwvWRkgD3GxVnUm0mbIvlTW2Eve3CbtD28J8ltTw7oiNwv/szmYWpzzgX94S8JvP0Rt/AHZAuc
fWu1OTCugoW0SxXw5v9FpCV4r1doFVqXBz/OKarpdszS9gPaLvrcU8ow+FdJacLSOBC37zqCeorg
xBYuajvp+mu62boPcTSoPtJSeIHmPC4qKRsiF3BBl8Kv6r4sh1f4q6nugHBpnuND6JIv4W4O0sxH
8RJGubyey8e9yNotzLzhdt1YwA0pH9ORyb/W0J24K12rKwsUjRkElwTreANz0fJFT7Kc4oUqo/ke
0xdafnAcDpXqWJqlJ2Z+z4HxsTSM4Vpaz+awo7OOxOJTzBOXVVbszY2ogi/b8Au3tKVhronfv/ty
7f5yUJ47WuNlpu8dCzHeB5DFcO1BnlgqlbduqWhvzYac89/i6AlrYdgXYw1T+tYlH00N+ZLKjL28
4ai0/wSEKVWIPJPjYpm92gkgYgD3c0JFN2rD7d/6cd68LQxpG6lFbFU9reQzAOSZmvV5C6Ll2fRJ
fs8oYMPxT6WOs7j30sfnV6GpGgioDTUd211u/eaSyboDaLcfc4D6hzadd7/gK8RW60qIS297fUKP
cUUczOmIa5Q1XSuV5RYwxLWW3QNb4hq3M9KhPlsQp91rK6EnbmHuQyrYP0ygLRQysqeiQM0v15UC
0KdmetZaeFuLCnq0qWLE34HGepa12I63cAoF6sROS/jWuJsZHMa2ZN9InTRfjjoq6TirvdRuvhIs
nRtObxXhUdPgIr0ZZJCFb4HbODmIVmtoanKX3YIMFJCqHwxQU8mouRVQTSLGJTmp6aqvs9eVczR6
YfLxBq+xYifTWjZ+GDh9qfCEeukr9qlR5sd0VfYTCMEBaXkQUIPdzuh+T3j8fiwEltOISwihWMlt
EVur1ZU8wTNl8M1Yq4ceaNKL5ELF8MFPWz3h7q3MK+XElphjlu9llceDTbRTWLAnGod0802G3jjz
GclomZAjVWjRPDngu4qarDMC5zF9KzGVL5WQyprRwoigaIqqvQLrohw4JZDP2/u/HRjeK4EouNV4
4wcOMGokgn3Ri6FWa2MydqjR2fwF0V1LA3aX5e5otM/48qAfNqpltl5zaY3lq/PnMmWCeUOxsOyx
i11N8kIt1lh0K2podRP6dBuSpcCNhskfXokzKKLIC/gYhdfqOY6JfhpFid0tID1//+YZcq1hXn9L
Fme03A2oZpoqqJzeVKecTj22u3E/uewhAbZnkmVPqkDtlJRTYtIDvZo7QiqlYy5tphgDv7EZvmTk
ExL4T8r4qn2/Tp64kaWT+IvLaCt3k6px8t8FhRpWTlT0ecl7zVbv1Cnaooj0rFxKD0XnlICA4mr8
PrHAwjztbztq4tzrJxLd3jRboYUeT+u1W3d3Deeq7TgiRvo9scfIRO41NnD/0Y7ctt03TYdaOPkK
bykc//Bvb2UtpiYFxguai1/sAJsC+KSuc96EvEnG4hXzbj/RUbXCZfn6DUbfIAOEKWuZoK51zaxe
T7R6CpUTQ2V5SEZ2ty633B667u1ZogmXrTiVuJdR+2V0Wu42IR+OXvGQRHe7DZQXUw8NFcp4U0Q1
YqgBs2DnEEeXfD61oj184vZJog+Od18Ec7mcr5XnXqtoexuYHfuhEmBc+fq+qgsBFGvPB84Z1xHc
eNMvCwnJbJkDnSUuc/LfFVXG6ewojVX02OhTKtlmhMphNDGlthNGDkSZZhBqAxEKpNPxDoBtNAKU
l5eTziVnHyXnL+nhUCzykQ2U2Vpkb23s8gldegECzLM8tVPGFwNMi1gHeDKnBX67fBCxf4GEp4mv
/DYj+2SPRc73UekyJIA8e4WQIwIGApbp9QQcHMRbOfTkuL6DFu3tKg0HNpwfpRwqtcKGRzquMoxc
o2stTMHAkuJ3b+A9W9WgoldQvqJRU+L8bVrdzsT0GY0dVTfWT/UDH2zRM9Z0Go+oEaWTn/zz2YAh
hwfSwraKZ3nVb5D0adY53SSxG5l+uKY4BP5xznNehQIIxkV96etCyS7R8wEsQ2X7JWGBEnom2Q9w
YmPZcbZ9NSMV1vXL9vIBk4Zv+PKb0XP2v9b1D+GD84xxfuxfATB35NmRkStds4Qd1wH/k4I5vLCd
LX+in/w2HT484g4GgjsevX/L7/+ND1uVtqs8EMsPlktcpOI02iPCC1RPgcmH9WV56Snr0+0py6wz
CXqZNp16+KmPZI6LxkpHey92QE5QafPv9y63KJlhmGO/Ce+1wK46oXpJDYE/44vU+kLO6HlhuSz2
U44BzxgAUDMTE98VRBilbeEM/Mz30QYuw8IOCz5uPeOfkIq2621zT8WrI8razQkNWFdnrbKImu7T
GD62Pvwyh6mYMIEYZ8ZxWGJyfXbahxfCMtyCOpixjsdKEF6gdMgsKlLC16TlxoP67U35ElIcl2gr
KwYBXSU992amIi7qkiF+JFBonSjil84nuNYrNoNgBN22DNSrm7GmllTshgbLJKRgNDN+MV8R7sRl
xkDTYKXNpLPgTU15qrKWTs8Jkz195pc2FG6w1OmUuS3fu2TApYab4k2SLfCER1dE+skatiICvwvL
PXHyiQK0RKWcnxiM5mhybd+hxHmMRGsLTpfAIVZLbxJfX38KlpmnR7hgpyqx/B0F6jTGG+vqldnY
hrKmFW0vTs8kv0reP0GmlOEv4VGneh3GG9ad4AmYWk2VTKxS9M9ayo9+5812FxptfzplJMbTULqk
Ankgx0VdT9R3yleku4g4u09y5tXEkg59Eo6uNF9PUcoMZk2lchp9ocbOV8tdSPsytxTbv6zofw0t
1o7hRB0foo69lVNMcvUiWqlm9v5wjmyQQC06hXaqkyF69uje6p8s+FfhVzIJIdQJxZmflq6B4FoM
4pe/KbIvCu7CC4APUx4X+Vd20ScK8TE5sHozbwWTqiPk71A6IRuNsGVM2QdreqJqIIXyEpzLJ6WE
TmMQbFOrJFb9LtK7JrCsKD3EfYLogqy12jrkP5jd/uvsXBwo9He5hGMa2b0YUwg/KmwKuf+4dCQV
6GsQrlQDYxPne07QL7EIYhteUbjSLWETI0MxcrZ1gYowiz8ABrMwsRjohoUozWGRRR2iXqLFr6ke
FyGAIhOP3cjhCsFNYCjLNZq68Vt+s5FAW/Mh1EaCzog1lGaF/o3q+eWzz1KJBnZtqbAIZCu+I7bE
fxMu6LqmrcwnxWPeM/wNJQeApz1uQ7LswMdNJmK1N6MDetwdhgB40knj2L3wNF+LqHDlAAAf3yix
2PpxFW3r0UQnu/lsdbVGuI5JZKZ/JR70vshRmCx2+mT4narja7EB0frwPy8fiR04Aa4PxdK9j2VL
7snBsWfieFTV/sNpkIy3LYEYQ4DqOU+7c7QfvriIXKGRDqZyTUQjbHfxmuM6rHfhVlr4T+ODCW7U
D2k/3EET2yMA9BsBD8eAl+z/9bNMI6MLW0kYW/Dl6jUwPlvaVBFX3eQDPHnxRx55c5OrqCLkmWtg
PsdpFK3FnRtk0zMyCMNzt3vpWufeS4gn4mtv9KTs3tOcGIYRGaa5/+hVQ92gtTQV/SK22eqgI7lc
4BhoQ9CYuF6pbh1/qFnhDutBa2S9ekr2Q/rrbpcY4YYCO0cstD0xwIPh8jrPwRBtFY0Am4bf2S+g
DBKPP1KFBkFyae21sJsqeBD4bHoIIQjcaybvJmeU3IKHTxW0ewpHQv/4NO1SKPkCsGfyxYVcLlFF
yqNH4aMsp7y3W5sOIeBuCH9HfIT9Ztw6+zPoEH204U2iCTuXcmuNBFxsF2XhpLt6WWD6WJymHrer
hm5luFgO5CM6XEJ3MNZsolxN4MSE2P9wQq20lvDlZjw1HBUk+6yDdoabjpnRlCoHBmGIAJl0n8Xa
6JSKF3S+CucdxTNzo2cJ6W8gF2n6TvXDMLmjpyZGNWGC+O84ClX2abtA3LgRlWBl7eU3+pUHdPZ0
fEVftplDWU/oLxDLOYa6OKOqBW0hT+/RfSZn11NW0WrSJcloIX5OADTfAO56rIfTJHsuD4bLyzy6
44jWN5FyuTnnurVrTHrfewOimXswhaP0nUeilagwaUn0FjOFvkogF+tIRauTiaU7tbfydrba4mQI
hjqKSFmnZUF76eaSY3J9HV4BIL0RGV9L7WeDTGMEytLKj51O9hrqtn3mqqjDe7VZLildFm+DFGky
GEk9e5ndIzC97TV1EHEwCIWSsFuHfISzI/cdjkO9ehFLS/foVxZV/lugDlZvvGVDmXGpCBVMQWqj
cutyJfOVPKV1kX6N9xMkgB2kdE2MuqjP7lqlR6HoWqZC0cw0xXaGRgDIUFlYNVPTqiJqbdG/4zti
/azQT8QLvO7HzE8nNjhNrC7HCc9cL0wcWBajhGc76SPE9ECj0udEZyXfTJjjOsq1Gm2jrQo6Li4N
FgHOKs1zkmuMPujnonY0rfs1XIfhNb2A40tG53eXjwI3VnU7jG669kerk9PO66UeTU6hqicKt3+s
XftR59OziWLJef0JwGVFmiCLt6R8Qes0/V/0P+FUM6XRl0mAyXLJtJxKY/PWDIIaAMTKuTFekzXW
8BqhqbY41qOcz6ZTAqGMJfAz7mUKCgDZaRlpVYD2u78x35o2eNJ6F7T66yFwObRpqECs8Q4uRddx
vGYoiaDzT470KH0e9aV+uidvKgNHmJB7sUp3+7520Yac3ywZEVD2ihhnQN1kqXHVcI7EwZbyCY0M
HlhweklIh+RoN3x3Kb0YNSyZKmpX6o4lUl5nOUwRM3Ug0jwjdWf0c3vHxomEKQWEtIab+WHjqB5b
oY7VO/OGmxZZPYRXJGIDfZkp0W6sjU/8a/2/5Bo93ds2b6xmQ0KZBQj5s2mnFAVsxotzTVgHiXHq
wse7uxpB+E1+T1nSvy1+uXLptndOiR0+lfRBrytubIZXCb1MQSe3jo/A1iCvOgbU8gJ7OumAl+nX
mjUaK2rx3QVHvkK/Di8yvzUjXq1OckWIPslk7oFVV4ZQ2dYCvCX3s/4uaxi/t1oudTM00/VokYi7
eoar2RUbM/ZJ53suRWGH/PXFzig58zkkjefFNfrncG1EAxp5WhIZw2cZTBZQQYR9bai7KhxcTXRG
KIxePGwRD0N09oawN+rErdPGyCp/OVlLKywfAbsEyjNDoA9yffEqOKBLHd7h/AUkddQXV0nOWS+8
pSBhM6T9ig2juZ5P6V4oXkRCR/wtIcS+RappD3MPiTPcwnkWEjzwSuTE19PlFRghqVpqq6PgD0jN
UoeVc59PHdfR/ED1w5j+fpoLX9CtCi+mdSYZ4J83L8UljAZZtHmo258DomG1+la0QX1k8dWokgZK
bWOiZEqNvdUTeMKVmZahqpncf+dFj+ZVhaWq+xfes9Leemaw7zyn11DldMJ+Ij0JxZv3YG2+LLvE
wClBNoR2vTF5tJuPAuvUFgZ29meHjcRIY5LhsFhf+uRVALToxeSkNi2KSmpYA46thGesdu4Vi/xR
4YW/oiYeg69XjD7SUmd+1rQ2znKscIOcNDX+xsAkSzlUCjOwmUBoAF/cF+mB08C9zpVluFFD8seX
ksOjG7dE8exFyQCBL3Lklyh0xDCEL5Il1oaQw8sT2a8PVMbNQ2c7eBs7EC8qehMDTXpR9A/Iy/1b
ujHVMyvnaHTsQp7gcewtZP9xrlXWMd9KrqMe9hj/zckEmZw24cP8LhleHfeGacmdsxlk6n3Bs20V
fDc1OPP9XuM2slSQ7IvitFunzwADVbX8I+zvdDcaPiY1FAkdMhXTRu86t/NEp7iTenRX5F1sXdxm
3L/1F111D/FI5zmJckjHPV3KJkSUmFDTwo0pP9QKGeBqN2iNLqEo76tWeWRyhjTctOyyjH21y3lE
QEoZRYH+sfIbz0mKFx7EeI4w+4Pf79NqJRH1VGOYvq7JNaqXR3qy2+FC3o4bpmmYeM++JuWuvC/f
zOvWyIO4H3muY7rC0ixnQFuH05/lKl9REkPO+CInwfzlvd8Skm3LgpLLOIdj9tOfp9auI3LcoDrV
MahLfLhVGLeMWf2Q3/JpyoIULuTHGvkojUVthtmdQfrlCmlitdrbfyOH+K3J+J7RuUrYX/sMwtf2
pk1cbKHBSqnSYu8Sb38wJvwClTWvsAjIuqwNF8qNraXWQWdJkHbKlqCUX5yIgC0jXb+NTXgQEeJQ
MZN8mD0cblnYK2zahF2L//XOqBPhfGNAy8RJCWAVTiclEut4qeKhFscVOE6UceiloRR2LRZEJMcY
U/+jtBI2aIdAjb9U6rw0N3/I9vL/LM2+g8t0WZ7jB7LJcRPks5CAf6RUf2BQNmHPEZ8Tg777Knxf
wwWw7H+csIGvRMG6GlByBfecEILO//iGjXpG0Cr3IhjNeeJyWKOmntPVZMFZrtDVOi6UyPz2xFt7
mA40pJwwKwRrORWOw+YKK2uE9d4wKKLlrI1/UNCFgySlshwGfgy+IDTJcI/SxX4+keqmnS+M1gHV
j/rL1UEbjPDqfAjlDSFQ1vMVm/hTaYNfRP96qgjsMmTEF4FZPSlWOEl+dAz54UKBS173BdhtXBlJ
nreQ7MarPqO63B8ReNmLM/yHwBscQifbV22JMwsDoljAn3Tt02JJmsSc4iwZuJCqMgOybCvf4lBv
SjiNbyg9vGc5AON+DnUgB+WyHoS1I2zhby1X34eo/q0sdzFpWtf/44uku6Nt34UrBEj95rGAKfh6
CYuL+WAVPV85QaGjou/sen7Q6ShOnwXSG1sqxt+KLyFqHVV1JiSNZ6sXdtKnHQosMGKF5roqSC22
0ZtGyCxbsmKxl51lehrt8xonOkLLAfXo77BvTN3cDxxGyaXI6O+53BhFnq82DuY8/WPzKC0D9EsX
m78hHIeIkS/iE5wfZD+weoXjLXY6TraXFWwyL+wQrD9waKuvFYqGL6UZs61Oxg5TceV8/7c7FJCw
klPm5QY5meT6ObjNCt02wlK9e9d7jD5af4XEASmhlWy9FiNOWXT//lbK34pTLM15L0YlUyU1ykOp
P+A78oez4/m8JQqtY1I1k7Vzs0SLPcXvxGzH4xdfkGx/K+uT/AQZDjTx6d3yD3xbT4j4GNPF2KMd
6yPj92WVKZzuzOV/yQbyq0uo4d9S19yKLWkyCYjlEfSv7m1Rn6cjOzIakMPpmytpHYWNMeI2QXkz
kNJL3is3cmpevszyvFJIe3aumyMvVS55RxawMp1cUOBDl82Eotv0Y975qDoEP2YWIBascpxi8Nm1
+JxbSLZHp9tFnAVdq0wDt7zkOg39/OeuVrBFiw3iLPkL34N9Q9Vao5KPHzxu5HsPe9NwsW7j3UJF
hk/O9H1Fbmgwt3AX8YMUjhES9mRZA4jHj3U+jhFzgSDpShisipWo1Rrg/rvTjH/iot9X+cocSDrW
HsxnOpPn9okqAHg5fixBFAU+X3fcCCBROJBuCuJDR4MjFZOV/I3xsnF/yL1YUXdvGSHPrq7va7fF
wCLm+Ejx/m5XrepaQ1F/6rbvLasn/W1QKJ8JQGXIYCDknrYqqPsi/a3k7HIYNPNTg+2RR6adUZuO
o4l9b01hrm3boYZYkLbEbYFeywyr11ypHxIUIQEByA/g1/DhEKGbtZO6ThszeyytThkPxLqwVXax
mzY0qXg9bR27jZNBbXG2t72FYCgLLuI+dHT02NxhiEryaIHx8HQXfQAJ0MRRxhqj4wGNHTZCMG3q
PqPaxdqB36erB3QsGwdfpPny3gp4DqBI083D++p1s06i41xWzSfds/aps3cqW5HhoRp3cuzlewGG
wkz6hH3Y2SkvLxduzShp0yfAo6v0/hMpf1FczfC6feBIZKVVcxYs32L/F/UUAu7PpMwdRUtR370I
Y6kRuMjSIod9R1cMo6SOMfYk3oJlfmi0BpjnlD5zOBQnYAvIrO1eCYncTuUUNCz6ZxZ/8MUVIsmi
9VXKC9wSfUkqIy5NsmNJnX/aXhEgaaqpf/eFZmRnvig4CtIKrvc0SII2CaM74KAIz1GSu9WuzMu+
SGLTFVlnT1++v+zS/YbOnTZGF6N42IVSHOEmOBUFHxkxQyTcrZ4o9jXI9Ft33gEVSq29oPfNrxLa
x2TxXGjEu1Pn8rbqJEyHDs4X8xkDKaz+mGfH5KwweHvLD76HMw4WFwl9xMTZK7kwGbPy+cjJYf4q
+In8dkUmrSc32QfX4Y7BSFM7iKt2W7VB+k5qmO181eO6XeaGmp9pFXoZpCLhUbMJEKID+/T9fpKx
9LLejSRhB8OQMWocgsFq8y38gS857ucyqwapriVeZOtxVFlzquEOv36/jlVPhNY60dLZprNZzVwU
UmocWcTjPFvCz93ARM6gBtKuwXV6+f6XnVs63RdRjUouAjVvMKyJiOiThcXwIxXezJBJjDKP5jt0
KqnmnTHniw60X3tgdGCGavTjeDYZhRW0jzzLwmvaleqsjfDJ3p/w7f8oGxrKMDLcrvX35i6i+2js
CdtFZoAIsB4097VVUPT3nHKvTb1oL4RNzcNCmH7eNplh65XoWwevv1Av6V3JrzF7fng0/6IJiU04
mYVzUcH3CPAtm9tvKBXYLozQGawgarnSGtf6xHD4Uu+hacW2alHM1ihuENgc2zw5+7dtQy+HTv08
H2Zkm2N+MvZwB+nkXhY4TuUqdtvu6LzD9p/VHG6f6Jw6GqfTlybw/YRE4EuexzeR1DVrwyj+FGoT
n6NDBWYp80eGwzARZFHGWiZaqMUeNMHNcUhIXVbn3ULDTx0xMXRii2GJgTIHQDL1ZT2K11t9H+DF
HQSVy2nSov9lU8vYKyrf0WN2/kOJ4Me7HOvl6K6ijqYCd9M+iBhodKDVrMNzjK251nmRaWpRqqPH
KZKR4msrZBY/IMsNkxGhdLbxTYNgcJX/0u0H+G+RLY/UcRVE/Jr+9Yu3onSSgQI4DYTdXTDlCGDZ
wy9dDXmNabxQXpnOFD0J6DNKjUn0N6P2BKAH9ouTxgA8SvPdPoSQlIfgcmokWYF4tXstSo41ens7
6Jt1Gdh2GyOnB0kLqwxUWKkpl23ACSmM6iG+BUXXNxCayPyBHbLDqIgnK2kT5Pj4NPazK2pfTnuR
r4xELZQPMyYa/2A+HUzHFE7bWf3ZKCuMUXy5oORdRR4v+MZZECVOTLHKF5RJ6jQ2SsUUg8E6IN5d
kN7UWz24eXwUb8m+sNx32PZtip33vLW7qaIF02CJ74s5H91ZLWqhTeRR8Py5F4dNwmRkW0bXgN83
CTOzdLE/TVA7zMXqt9q1FII+ciRLqP2LzW85crm7TnVIvjN3ltZ1MxZNC9/jzNdRF1mTdE3tQ0fO
mR6MHJCxaAFbRtw1cxAVmv8NOouVs3x+hBKC2pSWcTJzbXDSIwRSmPIb+iWDwkkfphC/w0QO/H0L
KOuidCbAXjAZ8R2DY7slHI1PlGxSyVaYRg1NzGfbY7V+/A8INp54KbZtaWvvVYuZr0Mkfw8N5HX8
WC/kHgvN1u+38nRj4mMJTpHYQ+gmZjCnLdWbBdtjzyJnvKYC6zleHdmWzoP8k1vfLPdP66VmXVqF
bUr/q2K3gKDd2HpyyouMOeNGHu8Pd2KT21tapXICl8Q2cGNL/eqAiM1AeAYSt70iQJlUSADZiN37
TkspO99xcJA4/WIbvKG1quSVlQPYubbnz3d+f7rF7tA6DcZ7pviylokAsIZFL/1KOjZnJg0WQZOV
TxTkMwI63buPCTfYyUnYaiFyBIbbPJaH4m9Ot9Vb1aw4PJiWeUxnqRZU8DIWBIJAozPrfvaMjK7/
gz5aDbfWI7ErgeIR3OrGbu7V2y1i+7kPgVQjQD8UGHUEQkcYehoPKicTzq1i1pacEkSYyqGVrSh7
UeRSGTb3h4piwAI+pUnXy7yIGpbVlYwz1X8trui/aIlfHQbDFe+rat7Yws4ovXyOF92A2P05a4kH
WHcPKZavrMEZwKZkCKN6wOF2n06ofPV736MEtnPF56GLYUMroPwMKBPn7f/b/eDjkGYN/nA0aaCh
qGpZRXHfUM9tE2OaZ0aIfqe1Zx+dUJVaFEBkjXlnrFDDgCbSf/oF+TFR/NLCmkHpWQjLhywF/Vj1
/Zrol+cevu+F9JkUEzbmxdGjAanPEV+B8Z+rZgB8cQk2ZbjHh9hmtrCA4FkW2mg+Kg+JExx0VI8I
Jyj2/JzUGshrhtF5Vtd1lsHkOdwfZ+l3lJrnWxuoWvMq5orO0vfzazvwubWF7cCEOZTSXLqcwbzm
bLP+42+v/b9dxDTkLPkdemeT1u4MgrU3QYvgjVo2gfWA09zU7Ve2pVwFERLF8le5sORBDUKbOMhQ
CYj7tgDKm/5P4po+y1nEn2uJios4s0vbchKstd0QHdnybjSxo0QnPJ5D8NgIAG1ZtIGb2oG7Kh+k
roBdI2xKuvyZlg/8Gy9RFTt8GANIe7Rc5gDTbZVZEtlDdWSfUE/n0uCFa9/IB/3bjQ5FJHXFGXt2
QfgmFxl6KUdQxgwTJWN4Jr+yrO8zTw83yEVGlSvjDz2EiXflMcvrPRznV9eDeWRQmXgZ1e3oc4xF
9NNRG8GmJHlPImU9dHXyqMf/o5gVIeCPsx4GF9QxVWvTHKI59H2zjSsxNDb831A6s9P8NyLbVXlf
vkqvegCXMD5dbbNHwY/99aoCWdQ3z6wjHC1D9n2w3dSS7vbsDqoZCcWCGFN4DIvJbvTpkyWvKDI3
qb0/GpmbR4pYnDf4t4GXiFsyneI9CeNUowPRy387QDopU/b2trKVdnoAszmdzTgUSLQ3ZtCbTeBt
AXvqaznCyXB5kMScGlW5XiDZMo/iCzvmdFCOHiqyuaskKA/7J690/rOf0L20wDZGZWBYntGMijj/
B0wAGyoza2HWIRPQ5KjPlRzBQ+ppJ1dKeWORtjVnR5luhbO4jf9pHT1hZovpV4jveRRT0FxOCZdw
BomgtEfOf7wj2ENK8w2xvDf2wmYixwfWIVcBjUXLKu5tpA2UfDV6gVbEs9ISCH/CKGPQXybxbL+4
Ih1EY9/22ebAg9IZUujzUdup0HHjwso4850mQ34qt5Bz+0PA7Vze3H2G8n13dCmuhm1dx+Ge9lsG
qCtzDiv6bxdMviy+zXgQKw/+lqLhLYj5l2T3N79445SL2CEdZsEMqwFQzwRwUGyrGJvP0vuVGtzC
8jeQ205oLMm+btPGW93hAJ8dyreobgVEzB2R2e9aVbIn0899F/fFcohLUU/HqHthY8tvgNA3LxzK
MuGXqQCjz70r89XvZ9gz28754oY2IBQViYOPLn1tCagF9qXNBOvkuuvBYP50NjV+YCxCP/VQxgKI
c49Se9RYFzuYpMEby1cFMLixTWXjov9737lTijxMBhRjTHJ9bsrybBV8VQrHRZ9n/swA7RL/6Wr/
10b/AxqElMPT+nzsZyt58e9iwSnp96+zkIW8rnjml6SxhGVtlFvoA1L67ZldjE+QmKyScbvQ0c18
1hlZwHBWqqmNSXggFw/gQASA5MQLEQxVE8gFbN/+gYgknYmPtvyDbLx3uSGQGr5AxzJu3XWrDOdn
8faxXwGQrwdAcX0m6xfQiKaCFix+moXX/Kx8zg0JGb/oRp/QjHFZ42/y8q/bNBCdDkPv3Kg8YL40
j4qJhPELzSb95RtkMKrcGT48BjjMHd8p2fN/pbiOmYA3U4AciYV0eovuVwLA8tZJOdiFJt+s7Gk5
9fJVO9WTKRes4jrU586/cFjcnjHaJcch/S5f2jcmBN8+i7F6zgSugQ70phjA8SPMBWENgLN4oQo3
cLOyv1LleC3sIooGzAPWTh1RieY6EKg09oDkqjaZn1XV6LlpWjQWFfStLxdZaYhVxuiDNiHSCH04
WvxfGXdHltTfWpDeh6F+s05fSaLoW60l0Qobc0c1gK4JLf3ZLpHdmMzrsAfm/gv4+lSwcKHqDZFH
Mrs+Q1UjE/OX5S83Wclhe18+GAKG6TNIsc+RUxZSre8de1/k6aAyHgYtSykgqLs7Ygi97ZXwzooJ
PktOQ8B/Lsdc4ex+hCQW9sNf0whzH9hM32U0dQ9TRev1+zb6l7CQzGwT8XObzGPVSoJeELNJhtLl
QjLq1DkSOyLiTuhJAt+dFlZxZ2TztIQ6u8BqTTX4Jy/hptSPNJYInjTg0zRkv+I3D96lzH6rQvv2
pVjk8qD5rQa9uEebh1jGPFXSV4OsK5WU0G7yZe1e+ghk5TNDs3I8APVJYBQCTGOcn4Sk9ubeQl/Y
ZyRBy39vSFy0HTr/P7V9ceUukkjcxfICpRfvsOiW86jVndT9R+5sDyl1d6bWb1eSssME31YU9AlQ
VFi0Y2Rx/0xy2H+ypdaPQn532XjsmdjojLJu86ncdQqJdhUMZ0XNSNGYWh6lEEFbb1fCHAb8iiq8
vxat84XUeiwMNS8Ov5oZ9BM2ScMl5E58bGoU14ojDOlLmLvB2OhrOGuOFL0tHUWivn1112sZdP/t
kd6eZ4NabtlsF6Na+3usQcDrNkcxa7/trET8LWAj6FdZYh4PxHkfRvyqMksjBZn8Mgx222zeNfiD
WeKhGJzpLruX87FSdL0Wp5SsenBX/o1b1btkvCUOJq6EovVhSHO81kwFfkhWl1T0t+Xl/I1sGKH3
9gvwFEcYZsyiF7sk0EDBS7cxPcebMVTUVvJWOkBerHHuBUynpqhpdSOASFBxMZjK+HKuFLHudJ+G
1XHclKL60ZUsLZs411W+B27igJR0MlnOqYKuPPIo5kNfYM6IQdpzjqwu2u8/AJyo16HNVTKbkjqk
khbInrlXK0wKtsZclthfntYFK8A55vRrJl7S8xz2vWxXKf1CCJhZzMqkw+Rc31cH9/2gqZj99Sdz
OqLshh+F/ozS2HCvWM+mcVn1EfGTci0HI/K5J52o9J32QlZ/1pYLyO5R5QKN3k7K6NvdNXwfsraX
LiQgC8yY/bUMBwM6P7/g+q+vRlITMgCrwkT5si+DxBqvLcPLhANpjzcN0UrOIAgJgdBCym+HTK3e
2o5AIzjngJOe19meiDabdGoM2ybUMu2s6J5ADzmZMsBzk0TquLsx1OgoIrPnwyo7yr2kzLoMisNQ
g+SbtINIk5avIfSFfg4IsOQRkQAEqlZHWAbI5ELJ1RjSmtY1Hrt4B6p4SoWWx/tS+I9Ro+Zj4af0
G7aC9qBZEHuL917pgKWyEeQQqBq40yH262AQctaKJER/MuNXaj7ZZm4h+gY+HorIiM6SaInYxXTX
rgh2S0PmE2ob+kMshl9OMyJEjc+XXQ6bO0b1oLJvIELXN6X3R5ZbPw0JYBV1SiH0Ev+jn0M1zByp
9pmGlb8FypPVgcEp7npSts8Nce5anr++mug8MmA5wpW79D2sE6cBK4tuB7rZrZhgoY0h/N8hj4IU
ZXz/A1tSSkkFtGhiKNs4lknsa+S4jTRlQeKIQ43qK60zYFM8AqtfB4N/sb2qHQEuwHsTB6sQCBby
Sb/mT/WNw4Y+TWY4ivVsHox78CzqZT261IPqy44r20WyUwDqdyF70FsXz+k2wYZmJugBq3kpLPHQ
Vggm0+ZF8ummO0HXwB+HLrEkKJVVQkEMZ6LkYckft7nFMVl1qtNulrQJdskzzLeg6zk/1qRBO2wk
6DpIgWsU0fzq6aoKQ1N1LlnNlH3t9bmvXtafuVb7VLdQ2fsYcizzPoE32TLJYcv+6aA/y0Ldh8dJ
S/JwmB21gYLWGt4ckaYBQoeJEN1GzGRTpK9De8tDF9/L/wWVLX1O8YwOb+lOywkvmYAwa7u3JhBY
w+P8g4P67CM2wQS8l6rqUpDy4MdQzHdNwvcDW74xtGRcAMoZMJs+1f/Anz+2skQLGUGGRtlSkV1K
82wCSaXxps+zkY9c9aOBPUFXRNtyLtRlEM5JZh7TWqjW/RMtVefrTLjCB16p/vaIMU7cvy2fTtmu
Hh3goXMqDbgzztbSV0aMGRAwIjDXTQlPXPcBigikVgSecZVb87tQhuEzI/sn+TOTElgiwngzFhU4
wF9HKaRnD/zeUQng3r2WvUdtYCalvroKSC1McTMdb1zdxydjrVF+97LngWPa29Ad1+XdfUu0CDQg
6dAtGXyg36xNIqBdn0qGh6Y4R28TzsYTxBQSA78Jq5cs7BEURV05zxVODqFnemMSjlV6yVQRHP0m
/Gzg3Fz3gcDKKxY5aEOZ9BIgLNYl6eAJ6YowRrAgbDZklm2+huz5nPnet+V8FoeiXNvX7YiXqIkH
hHQt1jJhg3QEYWru8+RQ5Q/03DHKxJCRKTQaqpVgI1UTieK+s8eWX6Vr418FCGV9ymjiGsGbz9lr
i0Q25jLSs/upaKe/hS8AEPI0DGJu/D4VjlpMPIzoa1XhnOET93FeuJWFkY2bR28rCD8FOERdY4CY
Rbj+r41DmyxQ3vdplUy4RE7rEKH83MCEf4TfgyVArVZplisuZXiADEj85s9TuQjyHyXkioFKQYV4
gl8R0/+vfXnLnW6++zuuBS4eFgPTLfGaNWc+9uoy84EOkACcFKqzG8DO6D3nHPy/maMuBV8qf2On
srMRF58UdLTq4V1CufmjfV6hnFFHl+Z+A+vx9XeHiyOBREvrJjtmNTIrm5DTu53ZlyZb2JPcTpdV
fNa/kue2pWwxM3xGJLYAlUt3Bdw/g4vLhjb/T5Uu50MROgVkUWVu2Ee+GwDGnHSRmABFej+81utY
6KW7XlSf1sjb8uuZBmsE+m5Fk/AWOQUuGe7Dg/eqCFzgTG9oh4OkWgzyTXZgz4vyKAsM7och1DmF
wZPpmf2esh8X1eOEP5Iouapb3DQV7TRUg4er0k3+TT3IY7z+Gjds2hGsy/DQE2z0DweddrM3NDzh
0hWQxYc6ZU9HcnIw9hwgIvD7jAbtKsMRttC7bfgOXS+NHIrg6alJZbAzV35AOIjJ6TvruHhGIYOH
v4Jxnv8m+W9dQPhBzIZM26pC/65sP+EjA795fx1Wma0JeT5z5oFnBF9lEDvYG+sNgjnzcatU4wG3
eZ5Zy0cqUINzI009FISODTfNYtllkleSmoafRlcTjiZErjSReLY9cP/n2NYsl8lrbKZlSPgNMywV
Z8AuWn/MFDE1auZmJTrfzlUI/8DynLjRZ/waYSekUEd9TTFpHgf9VTU3VTrlWHb7LVy2HUE+1XvH
O3AUcZPQtI1CUQfiezkRCIU0usrSif8vQXQTjEgw9x/q/ZdsASXrnf3xc1EvUOG2w/hTwagqhWFF
A7L7vv6oil/ythrAgb00Ru5FvLGg1QCtSG7ls3RA5VTSTaYvmpACO6tM74+j1no/fecUDRoOEDWr
O3QtzKzNJFV9Wz1ZYDa9KdsGtgCHk+WuBZdztFPmDpogdCZYbwsyFd1EiYY3/Shb8Xd0Ne1E6UG/
0qglt97DKvrmlp3ANLi42AtdRzBbGfIwwmiGJYIium/DK4eoEnId3uAkU9SjDHWGjAQsw03CTT0H
RMzil7vklDXve9Dh0TVNQ+X8MaasObZdGk5tgFw/g76FQpPHXT/lGgph1owAevFs0fptztjYdqbz
XipoxKACg6ogMmMtKNsDbp82i/esKChaxwmVeaRjyapdw8eOBvOmGaRQaP9PmfuNkMwRmKKJCV2n
3meFUbyqHqszUxPuDqyuZ6iR7HJbFx8Me95pDCOfWiy5uEWDm39Q/sbdnSlohx9sAhYj0WWxLX0F
09mUYRAyseLzN6LtF5NZcypV9jjHCTAEFBcXBsO7wa4g/B2Kw5Z1/7ut9RL+QZ5c5Q3ABH45XOoW
+DLeAhxPED/gdFQ0hl3gmm/qcpYvALEWJ9pLH1RRMBVSHYjODch8FqmWZglOeLXwiIt9xM5p2mVx
1rkpXkUcE4XAqsarMdmJg+4nwkqHTstx83J5zeYkUrG10NqC4+0+3xrH7IAcWvaTWAeeCpt2MQGF
ibMew9xNuRm3dQ4KcgPopu7uAeJiKBIpTjnQp8bDFla6OfNXUqnN+S3yQv5dbsu52AXKA6isRSiY
hC0eJJzAAXV8YzJaR9jd2gQh+cfMiV5zW4KZAHpOVHc2M3A0IrDLxeUOT2va4/pKEXgTO3l4gFJG
XonO+1GB/6+c1k/W2zGi2whZTU62B8/gg5o7JYR6UpCwcnICR881FqAEU+tGR4l67vqT/Lzp3r8k
zNWyevGLAOYoHijwSqAVHdCxssm6A7pP6DSHJJQXin0TvqIUCcd6EfU5pW68KURj8qodmEQzXNTB
TOTEIUfnhylgnIT8ArSq9+RrlZNvZLDPN+m/NwBTOX+L4b9TU77FKT4VGEkUL17NJQoU3DfextWd
BgozbG+EAF/BBjnpdqkJFTqwlX8KrZ4FRXl5IUgNx1fAjbfOwEU05vRwAWELplVtgdnGQbO77mm0
OI1IN05dIJMnriTaI1FRMXPGEFMuqjWdPCoXUSV6zbTqnwJZ1Ipj2wTbsgcvO+wSOAxOQb+x1efp
ng36AzPMvvYk4SQyNoMOlEiNTctQblkFWNU4kzDZG7/Kr4lnXeMYSCXZvnVsQrvlfCK00GExdXE8
ZV8cc/gOiyooC6yNcZtF6j88ned4l70Zpy90qCnlsqLPiXicIpqkd3zTwDcHzyb5bP2xStDGjlKW
0YmCHAjCEj1DmxCx1VJPeAVwHm6X6OA8GvqPDTCQdzSq/7oF68n5wjVn4i3+0eN5KuG7ZpmZ1zwT
gequYFiwBymH6s9Hmpq4PdleFessHlTOZ0onfoJ+hflLAZKlZwoZUOQvD5DsKXp14vvJbPABUJOS
aHFfyozEEAr6JemGIXtcl1SrxGklJANfI8orF0NC1avL6dsFJDVYiC3V9KkDxk/NelkTqsIwL/15
kzf4o292z3xjq4Pn6rQaYOHbROXwdYtcJvMrX1AFH0CiFmkt2zBz4ePl4WmN6EtbKrCjLxTB65uP
ckNjX5x1VUTw86tPsJxrRcDQt2Fr5RmOr0/DbXu8Ay7wLBbGbhUguc9bA6mG2pDyqDq0AhVOL7K5
6TflAmuaAbT/I5Y6QBhJmWNk11rRm7hk46HF8h4pw+nkl1CrAUhTfgfy59fQ1I2UyT1k5DCpbBZu
hWioaMi7ggkI/veFXppv/tDSSXcwjqm6dqIILwCy4Kj7llvXfOyz677KnhoCv5T/oKVFG2kJHGwK
KZ+I8cfHNaqLe0gHLC78eS0pZjewcGZ1ykjaRLcUa1slqwltvhPhqZNbREyzELcC+EZyw1B0ZhN2
1lFQfmWnjoBp4qJ5ZUmR0r3Y0V11bif1hsVWzDNWnoeyv0mT23vq8O9Wbzyv7RuHcaEUXjgFKgda
vU4keimJFDu0mUejjw5MEghFyDPzfplXc9aMFKCNpcRw7hHxjUDp4NcShuroYZYIS79Yxn2ZXJT8
uXl/h8o/PgdBGaanzhSQu/IsBJumjlTAFIeJ7z+AT28Kv0hoZ6FVFwm3iicLSp/F1UulE1/tPkxg
7NgKii1wfwYgW6yakpeLdIa67rPo8V4zKcnTs6DxsqxImm76kyRe73/DiRHSp3Jw4hUyIApEhRX/
nGzAPN3jhSO5YwGDlr019/V8Vj6OzHvRNCddWKNlXbKBn18HZstrsOV8uneQsCFHlqLg0YZHxboW
zUDy9b65KuoGGFb2klfQCjqm6kSmrSkqzHtryZCX1twKr7dsS8DbcKA960+5TrO7TWpNf3VWqPuS
UrC0Odl0Qc0GRBw9dIj+HE495FMB6ElJ9hK/AmjvCMR+8JzQxu64BmlsVFOL5Wh4CwVbMOoRGODV
rT6FUK5R4jyPenBgiWv0GBhvb83Eer3tOkfVsj+FMu+h96ZPFjc7958nFQIYMR0n1/cbNt8Fi4ur
T2c3+wEy64Va+CxoQR9C7k+ZeS1207vy5ULoxEFnZAH8EX9qkJXimNvbx5aCdVxzjkkp1iAVR5xV
3xqO0sWkr3jUi00ecUOKQffQmLMqf/WMtg6tX3jdAyy+P9t48rdGMnaz2/9yFHa4p6wAFSK+Xv7b
xyqknJtiqO+nxbJtXXCF2Wvj4JxngeMGtnH5eptzxArjzsamx0vD0XWEqUszMAVydeRVTo8Ordq7
3DU/mMgddEFtPT0G1JH/hJvqZ2+7O6lqHao814VFfheSy1NCpRj5bnBsKv0IyLQiQK0DPhoatl2+
3thU4eazpBduLcy2OO281J8J3Qt5kssc3LUEjPu/yZAWYnMmoEBUXCbLBGDwASLlzo7fW/lT610D
AF6GfsHLadmqqDIa7KMpwBxx16TtubThZYgXjI+WGb+lXN9dRlZQCjs14xVfm3iPDEG68OVaer5l
Km0Y0XWqoK+0IGVOt0T6IS9GGxKcKGR/vGfaiGaTvINnDxZOY0JPYzfpUj6oO1ndUy1z91NlkuR2
V0GZ0uMca2kuBTAPoU88/tRxnF8gOgqqImgo+oMHYM1237FKuEiissuMWoTlGRjAMxo5IFiNYqwF
Ak49FVzqouzP1SqnvDe9lljkVv8ds815RBEcDEeqLBL8g3sk4KFrXjY2eFpNODdxtqT3tdrafi4D
HI5DmC9v3AVaTq9cqQXgmMJ4VLlSbzit1WjejwT36Ok/ICPRjkQ7GjT3jFeohupWQOlDqK0AYTdX
lcF08luF3rGnv1QOZLLbaKJr86PswAISX/mvySvhRKumJzsvu/v1DABQX8S7LbpuAHJ1SEX9ZMLZ
AqnhqdYstN0nlmulnmY8dYq7CPYctbzilzaJoJgStL7yaAO5ox6aqmzbARoxe3S4lDySyBKrWq44
nmJ8c2fF9G2AnaA/uzHt3XoR7v1Gmdf+UWJ/SmyT+Tjo+QnBcR/iAQKTwkeDJQomRuP4qDiz4Lh6
S5pu5q1Q7DDVgsoJxjvrnjniVJ9ywaSu5T5GAPBEcEV3xpyeo9iYBiqjtr+N5YShIkwWCM0QoVzx
Y88R2H+lx9nJBsT7kOBT5AWnosVsxu4APZgWr3OiS49KdEsi+L8uI7ztBpvpyHDGgKrQBRnu4O+e
nOqUg3Qj/WiSOkbLwCFpd4d2dZl/MOLMms8HAUPjzcDF6pk/Hxb3XofvMoVwkhqKZL6xHz1bMYrj
/prusECXo0ikixou8Vbi7dID+2QvRjJVxmOBv8gtbNQPLSseKEScwBRCGOKniJdI9I6uhsdvXB01
tdIq28ZZF19kS9Kz7OTPcymi+I2h76I5qWIXMH/p3jTzG6v2Z6mGPqrivUhrfyha/mqIciOkPcfg
ZHtEsMRHfeliTB04RWJZZdz9CFegGulH9UkQPayWSG+V5KnU7PukbbleYbEXaRqjuIDW5MJKOjKF
uvZEW4C+q5NOskNgCQBZmKszdhPEP2NO9Jcgd7EdHLKrA/ChuCMF+2LFjRv5bEtLdiAZb0aPcbpY
7vBetSwd6Ex0tfdMpB+aSgJ8KW+JN8MfKNj58DOY48PYxEw5JdJW9JTJxDFJpTTYIxEwEsUv+6oc
ENNDFhJWyWh51fUq9bTCh8X25ftfbHoOb7syewF7qc0dtbGmKriHUGujmCKOtw7o7BKlNRVlG+1O
gdWLv5neN5/7hGdmuBrpYUYCJYjueeAWs0BngVitQfxg6f06EW6CH5r4SgHJNSSS0jvrLAQH8S9t
RMgqsELeHPwt1R7kxQ8MgJVZ/QiNYjCwMmgI7/C2bjklDDU/9bvcwr5DwU7Jwm0zrbTlXHkrTAnx
x7S1E0mgMS+Yedz/DU0+RPWvPb0Zm9BxfOnjRt2dmxCcfyhh5KWNEgoXbregsqW5iKFhQT/Xv3au
GS6MhnoDvLZIisYtsj0taYyQ+gUYihNeBgioKcEdQ4Y+xh8v/ZqAvCG7qLvaWBHTpLW5DstlWYWp
sfXLMLpf9+FMGRu15sNdpsDNjZ0mMcIrEHU8DP2ci+4/RrMt7+1VT4wpiU4b/KVs1Sk72PrUSHGc
0fRwGm4Jdv8614eVWkrn3wyX5mGnsdwrcpO4k87QUi9uaduTG4dc4sFIKW07A6gsgAWaooOdHwch
Wxpuk6TSznXowWzR1DMjBUEHm7EwDLxziMrbIrmPEBlPrAHvB00JF76BWxGnsDaLqe8JBXNfRuOm
sCkAm2jO2aPCQ0eS+FpM/xa1B/K62iUTNhi3lx4xPsEdz9Uifoz8Y2/vfKad7G1V+6U5AHz/SXfG
+oJOecaCHO3i5vwDVxqbTS705dA8QhobUVx4+GF2t9IngJDyDfpo8SKGqGs+C962WdAPb6gi0LWB
IWhxkaMdEiMR9O3PZHc8/C2mCha1558c2XJVDKW325rX/wMmlZbMgxPiBjO/zaaHBGU/kHgphdvo
5lya13K3P0w9C1lAyMYlAPH3xRSazceO4iqQusG33fyl4JN5w3dk0HjI6hk+ir3tzMR3idObmPc0
haU4pz6PZ1WftP1yfvBZsdVMU7ae4VqxWe0K2XvSf5mTdxLFCnJ6lMmMhs2vDndYcRegMiRBCAzK
OUQCZ5eX36HMq4IQLcuFEPOj8ss4rBWG8xKYgTVOJ0S6JwFfHUFglARI/mxZ4b8gqmsiZvnDZWBQ
nL96oERePZXNcC5yvNud/w2RRR6v2catE6aThL8Lmn7EJPr1/+XMjJKhfXtkFLp7cOzMHGHPGlrB
gUOV6AbVajTKG5vAb+Efh6GlDnAXcIp8bqslUKNDx2dG0xh+QkRSfSsqwjvfdBDfkVLErO0lxzyu
Wnons1gkiD1LT02P0xjlLjcZqPBpNnBk8djTd/VJDDOjej7WZ43lei/QEHPP1HCS7XbPU/m5Ce2n
f6WOexUVUh9BR+nnibY5DGDJOj9b1TqxnE5TRs5WbUsHVFIxMFPVQY7lUM9Qt5wvxkK93hqHLxtG
0AaZ1RyiHWIG3rcxRj9fncjYu4S1GfY2iP0ts+BwIQeIXQR6w5cHejEPZGNtn37kYI4CbABekJXo
OkLSs7e4INHQr44u1MeZpB5sbCjtCCQ9kjwUramE1vh4ZaweeMkJvLUWJ99sCxkTrC3rxi3lglH6
6o5sGw6hrDiicw+j4O3RAj9AKOg5jQNGH70ZJqJlqmsSH1ZBwJCfztoz1INu9NdXeGECm3StFElX
e6ajRuHEzRbXDVl9hPdazDaUhs048gDWqBJivPliDpRS6tV3nvPUv62RP462k/WzXbPXGT7scAzl
vzqqej+xA5WJ+j6Ucf1dMBNCzP8AI1kiSoHMFFmwQ+ob8Nn0IQ5mOTwJ3y3M3UwvolAdsvyWd1yV
0qzJnX/TyP8Sjcf/lyue2xZu1YXwUYgLRyvm+8N46sH9QZ0MTugL1LEymLgCVOtzkiVKlLipnJj5
0tiSfWHoRZ6awASYHA0vTdR+9/VVFtLD+BpW2M8l3MWKJHg4N2GZ0sdp26BZBejO0UpRrxvjlpuC
zS7Ceru9ujMzYWL5zPxoh9X5ufJtyqm/uAqdVly7wONba58PV0sGtLFjF54+qlY28PSqunA9wuEz
RRdN/dU/yEmFtTKVMJXk/vcjSkFFN3yOWX/grFjz7Kf4reic+apzbZvaYarjFQgf6IUxowYbnbuC
p3yljWeInxx5jZEz5u/gQGThEbBNynBGh72kXuxLJHHA8J6YCK7DJbJ8goq3uf7a3ELLbsZJEWyA
lGaRktENkLmaPFZLTI1jV/3Bxj+Wlqvv9aRXUkTTm/kbsjmMxEf2B1EJvd4u32xcHjDHZUuHNnZJ
uJeIRH0+uP9VeIycrWREecFMnzwLjAQcbM/d7M9EK6QlEwnajQNwLg6oeqUp5Z+Z09MgbqAqdWQF
wMrSL5I7dwAk6zOSXaFPKJ6mlEVYp6Nrsi+62rzSvQI0Lj768NLpznaxYCrqL5t8Ro7w6T2hSXNU
MOesT1hQEp+LL3ifW416eyCp58QfIKojA5y3qetXCLs+Nx/FgbVyeVM7LVSEf4YfK+2ARnCFPhmo
zEN5P5a9lN26a/oWNEaS4LHHAga6diclm8qlRXENATQ0MgYnK/5K71xSt4XKb3N6jFDhGLbyRdGd
1eyCiN02UE+bYV15VNtsfjyDbEJ8+L6AKcvMCKzKhlWP+Le22uF9ueiM9G85/KZQ3eT3uOb0bC3B
rCkWSMLIHE4iTNfFZ/mcXoV9Irv4hD4fLHhLF3EjECmx/u6mUA7xIF0oRd7aNNl+JwVsTcorLvcR
rkHztCa0qqz2IWFNYbGr6f9k2tzVT8oX+aPtw0hMU7/K/A7Ut9EbqesQ8ALy9AxxFfyGefM/rr2M
9NCb/ArI0VTNgUbkpdL4LBdvQDPyr0czZWNQ9p7jkhqe3EyovmErxMdgF6TbAWD45pIXaKN6QdXe
/rl4wwZSrbHwvxZzI/JpbrA1PkIJJfqhWOVAvH9/PKZwJUvIlCbdfAiysJof5Jw8kzTFBfPNWiUy
0q5MncCZyzPRNB1FWMRSiMhv0ANKuaT6POUEcPu8ytDhmUIkZabDrC+JhCo8wJXDC/WG9VaOQ2xn
p6aD3BASEvt0Q9ePkJh7QUtIE0SVki9tuyfOcudLsEfgDkMi5zjMHXX/LM3IiaLr7CXn7kyJdEZg
ugGjSMdf9/zGtZCD6xQ+EUNnTYTa+xpFnW9WPsCCYZ4+20loNDxb1y6q5DDZVKWs5rOypfg3Z34u
+2ii3bgRd4/7P4ifgUXmV21i5FoiNQ0BQx+kMoUi1AKxGNLpjtLg4kohRMKO0HwLgLo8DuAi86JN
7mp1T/Rgba6ei7yZc9v9ZW9VobYFofR7AlgiXJuIKyvPRhzp2r2pO8cZS1V64BTbUOBW3VL//hEE
Ybrt9x5A9e/wrlDEDhnl+795i3XZSWnfVQtfqBrriOmwjGwPX/VBehWcW7uaa2X/sBAZcCFQIwvj
VZSmKJgGHoDD1IyAsOkHwPKXSPUocyCDRy5UwIBy2lG/Di8Ix9ztmeEQzY9eDHdAZhwsjTcOXud+
MxAILe14DWaO9hQWDvGEX2ObCNmLasLHmCryNIsqk9ijT4O78bRrdY16KhsZsKlFl9SlIp+1ZG/e
et19G8JEOac8CXxLxgoTC7ksaCDQeCf5VwQvRzbjXfp7BJkXgB1QEw8EoUYFcx1d9h2xHm8yoFd+
/03PA2fVsQxb/J+hexUoCFmimteHDwjs6ZIO+mAi4ugfclJhWnTMFOd4XIKtnxz1qGOrE5tUfZd3
uJHDQ/EY9ZMeAk/toVTGgjOCko3UAx7J+pA//PMg/bp7B49mGroUg/lPtOu5bIxi8N9RwjqxxG1s
iOSKBT5208gQxW/RCkyPXmbXCIIUGhIEcZBw42CfmR+xIaptRQxvqnx8QVQ9RPke2N7X1gPVBRsM
ub943+axUUfQ/YkwI/UrNmWljLYJQsynzJwB3dxTArRJ0RWF2APzKrxPMslCNmyHlT85LG5LvwhQ
vwVTL8hY1zQvY8El67TpAPfIgtqCstd9ifgQqkopUIDwLsAXaUkNmtdmCqDCmPPABOtHwCyMf1vx
CkpxSS6sXtlKf8V61G6LWzukv2+XroIMtY6zhfXA39Emp/L0cu85eT+0VlIuT5n6+1IP9tg5LdLI
FS+pw8i26kQ80mWxbd04oRAgXwgKzWFYFptjKR2DzKt1syJtB+uO5mhDZ+p/WK2HhvG7q8ErIDa/
Xl05jDsInb4iHE0alsQQKZ7ty6DESCFyTRlGMJPte4XI/CxdklfdWLjZs+OUXxOVq1NFgmLK+7GJ
JYMwqyPv/a0Se02T/BbTwSODE0rmyXdUWgFGfbSdvJ75X9vePRx49lbT7JXQSm0JgNYpaRKZoDeL
T1husFSt6dEWTN2LBVTCSLpPwc0JA/Ilm7p3OTIVhT+rHw8PGMcbDt1nUUSeraKMGJHTVZSBD+wR
Q/Ht+eyuOMwR3iZ0bAWZGHDO50eLWwmcoHmS5MsHbllgrGGNWTPv7Khsh4lVbFcE/jZ25zsRKvPv
QCDt+POLL/SW+epfGkY0l3Q+phMNceTfwWpvLgNIghf6l1QUlTA7J8VNkLyLn112dCiqYTDe4Kh/
5mRGpWXBgYu7YynPBFkXQkQv8HrjuCPIA5a8qLR74DD0eOQASAqFUI+ggawba4pExcJGaqFxpGE/
SY9RJkQuTxBxO5J+sY/YnTM15sn+yIX2acLUDQ7jf7pIM1t2gqAOqUyvaQ9Sn3VWxHH1ylsNhH8G
moVCFMK+YxL7IqcaNzS+t9l+Xhpv3iBjMsttaH288fcVcgh++pWcpIuULe1Lg6wu7ZZs4U9W2qJT
mxbM+x7bcvrGcmam3HGdXDaqVNvbAwDZwJRkw7ipyl9bNd4YSIUArib6Gs6LkuRSitr54L7++a54
eMR1bHsU+8BWiv/L7Cp1fkqy2AsQ9J8SMklq/xzzrvJ3si4BvT83u6FO3EujRWOE+xdmAnXjBLTW
C6QcLZ8mYbBuSAGNVbkZR4klL2cJvv2eVefbRqmZ1XiYgnZB/m9EIZ5O430qpBdowjoKrtIO7Jz/
jUIPyIBt+lt+qPcwLp4z8ELSt1OurFWjZuUr4bolQcxYwDUpRUZ+P858pIDLdTXGVpsJR78gLXfx
yJ6QuLRZ4LndYwIPnckD56l69aE7XB9Rz8atyHmUoAANAEU4gMc0+sgSz0+dUKQmNHo6vVQ45tMN
0cuZ427aATna5d4m+zUu60cwEPEbMYIRrO5546bL+t4RGuFZqkIlEGXCNOqz+m8/1VCXHZ5em5iH
CdiMihAlRnpVhvSpdalFca895USlujDa9zzoBN28uxXiMGuhmoeL8gR8vgDdFVUWN8e7S8HCJejH
AVosieWNUKVZzkGRuw2r3Zc/SlK3Gd2tE9YSUw0tS0DM4bjBWqkWFhVQMeAiSnpC/RyfepOb1oYt
p750CboCis/EQeej8qkCtVzw5/nfQ9s0YZ6GaVEE+z/b+IiM/1iFT2xdIz9lkIEdvv8nVDgglUF8
DFjuULCWqyFpaV8aebv2xIin10UyiTgfujvjNHqmYcIGMFQt2MBKMqm4U60Oqn3YlgmouOUFXTeS
GG4G5F2jQxh8EjCj2DuRjH5goJqe/dgdasMcAph2saXWfAlZWqYAY+SdJDCYastUplqlu3haI4iJ
FX8AbZsGSTmvptlfW1AXBjIH/ycMlvCEXexFAhDimsSYVIcO9rkWymyuNi7QfU8o1kTwlVzdoCPW
n4VLUkwO+3DZ2G/Q3u6M8tAFDP+jM06VFh9Lt8SOgUNNdQXgmKvrfvYOOj1tt20bWekeVgwgm6tm
ow/RFHuIx3Mr3lakFU7Ld0W0p50J//Vv4ZJb4HBjUasrLCP5l3jSV8XsVefpNPb42D1fuKSOPZnB
WsBFMhL3uk+2T4JsDvjiY8mubaSiHPAqSq/vgzaFgyHiVtXkNK4+eAr8TQbiJkqd0DjLcfsaxnun
KW/Tzc12bWmWyMD+vFT7Akfqda11YtyOqWiFY+SzngBHSGdCdqVrG2IDDTU11xVH5vdfwBmI1va3
crk2Rr6t70S04evercbfF2zCGFsIbACbMdQfOIUS2BwI8uPykF2Tfu4wwwhAhr51uXN9Ke50+TOS
NY7EC/0UsKum3t61DCLUGVlIWaXVVgkV/L3M5NNGkkWdw0nUVSZQnd78GosJ8OkLpoc8lpnKGOS9
vAyVrRz0LMtapWdqmUMGFHY3sAW0xr0632d0S/NNrUhCRBLJ2Fhz/TDaOHlkijrx1em+56ifWr2l
dKKSybW83zR0uq0fzyxb+6sDIsvfBKruW/pI3OGeC3bHheBaalE4b9cZBgDNhiXOC6cWF0wEXJIG
RuhmYL0g8hfY+HPn8OaiAzbDFkb4DAd69ka7zKce+9Pck0K1wmSG0LgLzI6d/s03I4dKUoNthyGm
InNjSSQNDEj43Dc8Kpe+ze3FbpezRlmIumKA5qhZsA05GcAi8O6ylQDS/y5vJkF7USZZmD2Tl0+/
CIH9YbDrQivr6ZEGBSl0OXTge/7OU4VhEg1mmxgfsLSmkbWAz5QktDIHEhm/svjFTqeoNHk49dbf
I5FXbLwaeHa8T9glmfnMuuafCfiprgKGW32rKyQEywnn+9uZ2MQFOFkAimYql6x+6/0CdN0HEr8a
datPgcub3yU95KMyinHUg0z1xoR3wREjI3sUW3uGrU534JoPzEgcfkA8izqis1i7S5ppJT/y6/Y6
HB5vwfwJtXKJqeW43EYCcF8IXgniOegiCuleEOh2FLWy20thhPp95xBZ0Qh/mpDLtKkL06n76dF6
R9KMnejpIOzb8j/X3duCU3WKx+EMo0bzLOlUOoWr6PuXeAtuuIAVAsyc0vnK3XGsmyT45r8v+Hof
AEs6zx73qC8LR6UwjqaGDHlVVgZ+bVplP2uo82LhSVaCrDCbU4AzRBlE/4cE012YtLCtU5VbHKPR
5jpU8puki8LCtJKZd4tsGlTnzDS9eqkx975AHTvObEvQkXcqd7EUM+XcNc9TUyTvxOBjg38MtLFf
xIHYKJIeNoXveHTrZFCrM4kJZ7qqRBSNgYjgrXz7+41NjRZ/g/z0OSSdHwR3MBnWAUBFGMF4d4m3
1sWmpWcWAJxN7ehjw4WLaRh/5VMaT4ivdNpf5TTCsS4wTVrSPexugv2irytZD2wNP9Y4cXHmuiVp
901+32rwcJJY3ebPhriDSANNsgNbmh4VtR1ISfKu4C6tM1IBx+Davy15HFksNgLgNLlrrVrTXLPT
Bb+RY1zCAN005MFX6Hc8ZtgN3w/+vWpW0lO1GCkS4hmZP35KdLs73twbyALg4eP36YKbi2by4YhN
NNTevMJ3ROqpOT1uUKldBToW0tcYbYF0CU0HgE11RrFnfY/VDgpXvQkpKahPn97WQxr3mAHCeVG3
+i3tuyUkdNyYNVDSkXZSrjcTIINz7+x2ovU1UySvmfrmihIbtX06G+bJUqW2v/7WR8fi2xpNx/Gu
PHqZZW52VGxo1oq8ALuiQtbKTnS+u0Ve4O3Cj15+Rk7kR2P+XDO7uGfH6fr0Zdh35GKxRLble6KO
ujz3eGFsz0xRgMacAXn79azjsrQe9aEJjNll2hMQJNHudNsTCcV7SQe/lMFrLaznSXA9hmpRPy2X
NvuodtaJnFV2hICNLi1/ZiUMePe/EHFnHqI7cXeYkG8LLJkkjs0cH1hkqIQlKrmXO4fwXG2+UA4V
SQsV1MrjRGBBEq43icaOWahANszIRvZl5rVLJaYSGsWgazduhBfT3relTIKkQRgE/3HPFFqn5Fnb
9Jculyew7xcJiRawpxgPtHZ/ofCJ/L32lF7qHeWZtDqFqkjTe2qmvkCq8XOdcPPGeCtT4f+5j/VM
ZyPJ4BwjBn7NmiYii5GOWoSYdatDLVtLQzbT0+I4TquDlUEJ3dU3X+pAElB9LwBGfpsZX3+CAXW/
povhuyEuVzLTu1X+apGIoiiPVYs0YoR9Yfdt0dGQEmbCsn7nvGang/8SKqwU8KXrgDoXRIkTcL6L
uQht8SNrFVVdYFHAG1iWi16l+4g8fF6p40SrDEO3jVL02TcrKsGoRlAVJ7Ejgd3eFV+7kXh1OXqk
yI52Xrwu3mwUvFEULMEQ7sv4XJqamK2NGnCkPsmdnt7nvMtctv/Uibj57l+ZPYyHQlTmMuzS6a92
T8iOD7yaRlfAU7ANfbRYGbkNktdQzfQ5J7SgA0aiIqZrmxMjpMMrQrBnOncn0rElYZ6TRTrFnOkI
GSalVN0b6QU1HPeyEL3FSPe4fUtg7auVzMEFBjaznEjVSWwMStMxa0KqkUikf639j0U3Sy8VbS51
wBD5JsrBqx06Sbgp0IBOYdlf+1L7SNs2cP2RQars6ZD4YRe7RYNADMT+AJyRnnVM2yj7KTbrqdPw
hH2AgMhLjuSnK68Gg1QdIVES3hUt1Hmrtz9fpXBe1FqHTiIhKTTtsZ3CRJDRMdcVUxInH1V9rG+T
oOI4YAJAtV9qiBO3IP+1pFkR6nf+n+m/Qu/l23O/t+mMUQv554IOK0Ypi6y3/zOaqyttPLkeKzz8
AV65XKPeu3fvaoK5P+l6SqWJzBWQBrD2rpT7WRsB1302tdaENOll0JzodgFcpKRjn2YdTYELpE9H
gTMvHKPATHwM7NU5oVOdgaf8p4J2X37K17dgvqgXBI3P8NqH4NLbgJDetp9OkuHmReDLFU6LitK4
aQsEO2zOU2JonHx3ijSQqCbeL0VmDqjdVyWg9Wm+FT/aWXgGQVpC6bo+6gMpPKrP4hPW2BfzNHFX
QfJe+WsW4FAChkryWzTnrVfMZbyfZi3fl9bIw8vbTi+hjHIJ9diAT1wdd6diQkBzPBJuakZWwZKS
BGbS9mmh7jhcXNWuGppzTeoJjGwoJLDX2mZT8Zbn0KATuMeJAvmJCUuUrCG06FqAsqCGIbEVi8fM
63SABYaYYaVrSLA0+vz9mjX8aW8LJJmCVj0IDbJbu8Exb0nsS5h+WmcSKBuKVZ7PSICglbCXOWIX
PMs8mrXc+cPPFsXh9bdp/Sj2o9PhdBvsw7Fp+GxFE5x45+/8atTNpeg/1nNGQIgnu7ah1jtJkvTV
DOlFiv1KqbdyUUSQwpGqrtqkvjvmEzO6Y+YttVDl6YZZLRTUtjv5o/FexJJQtza0lGVJciJNBUIc
IOgEyzD57KfPQ+hXgRQpNbeNev7uMguQRb4kHZI+uSAo8M5CZ/XimBGLpqUxpAUV1IT1iNF2r0+q
48kKUDpIE99qmPDQhKobZ2NNxRR5KBnb89ZxfsWIgxkGmrzUDRT5tZ/uUUjR4hiFJHWP1t7pmf52
ZRdCMngMwfYHd8lGqm9JlWVitxW08kZTmPmA8fiLoJNDaYn5HylGxdywYc0W2VQJ0sFOMVHG4O/H
V4ZOXJGYNzsEKgH6B/vn3TlDgSEhTI05zV0UB4lACkT9w10qRnodjaiyLSvLplD5KGQ8Qtvi4alR
E7rsZ/XXe853xOyMLlrypJca5SzETC+QIlMngnQu50V8Qi1XhtnyN76t5li49nOF7iujyY1DS1IJ
zhpkNJ5T7luwtb1DaupdW2CM1wvulNNUAFEsN93NxhRjm6M9ZfQidgszdlYyDASPwWfNn685Eopa
Adbh1hu0Rq1bubnosPcSg4DVakDxjmGbv3NvHI2tY6ntK6kl5w8oLQVRGStzvG0iFltnBtUMP0nO
Tg9wLAvzfivheo7OGRs9rqtPnP9hIcxyETVzXKH0tS8icT14u0nzI2rvsRLV8W4JcYfyMUT3JJO8
uSnD6cuIJqVVBNb8l5NPg02ENka2yhvmheqkZPQ1Oy88KovvMBkrMQSeQAUkwcai6vjiEx0uYThx
LJRxwnVPHARKkOe6WV/sX10wBxQNg6IpoM9MBi+iF7G8otGjOFC0hS0Ov+FiB2VlObE+YCx99FH1
LX1h+HszgZvz6F2QfOD3BBBYKVGwQRmA9+AuCapN8gG3L71Wno5xSVahSLHKzCEIhOGD+ZOTafdu
DHfm1DXTXxYDOw2BbjzTsU9IYAARRRtQeBPJLbl4+JKM3EMEOVXmvXKTPfEp/smmsaw0ufHjBovS
X5GCPOOzLuuoMI9n3z37uS4uRYLAqE/42A3k4J1MlOtOuACqYE2FLb9EJ3Aj+7N1rQtTWia+dglZ
heMIZOvEJ4YODZuDswTBHt3PE+2ly02nisGcj9U9SDNDaO6wmLNfiyX5+L+NRPl4pfhJt5kySmrb
rqCPVxnSqYS2So41pZ4dmcoghbmmdj7/P5vnhLbevEuKlkFrbq894VINteu/IB/H2HmpCz/vvOOf
XEIP9UFmEiEr7ZW4y9FsCn2Jly9iAibV0OOdhDUHdTMFnKVw5r8ZsxMYwkJ4cwBvLxcUW1okyIk2
QFmDiKGtbGzUrAmlJf5D3LGuv3rOOC9hhFRi+2yqYLfOBy2xmB+pPpZzoK7XIzxcSjXhrx29+Okg
GL8mR4dxUjLfkTzPP+8NLtCEz6qdasFYwKc1OlZok/FNgVcm67X8FG3Rjywb051cURu3/Y7ZEmLN
wEhIdvC93pZEYO3bARIHpwYUURf+h4yEegXRdtulH/XBirRFRilLli7MvoBPtx698YszskCxaWlI
1YfQ9jdoyXoPEyR+6sOrWNo3lcXS3dB7sQWa74pSjCCJstkMbgjeoBW8zZFV1wC76eAToZvjSYkI
1piZa4UWZVgmfvX71SKFh+InSySoP22Vwcgn2Okd1Fq4RhL7AB9d+yOOx4+zQyM6tHi92pIdhe4Z
kxpNiDzoKc8P4EE4nY+8Qj/wfXfSPDS2bx+9tkSbR5nCmUpgVUu0agI9jq1GCrmulF+MPjY1zljU
THZ2X2L33wXRKhWAxT1p8Bmsqx4NdcBGM3n3tTtHnvLe2wY7InF3ZWB+8umYGB7rDNquZ0Q+RPPc
+jgkagtz11CFrEmHYqd7xMHPtqAs6fgtBeLjqiBOwRnMrfL1xJkizEPxA78H+iUqd5mI9nYUzNUL
jk8YdYyLUOirFI6841VHrFJVophe0nCr0d1Y+M0vMLSjNAkYcnPpC/UFfjUNgR/stodxhGPYP3yC
7iotGx9l3y9MGT0iaYmIXRsUfm7r+Ct0A2nkmxcn7Ig+PI5D187tmE0Sq7jv4QAx6+rdcpOy08NX
OXTx54DeCu1J1TnDH3esNVv4RmPub2nRgxZOP7IUzqX9Cz9PTd4YNQRQS9+/3EJrS0pcMlsHnlgE
63BCDP3tb92iD/kNEp4xARxmhy3cGOhg2HZ1ZQVJyz9tnJQhUE4FHYky449m3UdFwA7gnIVmMBKl
FBoREV3g2AG2hxd0xwyDlVqHzEHU5deM0Hz/X6vVqLhEH7aZ0yL91ebhwciBgS+XanqAfJCqfL80
+ekgV6bqNyoi/1wadtPa/v+t0QUXoxwXyCmiEn0oH9YPpjG2fVzeeuLvto6YCL3EdWAFddNEbExe
d30wjbzjecu3qiNC3ByvO60WZ/SHBZ14b1vq1ZvEtiBzKsEPxbUg4ZYsVKhOLV6gDrjhXV50Y0UZ
MxDhPkLOr+hafOtfHFqiEnt6tQKUSQo/Hpz2zWhqCa1UllEYRXGKOlyM3ZtxbpcPyYbOourdlR2n
4GP1JpjrRcp6iXIrfE67ZcPGRuEB6/VFPEo/wpaFAkcNEsNEChEpicrlV/X7hT303BjZgwxxjrj/
1lXOSzAT7I3od3rni/TMwnyZGhB5jAmwM613oT+Ulx76tvd9Ft518p/p3OX4ktTielvGjbieA9Ja
yyje0rtaBukRgQJFx3+p9tYLLZUG0Nmk6uMdMYYyUeDEFYFcYw+DWonRi+PB8i8MSlh0GPLkKWHm
AiiP2ihPxvx9ft6oCZ+OY35KHTQOMUj6xR93BcNaKz12N0PDcjy9hDRqIz0H41xV0agmIHYCXDTi
STiO+jbaxbdL3k7LtlvxiLoIjhBRl/7auEOVzqAYsElP/YgBayT1FbqZ9AqrlkgsfIp28pbETaFQ
UMIPwAYVaAhKNqLs7ErUNsoJIphm5TZXFS1RVF0Z3vihyBYOwK9s2oJBE6Td318Bev7c99N8hjWE
4eqXrVlbVUx4h1owLm7dKaNS77gt2Y6idGnI45sa3PzQpgxgFoEAWooAkJHBLPLj744wo3KQyx0n
eHzNlgUh9smPfIZYx/qCTRcxiWcZwNYK9+6BvrPXgmSmokLr3dR4Tun7l5a20gduEWQ+tr0EdP31
KHxCducD/gDARR2E3H6fjh4DljiNpH0tXT5bmmfg/3n8Fvb2ydiWzLjhy5Bs01UZx2I1zfN2Y9Yv
Y48kp51K52y5qd0PaiojmK/hgJa3tETdoNoTRwM9j+bcKp3rFw1oVePGq9L5hFHf7XQ/DIrwDoW9
ZEm/7fJvQEtYshWwDjPZp0lYwRKuzUdQ/elxd0g4n5apdQCQq78m7bmY1H0BE4RmNZqdlRmL/wbm
XCAmjPMU3kHUDQEAS+PbJRp3f0H8WN1zdNkpgYH8cGKYp2E3Fmo4qdTJHD0P5OjrUleJdwvSLr+2
KGBiUAWg2sOwMnFTp6pkedTP8QXtoXuAjSN0+TLs4gp8RdNeh5PFzlaP4K8fXtNpS+CjJWe607Z4
1tFr7LT3ag6XNnrd1leWirvOAxg1s1SlHOwFwODJrtZvAwl3RldwjxZOp0tz3iyRllg+0GP7g+gX
gfFYmwDzq6WKfvWpsPWK5Y7z5Mj6sgMDcj6OQp5KfYaXCCXKQoaxRsG45PzGHrJVfGZYs5B80Lyy
8qHRouGFrnUvgMFlh0A0b1F4yaL34QISRV8Wl4TjHtfHRYXV5pW6da283AtUPgqFcIuFttf8WaN0
BlIegRPhqiU1ibv4AbnuKPO28sTrXb/5jA5yiL0C000mfa1XNSuEvzvjYYIejkI4OuX9IwG8kUlW
S/N/PqztUBzjBHPsj2e9Iojlc3yKkw9svofXEAxTaVLtWR6yzqPg6T4KXsBjFAjkAvxriEWs/dIA
kvJ/O3SdcVGY1YDFljfrLca4/rkMfr25r3KXpf9MhJsce5Bq8YRV7C1nAgpNNwMzj+jU0kzJV0EJ
Mn8Z7S52k0wHQulCyvI63K56NcC9mb7flKM6mM+bTkyThPW33mHNrYOz8mG/ovrhKCipM9YcFzHG
f6Kj2av3fqLo8VG6mAOgFSj7Td/wAWAnHzzx1qYbBuRO7+DDHe+qfO96BFApXGsGjMQgzAVOt5su
UcDJ4fgyGSd8ml0w7qj6Iu2Au3btAHwTGoh+KhQLDnydoaZrKlh8DeJxuHI8Rt5BvMEDF/13SRAD
u2I95HgvdXquX5PbMfUqU0AMHvlxKdl+JGoIV5rEDs6PjtKo9x0cJL2syTJzJ4UWpXC9QRF/Katk
Votz0PN37ekVelAJDfA+epuHFTrs0Uc/8CXNy7Sx26yzTlA0ZQPX9+w6kzQmuUZW8UJEtBJL2JCP
0bQUOssgyuYXsexHHfFc1qTdIV5MSGkFp4C/2Xzu9uyOXiKroltgdKbUuq5gbIFUFVWtdhrzB9sd
8/h+z442buEtLehCt/hRc5gCFmUDm7rq31SxuGhMYHTcTZQJqvh+2hY9/91ZaVgAhRMCtMcvxR5z
YBNUFrd1xRO39Q+8s9g3Jn3FaiqBqYNuhq7B8UGdLSFkB+jy0eLUBWePS8E4FbMnGZS3NPACat6G
fyUTHD4S736yXlmYV9/yQbdVZPvjyZVn3fjmrZQIdIJaoRf0fi9RHEndh5kgGEhSea57rQB4NNbN
fpc+7QDzWz5gKbNlnhuRJyvj4hQsaa7+LkkTpybSlwzyf3qGslUrjjoeyMegAnGif+ADlAR4dXgK
05MESAjlyqsXANmv7qk4E8eqtcc4lK74aAMwXH1Ti70DjS6EIPEUeoDNkeQRFzWtZj8sqI6myji+
mwWzVtDuXyLwrcnNYSgDtbIwkOClGAs/swiDe4UNqHO+HpIqhCJCXwIF/Ynpvjm65HZVMISPZXW9
cwuDPei+wPHRjnylVjSFydzBbT98qgi3ufmc6cq9oSeQfZeKPHCFc0rJApW44eSnodx7nJMsWmTy
fvQLxOyUn8lfLanfd0v9qnDreKFZH7qyUlPPzuNbgPcFXW2Ku21M27VjqgNHAtyxJLaAHhPo0FlL
/T6V3G1ouWJ+7IUvO/J8cRp5fLvFBWSjOO0OL3UuTftOtEEz7CXiLnbEZYt6GbzK2sg3hZA+ePiA
ABSveAMp+Zzcm032NKhSdmidq2gChvY3gJm7fPbyY6P6ckC9NnwDNT03RtgIsQtI4fP8jCVKsuCu
fib9K3k9Tc659Jf1utI/rJnh8N6jjru1oFz4z0KUOr7GaFZArf1u0LTHiCfHr8qHUkHB9jvfHzMC
bJNWVOxOzOCZLRDmO6nfzDCt4BB+lKoZ5rJow5sbvqg78MXNPASmMWrMQTNkVkY0DvXAGbkMYDGO
oaNAfh9v7Bac7Det9/mJBtz9VZ92DwDaNa7BbZUOvSJuhSlqCxvH9TgRCx+SShQT3/HYcDmhs07x
GS8hHH7PCx0CjzO//5/r1HSbqq1J2q7VlT0AhokZ4fUEfQfq86Vuq1dHJxxguXdQQ8EtYsUaQF2G
gGWVGvab0szJFpe1g/PDXAOGFz1e0/bMMKi42tHSmCHsRbG40/EsfRGorFr7grUc5Az92Aa7E1+b
XFesOkFH/LB4zC2h1E16rhjfLQMqUXRGA6z81Dik9bgF2rwRlTUslTO2YDXzAfr0NFkIqleOyOJY
PuX4iPN1rYwGr/21/zWasUxLZn8nX8Xl7L3gjn+YTOCRS4FhaJIGtiW+sBqOR9lWWSmw4i7bezNw
M0HErHnV8B4OgtDleMjAsa4UohSNWtbJjKMJNNGZsJ2rFx34IytPhl8igwqLNHrGN2lhMGNtiw1n
Xsl9YAZCN7taFPkVxcRwd7lagT+g5UO0w5fWnaska1wK3MRLYvd1QQZXxjPnRFdqkgQwYePjbTIz
0ppGB5xMoWKSJpQlDuWKJZFTpCrX4MKhQuPhmmihnQdzG87fYJIbdPvmAOk781MIYOGVi0zoXAPK
W68cVwuZ8maRwdpw2C24IpibJO20pbzEUI5TKIxTd0Y29h7Dt80bbsU/s6s20mJTp0u8/ubfT5kO
PJMzlojy0RpiShN9XDYM/Hns1YLVqcc47gW9qquIO8AZdkneXHhpXdscFNaKzvBrsnPZ7cWnCjF7
fv0FV213ZfS9y0U8JCz3wBlJwRJ7gHBBV63J5m85sMfNq7UjV5yaKWLGVoocpRlsS9Cqlpn5iv1v
H6cMiAWHpILqI/6ghgR+dXxvCwwSHZJotXIZKw5ME+3SWzgFnI12i2jIs9vTlW36JhwoHHt0HMcb
3BByg77U91U3Mt7sm84GUJOiYauTnstn6mD0os4CPyv/jI6iOjT3WnM+jo+cYXlv0TMQrys7cgxf
HhBF9mzzkmZUzwAB2BDqXapy5+nyaZrH5r4ATzJY53Rmr/NIjzHHZd47scUYiyfOUJfxaPVQoXSF
2yVX/fyjJBKY4reFZyl95MgCGryiD60tZp1Fl5npi4stSxf3MQhb/XJAL4gaHmYct7vyw/eHPBCi
PK8Fhb0jwEFNtXke4ymTYUBsev8PcnuajmGPbzZBd3/A4+j3GDjY0H616TcuArbe62jWkv7FQ7AX
GJ3CCm6pTauByhUMKvc+Kr/mpukTTYQ43vWTXeFmM4suTVZ5TvlnIPDTAmoF9/SD4rKRgUHkt2/W
3Al7GLlxPRrVXXrdxySqjxLxKoZRZnFviz5zjr1oIPjoIvcR7mpY+Fu3n/ZLPK/5f6W6vDNUGzq9
NmwphYxGv0rhmy3aLJq12FICC18XrxE28B3JGyqq6B3bk/OZ3vcTpCbrop6fW2w+PVrCLUW0jWRu
4TTzYbCmnpfBR4yzt3P+Qq2exRV0Zr7ZZqjNafohgUdgHXYvAoVYqPCbybZroKohwFKJTdca6llI
eeQojsls3bLC36/3n2SI1CU9VHQZmt6uLnZypTt/pcf7OoWnKC34cKV5I+VJITYCcKJGY++K8WiT
5AEmxz0Ds/2lyfuZxuRfVhcQMq94iMWabGEeFkYRnIQrqlEY1b1DpHSGTgzcTCwNPYDPYU5zjCZB
7cH4Gu6bc/fkfGv7iRIL6EubPBLxB+MskG0EexATICx6i9FKieqq6pD+5hTMtLhpDphAR0fO0cbC
UdPKiynd8wEBdsrGqmQV0TwC0krygXnghBd/syWxA56kbnNjTD4RnjTtjzGqcwz/umHdyZ6CikvJ
/FM2h5b9/o/z5kQ5gia9Xm63EpvF3/CzNsz/8p37vvZwGX84NuAJrfNwzz4pS+HYPJCZYAdW9XRU
nmefZdlq1d34O6d4UCoMOzvB65viLXpMBytytD5DxM8ciXZmGH9vonD7S3A9d31+f+dM8D77ml9I
Y347trOET2LSqYFdeE4+BujWrUNz8Gy84Fe5Su/uSqkfzyOx23d0JKlwld4Zu6f+s+f1qfbjAnp+
Xoe5UjImfoKMB7smizKx/bXgRpOA88BzUNEsidebzqUBObscArLoHS6veCdyBXKNOjmdMDFQViSD
Avkb0lhfmPETFJeLVVJsZDRgh4P0PwNscJi6V4auCUeEWQ0AKHEOphvtZxI0t9udVnF1e+iWg+oP
N+AJBydBBAXG5XmOIsw8yhaDR/Odci6RQ8ACOfqGCsgk8SiZe1QDFmot+8lr4c4DoXFtm3ePRdfG
eTnIlS58L04PvC174FRrjHpLHqeOFsuC8cwooElsI2BK+ScZ8vKMMpVLJh1tsbHGEBkAMvZb9fwQ
Aw66hVYXccVqgZ1gJe60aYIz1n8jsGWuGDCBg28k0yWtf1FA0e4c9VFFNW8CRHDSVYnAnZ8m++C4
W2+WvfMc+mGgpjlcY80rAvSBF0z4jEf1yAjs4jO5aQIzUmyY/Xc3qioOtmERMUEsMxN60wLD2Iku
MP8mPCAlBeWpSWLCBkUP+7Q3opN3OUr6PSuayX5Ux/PdxZmKwr0dF2OWBqUm3Zqv3mjQ/28wN7ey
N6vRVRbVw7XrpvOnrwG6PofZUlR5ULx9Z++TfLN5L5rK0lHlGuXWn+4j95pt+ai+4lcWjBZQNoBg
4FttAocW2O+GIWwcKLL4Kqwq1lwDlXb6TxrOhgkFfboQkloZfX4wiT5uww8Q2CiZsRfqFWHwojof
xwbDl/z3mQk9TThplr/QHNqsvVMOrPSuyLUl/NPcddwAbf3R6zSLybvBiWnvcrYqEPlSi4qDSxaC
r8pajIjFaI70Nc/3xBgQsjBRcfCAfNsmC6CAZRQcUQARFuBg6Kuj184DCT+2QciyZCbcWZx+rM58
7TD0KHLCQ7cPEFrgP6X+7SrHquNrYlR7HC4blydRLG6XbFYikBSkUGuLyMSJBkl+cz4FcZhpbAD3
L3J5pDcPaSQOd5LB4DfsxveRT0iwJLBQnz2tBRPWMdnbv6ZVmmhDR1Ex32W3iAJiFRI5McJflNmO
5S3kl5/8Gxk9u025G2Qauk7uX2xHBo8cnvF5aEe1ePlBOUOSknYDqI80/wKKlH0xAlyTpoklNIZF
IFuhaiU4Wj+TqNKp8i4eggJg8CdHkaVobczqEL/SULobDsfzHtr9NwaSDwhFnw0i6YrP5OGR6fBT
JW6O0Y7F8Rep+QxPOICOLuv3swbbfdqxT0YdgGenroZbPVRGHqPeSEV0xSwDcEsimnFp6WSwTpEs
uSg+Hontip2d8cMop9HwPybEGH0T9I/UWHfja12MfVsIHOTkdZtuRt75Ai9f7fuaDs/C+TiYItKO
z9nTqN/Ye57d3s8+guTIQYUIf+YE1XDdWxklibTzdCgiX0KmZ9AeLw5Tr+DWxK0oGbWPYWnGfm6l
XlofXoaiwJF64Ew8ZQIOem5AvzKPnqcoqGj5Ux/cZVMeTTpuOsdm+Pl5lJAGarIoyDlCAVOjolGk
oDLz3i6nJRsgIu1cHzxS2ELITSL7ZK7255fAf6B1hgaU8ubPXhmMzdYSsFPkW6GK5IIU7yMyBhzx
dzB2rWQsd02YWBLFpSTJDFqra/fQRqwhuy7gIWXEGuy0YNvkSlCm8Yi7FVyJ9ycLgTK5nyys8sF1
bAhJOT1gREDH9jQaVqt7dz3Cflayjq5FsrCe1I5w9CbrJIay/sMoWWfoeNkkXoufb34FuCX65/bt
afpkIaAMfczOxlVcVn49MSiDw7+RErb34XWOU8Qb4aXA3UQ33UAVi6wxz+xSJsLvB4/N7k3DDind
J48DP6g9VhFLEWf3XELl/WZytg6QqKmjCaajVYczf9mEX/c4NnQyDnL5zC6Ro64PaGn8+J05PZRC
oom33LAIImbqvCvDhOPEznRHAWf86Qn+s2P578Qrw0Nrf8Cs0m28vevvCSXEbjRqg4+7psPZXgIu
4LWwshRTGHIoHdjTLVxlvWRp98Tup9EhlEbUlDevFmF0ajIYpPS8Pm5AGgGew1rl4o8sVdQ0lb4z
VEeiHwgMAQOQn0tiGDPnvAXFGfgOc++yvgqjjybDcGxgI9q80nL/8OUj5hnnrXrxh6+F3A343twE
7vuWctA17zwefNManZnQdTOeCDy1KvWYZD4CyUJyabcagMMNAPmRW7A/ankkRxZgB/1+mnop0qEY
hoeESpyaOVBM44UWdEVLO0KDzPjUvPv7aXDh499SBhF9DTF6/lzvJfULljRF+aYhdirC1ODFra2t
K7CpY/HUcbwKTc4XUP7OuYEet4q5LeDCwr15jdKhRos2ngk1Ni39r29lDEjQhhC/scx+dc0yt34I
jt3mGLszv2lROcDjxRq1hIGBGfXmE6Y8FTZ8460OTzNhIpo0xXLglZqwJvps6/vciqMeqj3ypM4Q
CXX9vvPFp7PqyE1LJ043PqeKdvaezAB1wZOhe4W+iCgCJK6mKVvSehHuLTJ0jmllfU/bsisKwmKt
hTxRxMwjIciZQdzvNokvFirNeqqMs6xlbd6gtiliELq/IeCK3cAgkgoPC6jCl6OIXNZ7fZm+QvBG
b8LrU1bBvkRQZagVBBdCAXdNbsIzbdvVEd/gbMVQZy4DqPx0dQADuWPxSnDPdlguOJEM+GM60gu0
MVyYqdpb3R6qeFsCySN2j7U7FXdy6vS1zscCotrRuyaJcHvUWdedKAOeuUkzHsnb9fcSmU1zOhUp
nXA70qr4VXXPdenBwDc8qu9g57asu3/e/giEs/cmaFsvvbJW5RDUbAKF/0jbEJkxQZttU1SwsWlW
q4j5bN4rpXO2TcNuf1e20G/EdxeoML+Wy3AVEWhoIdRDRSCGZBPDiChdF72EKXI+RX4ipLbmVtqP
sFY9mWK13U7P5R8V4hbgnqdfdhBceN7J/KnDZ9XkwiveZoJlT2dUG4jaOzq3VCicP9F0YcKCVUV8
LrWFd6r1QyJ1LCft1GSkC4svg1/qFQay2aFRsxhVjBb0eAfv1VF6WbvVebTpq5GqkQbc9xUCtucX
yHRxvi+is4b8F7Pj4RYhS7TugaBZwh06hy30+pQ/VGaBswuWeEqV7uc5i8r7ZPOLy3/Mc2Af3pjI
Gc486xrtVZOLG8xPvx8EhC1VpGB6JO/6EkPrTZwH9nXiYMjt0QQBNkHzWT7WlYe5gjFvsvLyOk5E
oFmBoOH4WguwSgPVKG6Tyn0cmDWNpOsXBDs9/nMT85IYSfVgG23E1gL0YD34nMhNkTE995afGhDG
ut+b0w3ynljV/nSBZk15TDk8IvEIBlbDRX6W7sG11wge8ZheQgb+V8XhIFBn1yA4vv1jQ/eOA761
LOEgDL1qDikQhw+JBSVZUoQexWpOW1s0ZWNfiyviJyuI9O6AG/vPiPpEIBK0QCRoY/8I8Obwmuc3
WP2m3Y+nqvn+9MqEycIY2kaWgdvRnc7zupJabo919YReihlVlwetIBIzcrB2eRzePe/AnZGZer0B
z5r49RIyeqzRySjQXVwD+SKEVEHXeS4owivrSOBkadggLRw1niI3SbuCmgoztxSJgw38Mq5poSGS
vIJUizSbaabgxWrDIjv4z++Vp/M5WonK/M3ZHEaO2h3Q9v+KBf/1HEi83WAIXIZelwewoFPauvIX
4o8ltuYv2EEhTbIC9KEkIVR1K5L38Hscj39utr5NKkVWiVdfJX85wQ1GYD6CA4Gt93y4hnD2gpAz
DQCPABmGDeTgtGBWwOe4aJ2OdUpcVig7p3v8IeD5ws+JD5tqHv8vaSAKaf5lyEGkLv6OGYDGX3Oa
EL7LQ0bxtni0xnqzer/rEwWltKm5Io7qYLfhfGn42FwLNy7kS20fW7bLqWfl2Rdxl7wipPT8hzIx
0FXPAP/W+/yjuKD6BiFspltySlqLpbGRdUz7IgqyEG1ic4S3N8mlSqlIFcmasaHBCzt/Vohc6dyh
FWhdAsXElEwuhKvQVTzd7v6i7jfqUYVPU8rySQn2Ze03maw/wTsCYDIhP2wSpxyWHHid5Y7tm7Xn
hUmqBx2caZgtxxcvV/wg2BtgIBCfo6lIVn7ngjMDFsG4I4mobHVrEnuKxmCrvC4J+Y2EIxCzBIld
vMJsu4FhvlauBxy8s+wC/nM7giXfTo6plyhAIA3dkRNTsFxZbMoTQg8CCKHMAqaREfz9gvYQu1Wo
IkEvk2vvo0PjBoxiYt1OnQjtCnSODXNWqDNfA85GW8Zp9rQe9atXXlCJwl54iWGHJ7NMqF1pC2g2
rRE/GLSDjusiZY8eeqWrSWbQV1T0LNm4mu9hSuu5s2MVQ5A8gX55RPnVQcH87evRbsXUnW0EnjwV
wg9EA0NaD7aZ6neIFiREYFbZDOibaDhpy3UgHJo++7yCz3kmv1dq1A94uUOS1/+B4k2boeUdUpgp
nhj02CpWjZ6ddT6/akhLrshroux5kDx2iGaWXuTf6i6SJ2SK75mu+8BG8cLM0AqKHvaqDHdq0Sc0
f6aisTFM3Ns7JiVnUXuzg1X5xzl0AeDVZwIC0cUm/jaR+WKs84yq6CnaAxbWViofKtzAH8vqCQB8
KbWOKmBp3xcvut9J9Zrlrzal8rrp5cROxkfMh2WImr9N8RnAfHb4hcPXzwDmwvqFnTlMU1QwPGJW
6R7X8fBXzf/M/uw7/rPKFS7f0mO2e7KMQR6VrLix3dsMtUyqvYfxS+J2YjgTj6Q+VSwO25L1Psch
xyKGcbRUpETlKiOlI3tpES2jmSlPUeLPFyY5i85u8Oe3BE4yl5yH9eyuZF104rVL/PZPQaEdBDve
+68c0SXlLBQ8t3PG+o4EJbd8Yd2N0WntfPAPnUhov8s1dIPIdJFqLD2CBkYXDwe+wPioGQTg92I9
UR3PgVr3AArII9ebHWoO58feajVPogGe0ywazvq9b45WDgcY+HdLHruF0AEY9LG8w3WRl/z/dmZC
oyXFjpok3AIBZhufP8C2KJzzaKSrlmMJwgN0WHuIrjDRz6aTfxlNCKQdmPUxkijajZlTzpQ51iyz
eWho4uiKpjd3Sh9NdYAv/MIZmURHkfklJDmgfeTZ6gO2/kmS1PKkiHDiTY3M4FSERBAUmNHHFcet
32svGAWHszUU56lM3uU0oBfoZCipJzlaNG2XBnFzKjjcOErZXZA0VQ/+LSeM+tyxIeGdiZbNThBi
Alv56zr66AYFcs7cdvv1thmYvmYJMEp+G6Aq80ILmvHwmQ/Lo1lo4wxvVvUdmf+HqixKQ8aS5gx+
TPeLeD5qEOI3fdeyPIyBYH8HsXL10NSoEByXV/IRW2+ppUyyVbgRWvyxCaCXg0pP3a70sApT8EWp
qUr9v1R8YdRC0Ubaz9/grGgxckRkrtbwn2vuxjSYhGIOYhTTK28tZAlk3xAeKeSoYqXdh+ZXgddl
iGaDzOivc9wNbdxTJ4004LZV4VAAcBZfK2JYl+wbcthnlfsQVi42FYJ1o6v5PtYX7HgKDDBxh5j/
1WRTsMVep2ruky7jg4FkdXjkDk8p8zTcOiNKUFO5vac7lYjGTuIHdTef0KdCmOqdRYXESCLl2ti8
CP/UHhqSohEpni3h00qhaVLBMtohrMw3cWrnvGpM6/jtk+DlRNthjXfuh7Pw3NMf90HPUriyOS6U
dryrODevvfBFpFsqFvwL/mXIlcC8R8Gbxmo89URf4ZDpnpgp3mt4uPTJ9jjncf9oKX8eZUETKxHF
Qt4rE2D+Kwwq/w3DnU8u/Qdc4o851y+PQKRG4ujggH29W0o8p2rsq2EVAxAm2AGWGRTeL1Jpzg8z
qjkhxoWVP72kV1CyIfkOgAfHib6ySUmq3CGu4bsWxrQkVXLqjQzi4uAMAAtry3xldBzB3jAKpQb2
3ISprJRKUNnm/oaRH2yxySFTdjqx0Ved2FUE4vbLQyZyXl/hiNWQpUv72Ygfaml1jV0L2plaQeHe
4U9ajHKbIDoZMc6Mk962STxmn20/qOVlbdSBqUPwz3QxBRhmikMvlDNTMiv+Z+XCl/n6RJyxUgQs
JmITWNjm1x8hhmM51hafFBqd5AZXB7NtvWT7GJ1M3ICflMdoyQjQ3HPLH4L4BQCTqnwT796wtCVD
yi3pDoJ8C3uUd78U/yW0eBa1Fa8B8G8a6SfhFFKxmO6B/BkJ0GaT0WbKpnIrt0T0/6pYR9dPW12a
j0S5DAwx6gzGi07z2FSXLGcABPTIm0oJKNVLICpZtqtTRjoMPGRDNXgCWP0m7dPr/U6IQOyF48sc
K8WHk3IbT0BdKxIKmRxt5KMq4B9YpErsk1KR1YYX6+IjtjJNIlA7gwg8pRiUYpDMh43cJWvZNAoS
qPtTD/ERZzJNjlhPJ8CnK7e4QDXmT1fqwzVCF1/i2exrEh3VLQWBp3ve393Pjn6aghRX1HSe1qbp
FSut8wN3bv7RaRqQHmMaURQsq9bOKa8rO7FVDYZOVAPc9kZHb+xBoH4bakQCl3MnSNvQQCYz3sT/
qZmxf0eA6bK+w4Xf6nuWZH0N4Jy4dbvlmsDcCSKyddhXooMfB8Ux4DZyfNOzCJlmTQfmRvNRKhh8
hJB0KnvB8US22alZAKJXw4mB3OFuRfrdXGrBExmlC7kiCtvcB+bHoKpZ1GDDWyGBqIrPWtJGlney
qTC7sI0gBwbfeLw2AmEtRFQpFU13scpsTyBaJrLTvqTnq41Rnutr9UPewC1/mK3flLh/wSBItyGy
ABTUIM6AloIAPOKYVVIL5fg00/N2YqbYj88jU3RanwoZiimT54RptKoSKiDaZDQBVCuQkT5++Nj4
pM3vOOxz3+o+/vwhpkFejYoqZuSqw9r/gGSjvYY6DGAIwgCBQMTDUVes9nNXJ1XUQAcsU2AZ7Zff
euiRsiB/tZQ+0c6njH34DTySZ7kvIXBEVdrnzojJ2aFtZHKGhElwiMW9WCdBOVIBiqaYUH+SUgBW
PfQ05lIT1aITFq+j+JNOjPOC+qzcs1hyR88JY0xdGOwJSny8l81vn6JFg3mX97sJVI2w25lqtqQ2
WkpyhA4reyZtI2voBW1FgRB522jD5kiZZDDLEwPq0/bNbmBhCLFgYfw9PXI+xPVdZ7eBGyect5Nm
Yicbu3QNswNJq+OdwrxDGA645WjkzzE2ZmchoVScsjZ31TpdaYLfUSlLeLQ15GgBkNiuliTGnhpU
ML/TtKrNnH57w/LAifwa2O4ZbU5aiYZWjO8xNqq8dJxuBOHwIJfoFXS0p9RPdltFNVdRsl7uIveA
zXNIAaTxhFLkXX5Llbe7tfCOH7U15JsyAvN/1cQw7StIqhC2COsg7gT1yBlyKlL+VIRtDQttCJwd
2AV4Qg8w3PPYQbJeFY/XAUIH50NXBD+DWsquRMMP0ycplMkd/2DctAiLNUargryDCa5m34QFQum1
fOqWunyCKH6opETeCdxzxXGeZkU9DQOhvrA8DEffvPrqa9FvqkABkwywJJaMpjPNIBMcRvP7KsQM
oDAMdFzviBhQOhXj8XIHeB+6BP92RhGq25QvzQlaCJj0ToKjRgs6yPaLhGhUOWSFOCLpBSB0un9v
i6XijiChba40Rhn2PtavXD0QuUP9Td5FNs+4xX6qy4gxaFXvfguQ7ufC1vlc+A1JIa0BAMUReuFF
sB9r5Owa36vGbSgK4DmMMt8TrhvmfSyulXUQaU0EbNjNSXP/siM5CzIEeBe8OaChl6SbTc+9TvBy
so9r8Eg9y9BM7zAAhd618E7qehy95kwYiXdffnIuhPKoi6NJj9Lnfdw+kYRYu5AMG4spn/byi9CK
YPRnZm7n6j0Boa33xz2E052UtahGrRrGjlfbRvHtK5FBoa9i9grr3j8GoiyefNZOGiFH5QoyGEay
XUQcFR6y+2QXaDfdYObCXxaMOTPlKn+1zIvZ2tD7k8CZbThyWdwCoW/AVWk6e1RaWzby2RJWbeND
PZaokHJNEBEc2pV6PZi3Dvu//KRCHncSUoRRa4lTmoyG4ItYHi92OdlLJO5CRgtwEvse/UPI4zpN
k5DvrBH9PRCYYtZjjwhDz+058g+ZDiysS7XfbQg7YwTYnQO+BnzkHdt/F+xhSRhzH9xjLI9BkR/i
cKl75wKaRdNV9DpJ7qYbDB94Frk1WSfT9dXa5wzmxRh/BQaV6ZX4w/9sa3PzCin9XZDdFX/x2Rk1
wnJrj2FQourbXH22C77JaM2df8TFEYXMiR1KOeiZl/skUN6gFd11d5/Gxoe6hohVUjUlpPFN6wko
Px+FMKHRW2BCUohxojsyF137kJhPkVra3QjvTCaX0GBwsx+/lfXfR0TUyxpGt/2xYsWQ2yfjXxh6
8MSqiIuze65fcrT3R0FoYwNYRAqzUqaC7SEz0IyQUZcr1Lh5KzGhh99QSYYv7uCpofGc4+MPyis8
YmkF1Ff71THnb9tmJkfBfNlVfY6j5psmcFKNK8v3ST0L2TH6LTdHB6Hiusdv4sDHFW/xdUE7YQ4K
WayaPcprv2CbYYoZnivW8OjtQJ2YjFUyNQ4J1mkSh8ui2x8dQvR3Nj+LDPbL7NPHGY2NYVRXWKxc
b8+EBdvtmggvbl7Sa0fpCy+JNXFm9+xx30PM2tuVbbzqs8I5I7IzSh2f7ErDCVkPfaVlLgquKKB1
M1MpUjPMQ5Ewb0YKUET8eJaNDo+hjt5ivCWKw2vDEADqt1u5ePwVPHnKLsCy2J/fkyOOzZYXyiR8
ipSTDwIW4H6Vtke6gCIalGB9FZ00+LjdY6iqyvmklk/J8WiwyLrEV3Cq+ZiToYqFMee2sjU+lrO1
Y2rdbDIblVEFGQILU97I4MC8nW/pdixIkwI4xscdoQVDC7sg6uRd2uhha7dP/jF9UAIIdkzO1dAQ
cQcBiahiwlCqppGk9FPgo2iv0/KBPu5rzD6K8KgqtmY8TL94hD+tANbz0cMWCwfuxIniCsE8eLeZ
DXgvlJX2wcOINy7/mCKePEREj5//aGHgo1A76xlNtHSWeuy7R2284GMH4hrwN+x1Lcr0BSEUjOk5
niT7FyH6Go+oeQLls4hh88eMGqORVjrZxUOfsDaGsRkLT5BkqgR0oF/W/SLs2VveuBL9WVPnIJYg
n5ZOud1QpYTYQwIXF61zg/PP6FjyNq4ah67MjO1vEw+uLTL/rAsSIZCHuCFuthMQeqscz3LF1SS5
imQTw4KyudbnKHDFBungsFs1mddtDEWGUn8dJh7Rj5EARfxKjl4/eXt/g3So2T0ujSHtLghoy6OJ
Rr9+khAgEvP4JvCZdfL6pCVMlRl9VqntrgJgR8i81LWOSkLeeo+by82tfIMwVtng7Ch+pdlyb1Rg
g6qrWz8kZCMiAdGs+CYfvN/aYyIDFUrVnZ20XrJ57jjXFCwMV7YaOZ76TRGcV9C5YmApTMDfxU67
zXfYqFbcajLZaYS4JRAuORHD4fEsFX4lXGz1bYM+Qj9A68HqQDv2lNY1u5SXEcfD7wNGkRry1KaM
5f3HSSZgpgFNRjTS729o9wVxzX931Whr2IgJ5IlLSo6jdXfaiwlFuTZJj6jhNByda5BH1NQomBxm
sp7S4LFzq4kXC1Ppv3Bc7dd++ZEOBSw/pq4x6g7fVKJZH9XaTl44FfSJ7x6XZaufimhuctSOP8qu
R+nnCh67awpcXZ8oxrPlLXSxKnAH8voFwnRrEHTHuKHOdshtTAMRw4d3o4ULjTCkUju0wipOJWOA
uB8O2Pzh58qs5jITQ2LCLhPownVCl7OaIXYVOxrq6yeOymh1XJDmOmMj0UQ4bu/Yi1GP29rIY2Ba
NW/ltEpaEjBa/td32xdK4Dvw2pX5z58a76404Q37C5/uJ6FTdhPfbU6BAgObb+hVs7kLE7yw/OLI
xen69Nneu4tYblwX3Bq/WH3cbQDGJz7i5fHMrZGDrG0/397HH5W5PZdmiw27qwvdzGWjymL3wPXM
yqmtnALTDOmuiwdQEX/CL21+jubsgyubcxB2H1RlmFtsquFVwVlxIoHJgKTc4Q/Mv6IU/JQI1TgI
V+4Uqv4/e3RyF32o5Xu5zx8/42fbY9xX33I4JooO29006heC5ddeU3hBONBiyn+aUqBI5iFadmR0
bN83q5y8E0aLB6AqYIfHby0VvIGW3jRdzi6bdLAc66WShRZvOOJOfgsrlWtoOLsCl/eAc+vt3aB0
gqOlT9Isw3tMqb/6sE2gS4B45RuAxz6ynY6RFvC9qkmps6vw7HccFUJpXBB/ETd15Exw1zESfdDW
9AMzlGjyvz82q8osjOupzCdTYAsAGXQ1WiULwT38SFMw8XuGXNkXNqK2jLNx9ZQ6o8rcn5ny5T1a
RAINbAy6V3DmUi97d4SYVC+N6QRGjW4piT2v047AX/Xvan+h9Y9H1YF8pCDCzHHQjN3ZAO3gGqRd
/1u9PwEpep+Ic6oCnwWIHINyEspxqlNbUfSbJvFB9jbEgAl5asfmUxGHbxpepDY0HwRlaRPu/sC3
5ciq/D6f069N3KAmWEx92mESvg4acjcIgka8ZaNCIBPLEeIslF/DdQtmRH4gNWOFnIigaxAg1VJW
8JaE4O7YBzHmpJJLwTiw7Zd7XPRUM9UUYvNzIDOyYaJrYOLTiMjbUhjRjIqHfoAGbTfAZoSgXco5
zd+Y32qIdHHIKnugkdPfv214JmgUzjZ0WyYpdA9cJhW8rD02ix66beRxH3CthhAM6n/IDFfJ/vju
oJ/VWN0N3Pomcr0ZvD40/cdKn8ak3j+Rtq4t2qZrp1iaQ5sTL1kR+CkIgBa9E2lwFPbIKKvzg3lp
+M9q54GakfzAENr44EOvFSdfhQ5G7r4BT/djcknVdVRSt9WmcHzEZMgrl0JwQCokYxgZQpNOjAo5
ZYEcr4eyBWI5q6wiKxaUKU98GOgkymxmjFVw70JGxPgrEC3mxJ30xITFOa/jMqeOnuP/wmqdyySl
Bosw1aj4G35J9spEHr4As3S0+Fu1AfUzqE49k7EmF+mWjbERDBFWyc5iPle5LlbeTTu+zQs09Fjw
dH7mOpr8UZ9/eho+KiOR74/cxOY/WrBnz7DSsbjW2nL4IkcNEu/+5GhCH60NLyzBXt6XGkjPamEB
5WjoJrl9/lZqkd8UhFFM+sG9sSTq4DVdif/8r3xqNjIcbDEM8W0fG5s3IlxT2X4uNmnQWgnBsDcX
xR4V1Wzz7hf9gWqPjJ9/TO0Gk5F8I60Qs/X7aucGcq9MFzDk4hig9RVb6SgqcAd5eWEiFEd2gk7m
WzB+pg4oPGEN6jKwxaQ1z7tA/7SGfb8P9Mq6JcJgG6p3ln5g2BefE0oSDytcg0qIKhZdAX3bD6g2
vNuQCkX+IRwJGVHqsAjiE8xHeZT2GGw+HaWnZ+oUT2DMkKekULtOXrDgglO/03QzS4OEV9lC1Zbl
OC8LmxG9QeoBR/ZkCqW4yq67r10ujUSNg/2S9ZY6YoBU12vgtGki8mOV8Z2I7p1byyWNh9w9LBV6
MkDY+b8AW5/0ar2yVvcJpS5W/yIOQzb+sqUokw4FOkampU5k1vJxsOto4pzDeLw78m6X5e5Qdq9D
byE8x9WXxdfde+vP+1ebpdaXKCRickHZroocfj0yp4pGgFiXgDalIsS1bIehfSGur7dRrQu+I9Nc
ehmP1kMaGrqyaTiE4XWIecT+ZztK8qchkDswn/oYel0TpZJ1mGA3taKMY/++tvf8A3l6qdeyHbJ1
C7LNR7uPRSNnq74VtovITPuev/3h+Ir114ecLoLk86bb4zhG74kSmOUqFrjYGI5ylN8rhTy7tq61
iWgAGEr0GbQJXytcO21DEHNG0esE3vFLxhMcvXiq6KvhAgVCo2Bqw2o4OMPWSQADM9KW5JvIKgkt
H70OBELbZoOpkW1U6mXF72hcpEwICbwZGSjE555rirXjEQJ34aBKA4AtY1JtYyN8IxHFsyOKpUxE
yKlPC3tRQYLLoAo7uQ/TpQVxwrTgMs6/P4WTrFJTyoimGSoOMlnF8lug+b9SsK7TcoUL0z4vDbmq
xu7+URlmtUTSU9+Vlg3H/HF+N6u2k1wOvn6jxB0U4qtnI27IUIgB3QSwlg0y7RI/yl7fD1QXHcl6
b4/4Ub1lD83n7ngd/zybJIj54M5alXxsBPuNP4iwjbt2Kw5oT+zzWh+VedmJiA2/oH5KfgCRZmV1
+U1qsBgDE+2Z9XKZ6OhbWz5/90ZJO2/U5UbdAP9XnEbsvhkYFzRCNR47d9LljVirE8L1nSvNoOGm
h0XxgqT++lLdbnMeyMMK07YOK/tkCrF3StCboHQ9AuBQOYtt1kCkPGdfIteHizrt3305TTo2ocfJ
uOY0IQaZ3RejVrpo+/+d+zYcQ5aLTQBOwi9Un5aHw140j9Bge4fQXYoxgIpW4oIrJqkMkR/CatXD
pXPtUPB2cykDPrkxYdggiCIuix00SFJhmwxjU/i3EFvtsjWsQUFVE0dup02Dmn9EZ0EhmVLBLe+U
9JBKD+r2J0Q4wWXMnAaxHEzzckwEubjS8gRcZDjUeX+GalGQPAsZ1PCXNKLB9Jvc3uOZNbIC9S+z
Rw9J3M41k6qUzfAveUUoOxTwyx97KBxSwBqf/j1gFn4tLICG+dykNn4Bxp8+AQwGSBSp3KubNra6
tIGhXNkk3WzAzZSc6Ycl2Q3/jggSznGCXkDabCWbNurYmIzJQ9xoN4wesrNdxI/QaXl+PEnHM6NL
pjDygi/ypf/R4ksmRVrB1st/uyjVOAXvYDy8+ldVzGsaWKcJry2/rUSjKO9nf0/ARKtkFOxMcNPG
8Qij//5eeM/i9fH7FPkPNsQxkcdeNyBX/3DGa+e1sRxQjU0LbzaWkK1l4nO8A23rbA33PtNPfdUj
/aRMhj0wCp5QDJnTik18nYJYDDM4A4HbFmP1ASdOvI/uUO/XWofYE95eULSvY4Bp1+JPsrUF8vTZ
ew8kzTQgTzbh3VJg1dwCv2enjoVHgN4WNowW6r7phgTcr6AOFu1HMM1kak24g6MOvUaPxgpxtd13
LGBJKK4T7V9CMFAUOnshUIj7iw711e8rCgrmHGdqsuK/ETP/wi3tl3gP3foSBikX9ljnOyfb3qjv
rFV3jAjFWFbFJ/2j2Oc6GJlePI4xCmG+/fqjNhhIPxHqkBB+h5RhztXnhK/IFbvUima6CJrxUQwd
c0e4dSqkDrSWO27OZtnWVAvm7CSw7rOUYAOtt6L9dPjvhDNIUx6u9ACk8zuX3IxMe+TfmoYoSeE/
dlqoOv+ISIZOobfUmUekgCxbgQZgZGZ96erWPvPHDdxT/gNG7xcRJswf6+ZNteqPrLX/Z86KQLTf
Y/6J752FBNY7uUQj+0YxukX/j6Rosdx3PPjNQS9Yf5yjV4GpEGPkR30gXzMXXXoYS2b1+Xi4Z5jw
su2+RP0PeeWNS/eUuvCvw2UFz2B+R87VFP3PKbPwNsEctmhG9GjoqpMnQJMKeBreyNI2zrtzMh7b
1+LSgn8WQLqb1Z+coW4Q67y9x2FD+JdN2Cv3CZD+BueuATUXEwfRFknGgpa0dzX5BjAiewqQDabF
ypFDg+TRseVAzFpTSlDG42j92b6lfFGxCDKt+vHVpFXAVW2w8o3FTfCQgDXkNs05mq1QZ9w/Zzzx
qIWhzVpBB6FMMfaHhY8/BUbGK61V0NUjs5Gb+ew+TZnFdzc2mT2y3qiUS4vm5nwd+90UM0JSYikg
dC6tKYwdcuyL7w/VCqKE0qKZ02ggr4ezY72oHlTfWbM8WMZYOnj14LiM1LD2h9iACz5Mb4qdPyWI
NS/8SzfDZ7JjzXztnnbBBv30Iv7mn0n5IAHSqbAWvFKvjxc5KRGb3fqhw/R96egiIBsZ3JsKfAZO
wxzJq3xG4a7H6jAvVGDnbkxvXkJ/VSzmWUrhyqctFDB9N9iomit0kPuaOY4VN/jClsS2nZcs9cis
cf9Rbmxk2q1ehv009aFgHVwKO3Jnmo/jk364LpXyZoThOYkGnqTPWSY4Ipmz0n0hoosoCc/n6zXi
kBK9xS3vmnf+gqMnkfiCv7y2QfKAtuqkM15azvK3tMZapVOYhp2i6y5HoGoQUkCzHyx7rsej/90L
JOqywhHH48bxPc82Lm8+36iT6kkv5jW/qMplGtDRP/kmc+ehw13m9Vql7CtDyQHTPJnm7I6WhM3V
mMq0lr6+sqiACbQjGWL/aOOb8O+22FP5Dt27I2JS60+jQ/1tcXSeSkezjmhEAYdhoRaSgT5pt+0b
9uXheGndHMGCRB0kBfvAbhfrHqNx/FfEZSDk0+6iKrJKQFSu/gI7KfyYtsA6K18GgirLfh/n+zme
2w7nBH0u2RpPneB6mBj51n/vqLlCMvOlwc5eI40ljC7DqJ2oClWC18/5rN+ujdLlMyAvKDQOh0W9
eC9op7xJlqSKxkLw/QSNkpmK7waOLhuvCIF/5bDbkMCWaaQwlVajCitIdF/dcFezsuYCg3Uyme+H
RZq8Yw2kwspZiDY3MmnNMOYdhEVU2AvcZKFSiU2Z9DC3rGksypF9+5aLZwltjq1VuzYqK7a7JWPi
OKuKFxoVf4xtIBGMUuQHhBgHDfEmMauzJ6bV3EBcWejMFbrZVtTzKZe6xLh+xSAsxO1CuazPYnXy
LTCQfARL7zaxfC7iXBJ1BrM7g6gBKGbPEyNbLUNkwIEW7EMcQkxvcP53cXvFcUeaZ0aIdVl7jwWA
cLYtTG7sIIKC0K7uZZisrmb+QgmvYxKyC58SyYa41fv3I8ARADV8cwNmSXYUvflwANNN8a03njoN
MCpxfccMA8W2HTheAEBdquT0j4RHjPeBi7BXag0lK4M/xIa3RJWedXiJThjaqYF3MO9u8ordlHpk
sLKlj5q15RAWuBypG//QhPoEWraam5SilLwpng/ns7t0z/aV1JE4DgVLxKzlgtxsVk8lPyHtDP+C
QyGKRDHwhjnW3v4ONMj2cDhahxKSPCOrb4fFX6VjmqKO/S7ssEtB6ozOunMoPTzx6M+e68zOsGfZ
L7som3kRuBg/tKprW+BAu/S/31iu8GvoV4i/8jS2pNKPrbTvG7CB9mK+ysiyMi9L9vtM0etqBxcI
8rX5p8MgssLn9vof83JZ5+N/ghZDvTeMAr+0MYUx6ZUoqAN8tX/ZkrX8b1jFF1KCHX+KWFoYTpSY
4kE/OggbVVwzfQi7TR1ToPp/z5zUynn8B4V1aJAU3nONSbKlJezV9sTKMThybaS2OOWAQR7hZnJA
AgHBDbVDSGumFHpD5DH/nOcvC2pMZCKRBsIawa4EkRSXFklBME53yWSSd2d35G4dk9yHlgjFx5yt
W+gKMyphdvFDdy/BZ6T0r1tlfcZX2La39x5rX7N+5c2IXotQzLuXso8wMETWJ1LX7qFncV9BIFsL
zD9kjf2JwwOM6e6WIRpiMDBKJ7St6RE92CCS8RolX+w6mS6AlAmKT7EWhW/N9ai/GQZtFPHYSaLc
rZt4N4a52PL84qjb7vXaXl0oMV1AwhGYjeIbOQ82fUgmNCaVRE7ZaW83k7lH2Z7Z5qKnNZAiWoOJ
tb5hElKUs2/e0SV/47ZgjWIwjlPa3wxbL56kghsKUidI9gCG5kXXDAJQlbhMdY3cHMAhQMrZG1Zr
uk7NpLKWnxCapQECRAeWgkchtj0twqgxgRP05QztsB4LGoCn82SHtITrI+V5dX90kczBP/N7KzO7
CRCScdQXwOdD+kqw+bQDBjoAETM3VTAyapcQqkmvr5jf8T6pie6FN2YLwvgWh5X8xb+3bGDHiLuA
XhSMyxawDhrfWS317UJoZgH5JW1Uu0NIFy7WeNyp/g2tX0mGtLdVDmbQqHhXhioZoWklfook61x3
oG6QGR1kEzRJi8w6v11Sjc4WJ7OkU8bNCaYp8M5sRTAfz/L9nPMZovXFzINqJb5C67SPKyePybB3
swQMF6hDmBYN8zDdR8co9ltVE3e8dRCmV4XfwF5Nb7BzZXbn4vG0PdYX8ECjiLAlYLosdOfQ6IcI
oQK655w/iZChbUJFDfTdgrJzmMdky7yuPf9WMByoJ8yF6EIiWHPCW4khX3TAfsCCvYDPHP36DCYS
KMBCpQlHNyJaTSnv88yFD/+g/vv6nEROxJQJH5YuQfIPLp/qcF/HNE8knlrTHAV9QDNAtgP9ijvQ
MM7vOMcYIorVO4QdUsI98umP8xy+p5Bz+XohzR+JsDrdN0wddEkaiw717Jw1QRTTT+UdQ5Uaqliq
lB5KOAxWYtXC1iuyQFIf7MwUJoGf391wwIkFBeuixXQVHOwB35qTTK3BTym2wkjYoC3BykG2H9cB
4ytdeXfqbZVvPpzbYg2AQbMID0XsCs3ILK7wT3CdHz6QYFsioEdxPWgAUtlo07DS+gvmgkwiD11t
IBy+aLkj0VohBbDVwXmAbns9Pu8/q2OR4CQITiqu17c5/5S951LQ4c+d34xSWyuR+Of3m9P6iIiz
dqNNc0j+fZDK3QPcPMQ9Q5eYTT5qC7N3YWJuJa1QmJ3A/+EzE92tAtd/1ekmLloSlCxttgw/JlZ5
PqWVc3PYlulBGyrhZ/niD3KNh8LWc0meRHarjuOWBS6LLVGeMA0EZUkefrvRKdkEAlBC5+ylI0zm
5WbG+T02EpEfluOsJMTWCXSJ5qSRkjuZyggX0wSwqCCiWDFRstmfxBHcQ6GonD5skEQspKSBCXwz
HYAp51ecBAszONepx6aI1MFlbgbsFxxPZzLsHf0DFVchbbdkXJn528yYjVWBnmtOldtp5oVUZ7sp
3nypFlbDrZBf6Um3Yd3MNIqvQPgQ3mmKR0pE7c8xTwYa5PU0vGFgjvOMI8tUmAceUbhi22jBsR/q
SK7/U+aKLoEgetZuMXl6zvcXxGeLetkbyV2xPX1ZL6hL08Bbj4aL2FWj2oivCv9Lwd/kNDxxMY22
SU9tJoAg8sbrslynMUZsyV5qCmUGrQZ7SYFwmR/cWkbXLIksGBOtbVq3cUx8V3I1u/CLKcDp/BnD
eHf6PL3RjYnyZHxHedCKx+z0z07jVcVoGUm4241SmfIZXMFRDQdrCJONkouEHxuaQxFaPyAWPv+M
8bNugowDLW/VvSAj51r0Ht5rLbol+M14Vc1iux2r25EPDz6G9unw4v3KStW6YdX4xcdxna1OgZD2
CyaOqb958Tn2JSbKSnRs4vScZJVXTlMmpeXfsUJEV/RBWcFq4sX141CR5gBtQzrFo87ZbUwH59II
mBvqaUoO78YV2UWhjj23lOBsqZHcBHHHH5jsrEk1d/4FFSIrF+O66IyUb683M/fNeZ2Try1bzAoh
TTX5jUduwvSoeUzZVXK+ezfqCRKHJFCbYtdUrpJVSxK6U7TwC2tpfbSqTGlkUWB8ZgXhZbbiLiku
n+xzhNMMVXWzP+/A8NckiXymt0aZSx0UhAKFAMDs0ZuDbj5JnDQ+c0QPQctZDqn+pVP1dwvZeiUz
o3FBS9oLTojkXSKISESKmdYT13bJdHI+5ccZDq8ZIMIhxtTMF2A9nHHvkJmsxd0iIS56YVD8Tv5W
yInGVldtIAHJ+C047lkS9y4TT67wwjNI29ZcF6/xsCWDuwbKZzcPqW6tpXWIti82cYKJeGHnQNye
K0cFrj737K8EeQKzvCVDmWUN0QlXyomBcQfYJWJ6wF4pBehdBJu+HnKGUw4i3glIpLyqcHHAhic0
4CxdGS4nqEfCiBC+7oHvfLhjuFwbVjfJZQ6ZeMfA3xVT+tHSzhv5iEYn6woxIVQ4giVbWG6Mse5w
l1d7S8eAoS0eg8WiQPqioSKREFj0cBKL9HyymEIkchG87YIPzxv/EO1LSxx9LxN5eey0PpZfFMoA
ic4Zd8d9OoZKbUOMPvXslDTYoSTUy18Ci9stbiwRoRKT/viWi1NfRwrqDZ/Pfx83sqa+/oGs3AkF
mMJ1hg9/C3LNbYTcSD03/CcvxZHzwKVTTdxqY72m/15NBrDrPE9WKJtiwDq5S89m9wId/RlApaQ1
BNye8XAazLp8wawQmJtbUJjwQICObBiopSDbqn6hDjFtC7DsAZr8h1f5LOUKUEmhXhspXh1Pzz8X
VECyrToTBuHLaC9FXEt/405Z4B0RwW0Z0Drq8v76N2Oy0D1hY9zEhPBIDJIGj09p8oEwKcprxZ03
bPzYdLyKSfwZsSGzEJFKcyIloqmhXlAYQUS1vZwsSS3iJbohzh4N7LDRXVoYbkRwq9Jj2c+SDsuA
Ze10s8jJOq7ENwDqqt+D2Yehpb0G11dAwjrukXInJzYCT9XNJhbfk9jUHUm2PI+uzMs+HiQoq0e+
QCE6MogTqN49948/AF3yqzGeT4dn6N/IE185HvExUbKFids7iS4F9t5w+pkZGXXlGqeW+ZnzLblh
EN9dXJ56Wwuz6h3OywBwLA6Wcf8JwOIK4gpqUUIRTkJo3Kta0GvjV+fi1R29iSwp1c/ZhlulJSLP
R0qeNHYUP/JrFV6wwhdPHx8RfWIrnMl0zb4p6YtkBYUcGskgZaFFgKY/xei227UnSYZDPFst/gae
4OD60BglIJ/N4caYsJyU0U31um0Mjxh3EgtmtpZuDQbI2TnEBVg4FDNVWHpmIhF8vlb5wz/XCJe+
oezu/D1f6BqPQDCn9Hnk3m27c8N+OlIwcsienHO5rCoBGBKyAem+DG05TsnHnacL9rpg6bRuHMkg
rJxSvsiHVLnaE05+jCZJQv3AEIrxY878+NkSaMQE+TlM3B3ngWoM9yzwOQweH3v/2Hwwi3PJ1AXo
AJD0YPzpRH8/ZjRgJ/xV9QtxEJTNF3fFznd0eaMR+D+6KDUMbVfsjPY5NzFGukayP6RoDMsY3eLO
qwruCB3xMmow8TVHIYGE39VBvQoVKxDMmT5UEhjMarQt/VI14kAqDyLKsCAfccemsZ3+0pQMkdqc
bBNWR98xyasH/NaVcKDPycYVBS8dh6IM/Bv66XrOLrg1edVCT+KG0xlYohubrEwtn2RfOv3U/ZeM
l1bKHPb0UmTRiexXl2niCE3R+sOPnlkAS1OygAHyPIYe4MSRb7YCXT7my6Rk25IFNkaaNa7TRd9k
I2Mn0vT3SQjMxizj1i+iW78iZWih697dvs0vMtIuYEk0FEQFfLvxx/yKf3bqRG9LuZZvcj32ux0l
WLZdJcSlbBkGxc6xYnd9B3LDqcIXDhzjEgbsJT2Orn38fGvGPuXLrBp7q56F0nj0G5yM3z54rVD3
ZYX361VuQYo6zIE7aCqR3qZ0fYh8a5SJk3biI1ctN/zk1k/gfvA3rLGhZfqnD/ho2wcU3nn6R4W/
AAEWqsbSrI3rAPs4cRv4Z+XvMmcduReVw39FE2q4e/r8pymWQGNGddQ2gFfhZYyIed2vBU5ev+yR
B+RCi71tTr8DvWG1BxGod4ebyEGVikbPUyIJV0IyDGVCVPtJCyAQix4S1lUOWFkPSMl3C1qagKEi
pRtuawbg8HromiK5djrlIVECx5VRLGTW4BxDh6BL9hY+LLZQ59Wkr51bYSZRXzqzwSZ0/MLf8C6c
asWYU3GXgKkvoy/+RQW7AvSU/oh/aXD5WwAqmBGUgH6P1CmSZrq4ZUk7UYs5pVXwfWGMnYFGDw3q
YB5KVrTmtoUw12jRAhN7wdW0T4MJF6Bvx0sPYgAZ/TKBUUSq1c9iTea37sbSPf/50XRXjMkjjgcl
BwCWQu1yHsMXMZNpv21H/bSDG2YHcyEU/h2Hgbzl7zayojBwGIOlAThDm8aAtCS5IzOlWynLslFd
V8sS7LSZsqHZJaJpaJg/1QL4U9TieSSITui39ow5pZWSECycwYCl6VUMDhSGBzyiNoS3A0yJRPGS
snVicy/OqyGuDJZ+GK3+cUhEydpM+vR2Dfi4zguI9zA/21RYSp0SUoFH+EQ2xVAds2SOIf0OBRDB
AsdeA11BYCxqUFT7Qph5wlKm2wzaZm4AyhqdrcjC96Szggawzdx+XPwCsPm13+/wzFegsJ/Jz3rE
Kfg5Vkgt8Dfv3Wt1Hn3Rr2139SJ3BmBUxII+yQpeRgZAnwzhOJO1Bc9tUAd/doJXjL9QiznqIxhf
ThE+owILkLtQ6qkrgOFUdqNeiMSVv0tBAXQNPQ0HhJWiwP+rgaPEzVRhPn8NRVvSTDrXEksAmdrd
rJklV2FsOwU5FmO6/XrULQmUztBVMAR/P8woODSuT2lMts6If0REcOc/4wRWP0oae12zXk2cgfxF
CXTHyM762+7w7JbpunnbTOXDoOGy9pdrOXbwdvYcWIgggaq0/LwGQQiYg34fT2o9azOpWQZ96LDj
GYWpB5tdesWHqRn9MqLHTHlhaHkgpmXJpHKBlsBZ8dcuVNOuDFqivtBHLAnJ+B50obbb+XIxuyW6
QCW2XB8NaOyDyGSdQKj7lDegRiMki0HrzWNSxCNeScYt60y9a+ggy+FcjWqQkUUiARQQAjDGxGo7
5jHOD1MGF2/TUrOIgZ/FIGmv5vu/1fxUnnnsPk3GhxTzsnYfkcWVI3ghiSKZw/AHE40bMiOn0WWU
xy8HrXoT71q1RKoU8UNi/GqfFZIdZntqpfRsUMFp9wtJD4ciq+00b3Ak2uWiGHvqDF1WxwpEsrVR
n5wS+tag8kqzThzR55hCQbFKGHjBEySJKnxBZoO6kkhZr8y+xzh3waX1ueVghZ9fYeDiQA2sb4E3
30HuiVX7fZAL6zBYuHLvQXtYfeNu1NSwkHHzZh3KK8pRkPcyi1SRyvy9arrYF+j2hWr80LzgmfOu
R91AbboVmemBQfS3PsV9sy6DuPMGtkZNESOCbsObo4EPi6bh43S11Xho8X2ErLEYjA8Hw87scPpr
HfvZ0oZ7tnjdx8aUzglxSPh7L5QhJAXSuYcOtnHkTh8iwWc7RwNf/nGqvudVhBnpEZZevk/oP1L1
o+ZWSTL41BySxJ/kC8Dbia5F2KzV671iwPGOusesiVS3HHr/BU5nwvl261A8E9tLpPUmf0gugShz
XSRsZOFxm8zJs2Rk4tS/gKYDi0k/D8g9IZ0C3e1QBMS074dn01XuuXD5W2GuGuKfIBl9zLAf1hzm
UcdwKVehlWN7uxUCegsF+pozlOWARO6leUraQM/o5kW2Ifi+CVnWMjFGyTKRoLhjG141nA3Q6Jft
na2U1JdAgSsgmBhm2K616X657aOmXP9WSptpLtzxe9yTBq+Rvegd61EuoUXAMLjXAdFo/fA81QqW
5o+/k50PA3/yp1BNBOLNefKGX2Bkz6DqROKJxQ74Y1coOYGaQdvQq2Jzg2ymbxo0l19413itNFsW
rSPUxhPJ9wTFtGZYAbBbhgOoW3ofgjoa6Hq9JkeiYDuB1F0M/jCH9vvS1Pe9h53ispTvMOI9ZiWY
9x3MQ6685QvqRxavEFF2gRvfiqp7606jp05IwfArPgnB+/8KjfZYZgjCUfFyzdDCp78BoE88Kty0
BcWTPQeXM9KKjLTPg8Yj9ZkPGsABknzkyPMId+afloYb61bSs1BcZWOlNHepigrnJyHVaDUqK17L
h2Z9UCQBLB/BBn2DXLNA1L/MxkgyqC62ng3ouKW+jUNKG2qDblu+zGcHkrhhn/t1C1PVH5m500fO
EbahKTcLK0+Ow4PbQDRqhU70B2L+Dm/NKcxmgy+kZL7xp+cjvhvS7M+5S0iYroNJxCZfUJkG51VN
1X0A5avz2+e69ktym1zlCvyrRm6yRNiRPLqBYDvsgA4f7eYjawbmjVEJHE1Fk0yVbUJZySDQpM2r
jmv6vya2EvetfomkgJG6hruhXQ2zKDqipYRZuOsmA4ZrtRgyqEdnoYku69so9uIOcU0x+kkP00Go
xz4kVCCuItZIv20kqyB5PGfzIiXA0OGijYI5WzqlzcDbrpQgpvgAYqRpCq+utPRoSoLUqsWW2n+g
uhhUAay+10X/Ai3dWCJRj3mOMUd/dFQ5+apIRoaejYmsQUOrlJ331UKNNFtaowwPI+6tJVIEAp7a
omlYoKdwLq+tuay5/Om19ESRibS0/a8tvioZ4tsYcV1a3aloBAPvtdTJsPUJHkgTC3AyXj7fSKDR
xFP8aBaIc4wX5R7QLQNf7LgHzaL6qqrjf9Z+UkJYOYiytf2lKameJCFoghncxjZh3Tv/KgaHjmK8
5EQlyB5N7Nj654w7dKuSFIOuLtOYZ3jesICCrY/Lze6XujClC/hOyiq5whMrxq3MWsI2YHfZZiWt
gD4T3wpHIhSU1IWGnPx7aADePzgGTQQqZUyLDEN9a7beKkZDma5kOTCKoyLDasMAz66/XlPKi5Zb
qyagSL47DV96K9tURQLdwtBhv5tg1l5752lHPSturWKfJ7354pHlYYwRiYOjJjGewqWpiBIoLI0x
b5z4jwx5DazRr+wpIOFg1xxwdTSQOBfblD9JrUxIOX8cbkrXhaYH5c0t2AOtBKOkid8YYhOtkTBY
/b/2ud8Hbl3IBsVEo0BLKoXQ5vGl3/YQHilT64VntEyno4wHkLLsAf9AUOjWvoNRB+TOiQlsra/b
R8UejmfsefXm123cnLa+YfPNYFojRaoVaQhkmOzt0bFv0OCRT7j6GbfMP1o+ntN19g536u3JLzxn
6Y8HjXLvys9kJeFQeNmNfjLh3xtwDhWTFTrsncSjg1SQaNSY2DB+XNH2RwJwo57c4B0maEpGFlL1
VlId4sjvD4Q8kcWNSJdYYYZtGqS345MjINiRglYWJfsI5HqMbeRH7u8si9KKOUIk/sYxnq5lnxKB
f/ZHTA/iM4nPgUQT2iVUYHD9EjHqhnb+ShZvBT3J+8qoJ2yRBi7jPWPh9wZas/HHBls3HfgYqGfD
zWk1+uh4G0Ck9WfsgHeguX1+gsz0khN/McYQN42NRInGPZgve+COu0mpypihGbYggXWCpDKJwD5C
vtlM2Yf6+By3rTa8bQJaE1jRxHVFqhITFVOFFL50SFgv9vKGJNYpG48XmcDgm4oB+EuTpP7JX45M
2wLgHvzdPRsEFc0vvFHaBoiPMHJzaos1m9E2uKRt4zqnsM2mQkW61YRhHpxj1NxXC+3x+FwfZ55B
YKt9cjb7VXtg2TTHZEjXzgmLMHoVLPX+T5w8jQ3atqdC/wRrUbTy6gTyyIEZhNzFtgOMFRlB3uQD
ULp69KljMmFZzw2jfZIH7GAVg+fckl9kH/qUawZUcXXLZLYwcXom14LtF8/F8UxO1vEgRelHCS+g
Z4hpyZnxwzVXT4yNbdwAvsIF/S7lLqJ+yBnW2exKjqafKtgZHP+PCfotvHk8x+Wo0+AkpcAsNpVB
xyeN0tBthMN8LCcI02bBTqQWsMGdFGCizwkuWcWeFYUmcnOGFAKW7ithLyLRq17OxLjC1onB/j8/
ITxc50zyj5hDgy5l+NA8bMLhMEDIiwxu9CZLYYCBnPUSRGubDa274keE7hutR9A3zyu1tD4q8Cam
++fYc5gTkAyYsMxRUPabeSiSrB32LlBGT8Asm6QaQP0mBuvWcjsWLCDi9Yr3faxVpqJ6pvCGYU21
xf2tkF5o79xhKwu/w29G125m0mqrlTv/JEWz/BrTWepXNAMEX0e+ZXL9/tnTx93+fYdCOoUfgTck
lwt7Ohv/vVX02+C++r1ddfvlglD1J7h2AuKlEqLjhK8KsZ7rFrM+aFKDtgtwIAj/J7cg1yM3DOii
h0kCaLQbLQ7f9UGsggfVPHNYyUbETViGbgDLEYqr6CryvujOUTjQkRzMxJsPIYq6vbOJS+DwdtZA
YWqaOZcgLSNqt9YNGnDhhmTZLvGDN6jLgXgkrswhvB9wwWVeFn1/9sGF7wvJCGuc8yn3TlE94tpF
i32yEwQnaGR+MSP7BTOcB6FhN51MZsMe/YA/VNAixWv9rGtew/ZJbGU0mpGSY6DEUTaReCk+5cem
QCuL1qO8zcham7EqIhV4hdSbZhgE4zzRUerGH7kB6uhKfKT+W46s7NXEl7aG8thUIxIzWdS1YcuK
0Ydlxep3GOndOfmhfC6ODk/MGhuZixIyc3UfkKf4LXUKgStJL44G3aRPKkGOPuNiqGJ+axgYhKZK
5xybnfX9oDxQR9Y6hOZOOa0ip0DD7gcF8eZAowcGHgQxThhFCkFlsFOZ3+xx5ai+fp953l/TihgO
O6vz64gqWZfdcLHSBsSrKEr3fgBhclnbInrBsVP7QF2fJ52B97kgkH9nyql8zc13CLL376FJkTqc
CfnqSWgyjRCvPz5agaElWUDAjE0VrIPaJfbmjRWcoRhDmD8/W3DulIpBbagyNsqfPc10lLxwIgFp
+4hyiWJk9BiI7/SjRK2QLnZOw606JcsESNWPeZewvWjWnmev0qeIFqnS8pi4i/T81p2jrE11FwBX
zCcfJU2gIaD34OO1UFSJVArI8otDLgNiaDcl1NafDJEndX9YENO1pibIJFCS26p8hCXwbt1Y8ndm
D+rX3dZyati2niXv9bhXRKgfcYuVMqDgKQCJXZ/qmyWWgFLpehm8FbOE2ThvDWDCm5hHVu6Pqk2T
XkNqccI8au8TYpFdWhxIRv5G4b2X2JyuQ731NwzUi1dipQgE36ZFNyhvMEYpTUCc/Hi4FYBOzB1u
vP/BwtSjy2vuRx6reiraefTASZWjqXUp4y808STWld3ZTLtqnpxkk5ZF9uj5+jDj/j+gUPb7CcCd
EekTJbOE/D+6kTKLVWRRDxhZdwvd9vWRNwjpZMr6+IKMGeNjefJfNDBdhkeMAhcxw6qoW75RcpbN
LdmuYtOR8q1G2sc73Ia6YyP9RSRwBCnXvnhdgV0eCK7oSU0lOZjSx5KpEdNarKR2b5hlF4Evc3QF
0wI40soaiLvo21ZvUxIVPJ9CTT2Xll9FoG+T7sFE+Q4vulAabSIooU6f1bO6Ks9oVaq/sK6LApZE
KsdlymVgv61pMAmsWt9tjBaSirzwFlZZ9QhHATo5A0o8tr/24BfKsPs5M+HoRa8ICCtdfs7oijjr
ETMvoocGVeRkhgVDlftGr/kS7qpvwgJMa/K5UZ7c+IzOoKcdwDbttA7l2upvFIPOfCAgdgduW0Ws
CZaiWszF/Kcd0rDOcx6BqnTg62dpXdRHrzzCTtRAbtZT6jfC5TkdWqN1gZ7ChW8zPmndgvR9bqRo
NJ+gAiXJX/p4rvvCsnHJ7J7kJPSZOWS7Db3h/hxkVHcPaCjDjzsjBwjr6EPF1Yv4mjbwkLd9aAhZ
lb8Xja5zf9ER+BfOP2xeXN0sdONBC0q3q5HPc6raa3PdULInt3KV3A1Sm4cOuc8oGWy9B6kihKvK
ZT6/TKM3CCTAAF26PNrOscRcTAdT2KBUmRr5UptFPr4KUAW2HcbGmtpFDKsUXipEplnnt6iCCG7f
VosLXT65CIx1zfD7ZRrKtyI7IqoGeFzwRxfgEodMCzmauGawKaaM6wqs6l3LQslRxuP17P4UBZV3
9LLiFylRrMrza6/eI2Q4WjLEXXDTu0qvSjhvjNka6NBsdUjcuGmxXyzC2fy9+Een+HdlhQNch87u
MO6X1zMbbdJ9Hm50zWp3Oz9c0GE5cbT8pVlh8Ml6M5efUuK1/ZuwwpyqNNo9ERXfJR86Pirink5c
icx1yqtvtRghSInA7qKFxVBb8wpm/KWYj7pyaDyAHIhyqs/XJ8CBZcvaL8CTmOCUnZ2c9IZV38yC
uWG/DmdqEvogEYyJW9gMsDdmuB+18gw3QV89fteZOtlTAA8tDM/i5Fjj+OaqXmHAVa17Y8VATR3P
PGocBWtO8fvfAbv9ncIn3SafhZgft+lRcgSLlVCGze5d+yMkLGw9j9SsVpg1hN7FRVus3B972oC8
ZI7S+A/vg2zKS/WgwAMu3mmEpowrbnxr3Emway4wiGH38iyWLG+wHwo5vrkWhcZEOZO6owayb5pm
CcMvkuI1GDiLNteg97iqMu0lKPheF7iL4+BLOV3MDBNyAT3Yvag7m3k+EamikGM7En25qzOzmrjl
MaKUajnyuZPAzLjgrtFlIE+iHEPCoVY7ZJiGdhQGhKwbv+oDyW1zgp9b01Qw9K/O2NXTwOhPjQYs
TtI1fRqcechD/BV2CLn7NQ7u0VmPg55EUegCtdAmrrEgaPxjYcRUft7uxtUwEPliTb4QkwJ25QSI
9UDNs1Ifh/voc60hZ0hgmG5HVaopRO/05njxGl0eI8m+moik7bGNIRqKU20NgPPnaHUcUiTWFoOX
0nW1OkotwRki49IkeGkmGj/IL/dMS7vc97cV6HmsfZ4LrjP8hJAROVZXHZhZzSQFb+9fA8VNvyij
J6mF7iBjoyexLIEGjOCNtoG/d1j+sK8FYy1ivcFgd2U58oYaLwUKbzxsnt4j0cKyiK9xck4/6kwI
DxbCIqIUNNp892N10pTdYdhuxiGjiiNatdmG8vk7/1sC0mK0dpyghhKjr4/BNYa2uSfAqHCuPVGC
Q/ttQG6pYvLlg7h4RCYJBSOtu/QIe0X7LWd2fuNQcNUR8Qr8STkw5wUDLV/8ReVpVHiq46TWxim6
DL1zy/xHAJ29IQsLwWZ+P23EwkyXdaGIJT4pQ30GzbEFlMtHhL8vWQQJnScMr3vp4+HHroyN4PW2
5mggLkNrbzxNBaEWYjMui4U9bpEFXJ5jfQPbVi1Kl39a92if/5T3WdDIGyddq7KAVHzShqXYcRMN
SjIsCNs2G6W5LbdTGxOd4px6SbTzQCnL+qgy72Isz1X6Ks5JXyXiaevd+t6e4nMK7fcwZeLojJpt
xLMeWRFlN8QF296t1Kwec0XUGZ4y02Wt++d1wFKGPA60UnU/v1bDL6R5BI2xP/URrIvZK6sDCAUf
Ebb8Ycs1ho2egmgmUVpybqGuiDUB4lqtqySTmd5olLpET2cpo68a0KbuRyx8R58NyxFSsraSPIXK
wKNK72GDcP/EqrBKmAmISukt8vtSyqGmfGko8twGy6JDi+twtSUq7/SVO8P7qpv5fya6nfyYNhzd
CsFfUEu2ri6LblhTYz9RkIQPMfKuv6HXmKIN0vB/LhlKTrqgRh13xl3R+ZFPSPqOpOfycO6Y0Qld
5sqpApUo0khePfduAdi68yN9SSireBfC1k7IBJIikC/uGdxZPmpeRUqCb0LkoH7aHhtFNfp5YSB+
qjHBmX+EKP/yubkIdsqezhsip4/wEefn0JsTCghyM2tnDrXxBQGeXqG+ZD/5Uco9XMnN091eZBhl
1/QpJNxw7QbuX/Ak/9uQCyb6oXnDClYAF9Z44a/ZfAQ8RrniiIX6RGE+ABoJvc4mNbnQXNMVH2zI
lq0lKwAE+6A+GEzvF/cesR6HjLgIjJZomLAkBPep0CBIY3fIn+lhk3NS+e0EvCMZe09yiHYmVTHC
gfNCkiLSRWSc7Ez4tjlxjXzs3yNTmi13aIQWDuLeHvGwZ9PCiNHWbQIqnGOh7Bay29jC0qTdSqC+
b5dz3e/4rkdD5U3kpwphSTEZWUz9mvuvcXsY7gpjKr6AAt+0sdZtUB2rRjE6eNhLu8+TY4pgq+C0
hv+bE8vvY+TYOmD2H5AY9J410Ufg8xcJXL4NmQlw4f0VbkJN8qtc7/tQGoTJBBmOgKwUmLRksyUj
J/x+OsxjkLwRRzCcwy377OJZgGvsjqF+FmWjUn2pBvSkJ8huGRPTc8FV3aba4T9mGkIn2ZdZizVA
Mkc7CHLF+vyEwK6IEr8Rvr3URk54zyJIUmXSI+VH1fxB6BL5Ajo8P2ySLcowCd/WNIOoMbJISUPw
uLChnNJHErApIbTWWLFGoio6aw8Vu/vbPYAWN42QkYCE/o/bfMOeOnlH1pwIYRFOIBCLVeIQGX/9
IjdZk3vY5ZdgJexd/3U+dZm7/sfm2Vn3lL2luvezckdZNe8IHjUqB2JA8j1grGPOBWKVSUkuzpeH
hLkBZMKtrycKlOr4e1CyRpemxtER0ZV0eWNIkLBw2zs3VD6Wnn+Pb6UdUAlbOpkPD9aNvuXd1WFT
BN8Vx0javgzlwbsvSrEnFSme79k6taBlmcRfTm86FVX1oA1ShSUSa3e1PVbX8J1sp9iy3JlkKENW
Ga5ISeszIoosvXsDzETDVQVzsHNdW+cTMnbkWsRxOIwkywjY54YV/eNQBvPD9EB6Y4Mb9jpzUR9D
/CXnMw8UGBmffTyZrT0+cYsWpWSgiSQXbLgTE4szkF0n7PUsnjGj0jV/W7fVq7aA0IvpUTWIcjBh
8PQzCd/dd3yJQQR+OIs6SZ8Q5vgJ7Q8XJnY+ImlbsTokfoxial1Xcedv592z0NUGMT3oTwTiNaBs
r1Vb2is9TbiA8+wFj8LkRuXs7mFlxcc7YgYp61zavw0y/sPAWsCB5wjoFxjrKcYZZ/3VVbg3Aaxi
ziJOzjm2fkj5C+nS+p0bEQfTyHerpzx5+14Jr6NNZaMuyt7mMBy1O6MuY6nTNR3AZKukoN7cGULy
vPpPO2umRGhdGAc0FaSQcDC/WBPsZ3umK88qtRoJ8cxHroflwebuwEBvgyYTlEZ5ZHp/ey3yTEQW
fImzVupkFEOnpnGhuVV/QXYoIdmJmQDfg4qsn8I9WbSvSD8TQ9okiRdCibWZer1jgp9v9cu5Uerl
+NzalBHospem6Mrinfo4vf2ADJne7N3eswtoivZ7IVc6XRDnZFW9/VJ4+qzNPavgGXdn0MEjkoR8
dwZnrjCCbQfdl/P/5JbbsJrxAAnvV8rJMGPZLaC4fPkt/67OHj33kLtVAKJwsqNum4L4ah/1Y5Cc
gIbimVssMADzB4YeP2pTVDUeEU6Rfaggon8XWt09q78y4SkoJHLYt1ItKLZMzn4g/ZbrLs0icudI
2dIvNoYI/jbWFLy/xQzurkPk5Vaw6xAAqDXXoHtEXZqUisaWMFJDQXPfcY1QbUtjuIBc+T0VwAwm
I79YLZrVGpjHpH/0Mna6Oa18B8J0BMXdldkpULRMgjvwcScQWN2Bhsay1bopRKqhcspsSqcBK1Tk
/dsuz8ys3VoApS2zNqHQVq0IGzBYloorOb8IPIVrlLVDb35lC9vP5pOoUzIjr14tBVm07lDsXox/
jl+01auq/opGivL7viDDEbM1ek/oHIDToVp1d54Fn55gntGDFlPBqORJt8f6tXkqWBs+KlhU1KV3
9swOOJLtZIhZM/O9wQzRfXqQyLHSQKFx+gJl4yRWUPCXH2mirbK3e6rTOGBMLJkYXCU14eW/c1lP
qHsmrKNZkMhLfPHh/0yMhhMAWIlztTDGszEZ7xU5JbGcGOyghMcewFuTbtcrVp8wmKGUnHJ28/g6
txdJxL4L3NevpMA0ZooENB0irw/pV1dE2eOz5mkfTLXHNlTqdKq+dGCpRArBgHe98lq8KYrXxUoT
aIx4lyy+QrqBSaSLu1XLVDCLoQyMT7uQujQmIUqWAWvarzB5XZw9bIKbf1o8x2IOHSrLBDy8vg5W
HYHL4P9molsO0UQGc7Nk5Al/bFucmrgH/5yR6BG/R5menKVib3zlIyS2Q7GiTfYpJ64MccGPE9sA
+yOwoyd6rBUONvHZpgiEHGo1AuiqYo66E9gmiXYRNU2Yz8/n9RK4algWObdjEk31cuUc3y/l2I2T
X8j4IiAFWzcLnvu/Py9xmJJd8+7woNuBD8JYU4Dnp8pMr87YkQwS232/94wdJpZfcmwyW3X3a4MJ
NeytETqrtE2PjFDzSrx3n9TN0sNTQKTS+mDWx1jhhuVHougHrUORN4+LCTZLx7IJwzCTTVjrw+S+
02iJtg/+OgJG+lc8a6bP9oVMv/X5Su6wavWFsKqaQuzof6L5cP/oyXvUlrZD+jMbJ3TVfWY5biC9
tMQ0id+5/0bNM/fYTotaBpdjPsnREWG6rWmk7IYP2N2wr6MNrtHkaiLWwKq442H6UuizgqA6GYEm
X46NtiBBUiQY7BA+/KlnjMcwgtrfjsRTw2h/rxyHy2i54l/fVjcL2CCzqMnraBrJp4zEXgcT+Vv3
o9KYWU4vGUn3qhuz9+4Tz7Sc3wkytaZ8kQmEvuuGErlKW3q4gElXmIE/sM3emTuYW8lMZyHdNCaA
71eRjSQ1VYD4j6kQ/peFh0Zk/c9jtfNnhYQXaaZ+2IwYY0KycGIr0ve8cjRd0KkDQ6xxjOweeQ+e
gEC0//xZFXhBjAWqGKTp6CZaIllabWZePY+X72WqoohIdvv2TtRv1hqbwaPaqDnWSMwTxKBxKFCb
j4aaI4+8U/ksMQtbKIQAWTgwWc/Kyu0z9QCCav6nmUf2IDWGURw5ZfRgMR2Wbb6eIIO3E8PlmH5F
txWBYKuutxXmMoLZd2Q7nNtirIb9oB2ZFlFtNcip2iMQJ4/2JUT7Sf3+1lhqcLlFBTiaGrBdWcTs
iEVI83FgylkhA5ON+dMTkY4Z4sXni1Qonj+NkiYG5qhm28j7HJ3yT4tfTFXLUYSZ044x7S3Rgbs7
1mzMUZkqBuK/SllL0EkJDVgBQGcyNYTpGlElWRttPSWk96UZKAuNFxGQQF6kOy2DPE6LtQXAasZY
NfCajv5GAwUL+J1PLZpgITNs68vVEW92ly8Y5ALFLRUHk3VH7T6AmPkV9LPsLcmXnyls8d5odRfb
I6+TSysAwPd4ZWXtTUnTq5wYFgyjvBfv0KhfZi1H3lgmjVnUvTxRfNEVmFcYyuH3hpsBoVGcgnzf
OCxQATJER7dsY0442zC2LKD9/AtFcjFYOdcFK6exQ78c/XbrsxL3ZiJNogGnJPfR4DiCKMbNIgFH
V3GWUvRZzJssNvfCmNWUnpm6wNnFb/nlugXPHZEaFn8HRfu8Av5yhK5omDWomYzJW93f2zpmW29w
EkfK1ixGwYzqv+xNXvGiTQyrJmqIx2y6NC13A3MAitgrjk9baN5mGsL1x8G4YKF0PlA3+VyYz9KJ
2Hgrqn6UXXwozVYe7x43ZaHxe3Xwzxd6wt1HEWhKrnLIzRK+CzlWCPFnzXd/K8enz8DGFru+ATLB
A9OWYDt9B+3tvjw7+FhpLs+XgqiQ25zVV0wItLEeKLrY3ziJxiTml74sY8Sh5noYG3WH+1Fh9s09
iHWqE4mlkJ8d1YfsUdfV+SiXDM2Su/xkqKQv8NiBIsb1QPx+egb3UI92d63J6yZiqAbjQVeBZu4B
caWVtEcLYt2OJpASyahVzXkBleQKHG2c7R2wI811HJGYEPzLaDnL/mU5WPvEj+LMsbA8y8ONnqRs
3NchKFRQKJsVHGFfLAhhw2i7KA3vQHsRDcVWGkgzRWjJan1VsTbVeCH97jaT0yFmI9253uMZImnK
+JR13Mk/4Sxy6HmuK+66kqIPW/+0KDejy9muIO5BOmNhIt0NJVyCitEuADuwZdPjfNb+DmCOS//t
1iQLyrgrSQrXidSInmSnrc5no7Ftk759q5bGjnKG1F22Ikk7oS02Hmea2DpA/JjzUo0adEAJ5wjy
JPuSIGGorni4yyFjtq7bctIDJMZavScUlNJ80vbXRxrnQfLGdZHY8SiB7dZndKDc8OOP7NxoDd5T
LsoOKcIoPnuWQiXOhQp8tKvC2FkXjlLhkBV7AXOtQhjk0a7qTWYHPaSdHB1eBfbw+ChDsP7R5ijp
f7UN5G0f02wWN4y66LxBXY2FI8N4woTy1tE1jYb5dLN5Hp1SqooBaAApSs/cG1YP0D3scSEDF0sG
Yu0LQRg6+h4NA2bGINDJQRtpPnw9C/5zfzVMUorCSYlr1oahcULuHnVILw71MZBw/Vnc2yPcQoly
cG8/BhRWICC/b+RZGV41X2/QO0wgI1tj16KV6B/vrCJWxmg22aJ+GwIv70wilop3OOj9HGoFWz+V
7DXKNy95/5Go24H2pzW/pLrbjjWtxJrbI1TgxVS+gomi+gy+NC5s4hvMuCBnknV07JKxECrk+r8A
Ijqn7/LvwVvnrol++Zw69fygW9ZkbopmxbAIFoyRc7PXObsDyqkLLEZ9Fu5cj/OqJ1xIgYRAU6gV
AqOTGeAgnmwF6JCaB6+caN6AyXbkgm3hj5kTsNYINxWV39MFdvTABpjfQPwbdlxCkZ+K2EF9tVX1
SUPaRBkx/nb55FtN6AxE9XceOisK6u5AhbdO+SIozQ3DXEy0QMPUad65qNIs9naz87H31/VaWMrG
+VjdQ1bPP4hxVpNxjCPv0XBRFydhk0goedQrFpNKWC7xDGj9V1JJcj2BOCKQlnoG7WKGMRrr1xWP
bUWTfpdcRePwPrSdEOCT8HntkU+YrUG5J5KZmkoxEK4VQ7mmf5yCzVKWI8zJiwq99pN85zK5WiT5
wDhEja6oAaAtYe0iuh3H57GPGHVFUZ+DY3jIMIDd3tntW0Lnqxdnib6UdG2DmiMUZ9+H60uh2QaG
viAtKW2TC0+DnPaN5PJYjAfHegNZqbQehzSAKCBODhp/8ISqQzoPtfFYjpqjb8817X1n9yKVljFZ
8YIJWWgKvqQzNI+0aSYCB/6OSeLQwTmlGCw3rMkr+r4V/pYRIxv8v9y0HC8EyNcPRApDtxGWHO/h
E4rAGrLsk74wEhZTRwxXitj37q54AmLvCVaLZ1qKoblCbwkZaZuyLtP7k4Te+9g+VhbOMjZFlEHE
54eIfk86cQXnsSw5lZu5IyBtmiDQII2OpSksZ6f+nWF7XLb+n1ql/qe0c78fouvnU1AOIfRxIh/u
ZQ9bIqQ+b6zUpGjrtD4V/h5ylvLuth5Wc7prPFOiPCtx+3O2SZzzID2Y21W0a96e5KPSrIud2zKd
Rsfpb2UaFgl3iBlLgaO2nwigSR2pUGWEDsjCGp3jGmFSf02lQc4oOKCwfUjEndvp86HAYzDCNQ1L
Z3LtL1h7N6fmRYmhF/s3z4GnPBTasBlXJCVnie1s7ICrQ4EbAnNIuD3SxhL5ogTBc2k/zOmTdLzB
jAq16UNjUpaFgWMXlbibGHxCNwhASDuf1+P/iQBUih+C2jTIim9GeC9SfjDRBsmC1VGdC7yhYOs7
ITu4RGS8ySOHHpBvK1TpD3OgLZlPc9FBipikaV0b47TWP+gnFjiDGp/34ueE/EifyLtt7jFM7Sz+
oN08iLf1ZAUesXYRJlJe+3CzJGDFwEgOYw1gVWW0E9Ojncs1cqofA76HE8INh5b1GDmNAWWYyhSt
BD+nWMprzRFc6y6FSQykTahn8bJn5VNukHOZYZJ0WdaQ9wcNJUb+KKG5Pamk7I1/S5qqMe/1nhN7
nTYVozxkrex09moptypf8lsAzN5LpohvXQLe4uaetZuKSGs/vreyGZkcHWfejEZ+w8vUfmPCGJ4m
b6DP7KcIe6jUhDgngVxHiKeQ31urE7sO6tUMuMQ1k35qtHL6ngjTP4Fh4I2okJezzplvkQIuC3DJ
NNnQY9U+HSgl3SXROj0bfGzICsGLOyo0moWYPdzAe8SlciF7BZ87pk22FDpfnVp9Ila7csn1kPtj
1dqVD+aw1vNv84jgWU1ZMA65zUIoQLpbYuBlpigw73E8mvBgFLjqQ48C8e3eklBzD/jKbqTVTcFp
d7VJWvA5PtbndePRHaXUbazpDN5kxw+LZXU82/MuQpMKLM6jfvAaNWFNwGNQFBTcWMFmkLuthqPa
RIBcX5NV+oslqbzQLK+v6IhEMAzvO/8pihymk93/pBPyMd0bC3rlnaUeZeokMaClkIQu6Q1KZXFn
SCsNxjLtS7pCP2mHRQr0v4nJhEMHWNL/J83a44GvsCcz4o5bkdrSBMvHaKyz1LbJqEgHvsUu33yA
rUbskMJK8342ZU0q0ni+9JwVSk+2/1d4G8DZbW2k0zappDeMsow2+V1Gv/J4WUvlmU1fKJZZzVHB
X4tXjnBfPKRIpOOrGSyurO7GuoC4cq/aiO8WKmwH1rfELYpmLpTQOBFbZ6nWLRtiQqeqH4ygKs81
rsMoIoZGqXc79E8g8Y8kbSPNfLj1ls56NpyvAwZCrCtxL+zNB3AKbkrbJX1qiLNppUtoSgJ4xHte
cmV06G1VxZAs71yIuuBOcCWlafw4fhZ345bbjsBYgaDYMIxaHu1jvjT3PuVbhpmbTTL8U99GmzBa
y+pLEw2NZ6da9VkM3ZmMXwllMIedui18XlbuZ20QKqEtXIA6hdBkQexLEO/lnsDVknCrBfkA3cEF
NfuSt6OKdEzpEqPBIW7y7j2XJfI5s7kiJhirobOzNO69jg3EpD1dQjPwMrFRcf76VWosZW22VdtC
TXkgulfjkxxjKV/3+770/6amcmz3b3q+NKVrjoXmo3sWQclJXC97m/czS/QVeMyVPxUUZviwj9/Z
VOEd7szvc9McFo1yzIr6IrbgHnKh83xmL9L4K2dMQTg5CkeFCt0qeJ74ASN6XE7S3z8LNpnrxUvG
o6KqqPLd8YoF3HaXIOVdyUa8RiA3T/w9n3kGjDVxLozSMnLYawrn5O+XZXtbbzwNO71JVhN5hS9B
Xqlshw4aN4tCLA0NtOlgYXFGhGV6U/RqpWWlkxJOzZ6SidmGq3VJSvuctqIVkqOTLoBGmA45PAF1
QkPIqulaisKaKHjfWfh9Jf/NA7a+5boEJBWPycILuOBjFUM1IDiU6H6DKUznk0LcOvyPfrZL858a
6XrnhEKwrCCQRKRrsc3dbDtg648p6vcl6cNzhMpgXXkeffym8wE0AuM6QB8/7SsjYWKm58KqG/8u
xdJfyEJWLA0YaM1/lvtES5a03GwkahjZHlnepDuLp6efvDEJWXv7mGSvA/bSusmjwBel43KwDe7B
YPikd8yaunIfOpQv0RgtVGUUgiE0sVxcRNvpM9bn4ZUvBuO0fFCn/WaplMLDlbnlSA47rSJrlZzt
ZYiQ3bjLeQre2/NZUJnLBKeapHAwOMQTRWt5uwXe7VW+A+WP6gnqBQrt/DJMjAfJVKr8GlxubVS5
9hNFW+FyzaKT2d8Cdyog/84WUUNP1HLdpuBUN0Wy/u4JsblyqauhKsigC2c02pqDKYpcS83/cxDm
jdi+TY0wiLPeLZB1f6hF8CsGYalM488FlZNKDf3wNoCdMLtsnzKeC6Xd7PkqKsosMJcFh+U1m9My
/crRwUa6oUExIzLUjfK2B8sf81UoEVUk8JFfkw6NPe7zETSqFzuFf/LqNPCmavm2+LTEmH/B5eOM
VPH3+p10VDgo4V49dpP39JgWh0e+gx/7F4v8cz+5tYHOn591qpYdvsA+oosCimQAvujmsuNQJEGb
+EE2Ol1W1rRW9iW80rdXNW6PZg+mir4T1/YleC+wQwkPqkJ5zgD6fKioFk5ZJOB3NAVtjZRMT5c7
yGw5JCgIOJzMeB660w0fekPxTOQ6PuESrjAJWPJJsaJMvkbVeR1EJaNRKRfOdemE+dffrW35r/9V
y0eXkprILSaRcoFRqANe5C2eRwD5qhwnYy/uTI4NlrycxANDIwGJ/q+21kUbdkxGfhYkgumQ4XN4
vkysuQLNSYfzojh3hl+LIXnOMXEgNLLgpm0T0aQC85D4Plbz1HRQui8lz6d/vSen6IjPZXWWrZuj
/oMVmCM5wdzOvyevqh0gF2vJrbR0rmnbASxbTvXTJwYqFBbcS3dq9TPbpMfbDdgNdGas3MYH8PPS
f5lkFSq0oTc1wR/5F/WcXONVd39E+zHR6JR3unrPS0MYs4V8yAia5fdz6MDQlFZ1HqDs1TJxa0Wu
aoILdC7WBWfnCFo+qnDjvhAhP/pshiJnK/ONM0EHeuznDGZZ5yBx4Rq12ICnkHyDG95ZBf+arqO5
zrWPwZ4YSUPIVOY2dLtTn6jYi11uYqhFGkSaVFO4AwHnIT+skb+mbJmhwjd9RbzVgfkTEgoJE7yu
6sSKl45jbsfdRcOSdFi0YfDCbMN2o5Eo3pa0CzxHEVMbOKvcV3rNcuECAA+Bw5U343kYuplGLfqz
elGqXXROR2/DruBmTAoAbrR5YsJ1kqGsdI+AJWxj5F4IB3VUmK0dNuuRoBI4kMuNTg0pA3bsDOJe
VhAeO6KRvgsyVenDK2G/6JJSEzUGoWtiGVmIo8FZZV1EqR7MxZYipp56NahBKcAWN4Zc71/BmW1F
RBMaqUEwc5RNQ+6uQ2WWXGattVwONb9G/fnvgEJ0KqE/afPb9h07dFMDf6e6b1m/RymZjpMWCe6r
rAxwtqHzAideyW2HPGGvXDAvoc6hXgvZtYaIiUaloidOS9ZNKEtJ+ptPgCpLHeMN8oU6CX81wVOQ
udmqDP2r3ZXGl6m2+bB1GtVCw3nDV2z+X08HYNrvVIH5Rt8Liw2Rnp6KyJw7ev4tCtL+f+zBnude
JQorSxPy6b3a/9KVUHJ3f/SKgy6dDh3CuuQGVWyV5JJ+yCKXxql4lCgvY8YnvYsWnsYk59pmhQL8
e2VUTbG66KDY0g45j51xdcYL7WHZe4pqHeRcLZS8xs8VlIiCbTtKoK1zG77x2KnGd5jr06IWW7nF
IJKAY4fFdtoNJmuWr1diAp37YrmTRJks/6ojjsZFHur/2sVIUtVa781Jix9c/wxj4QnIsuLYSlOz
VcXCrbJYDIglKaZ9z2oqpRIRYD8e2MOPg2KieFaYFVq1fAnrZtchLapjuEjDC6tSO8G2Vo3Xy0bz
k7fpuH/b9WBSg+SxrDWabQ8JoT85Y1VRAT4+tCRSumeB0SjtKMOZvxoyGSikGqtnvgdPiNsetPhE
k/KCVqeMM9e7wqZby6nfKZ2F2qiKoWILXzPVry5QNZ2WbRGAdvBp2EHYVNZvofi3C95fXAMdgJrM
+hiwVwKDKqRPGlkkg2JLvr0GVt5m5hQ33y6C5Oct+Bk85V1pytQGO79R2EIFl3cB+P91e2HvG49l
j17PG3WkPWg3bPUs4jtNtCquyOBO70+5qsc9LFN9ygOt4Ml3SCchqfdHfSjGR2ybRIRS2IeCiMA1
fm6oLpE7KA+eCsk+CZJ2SUChVYMgUqVt8LSZl9SafXOiAq8HNxyudoOWBXu0lGvk4nLX0oTgQD0H
HkaUZpFxxmVBriYX01pv04o8nsL+jJU/TdSo2aS87+3kkXJpNyHw0CqcRY7MWbIO6D6Qtfl78Kp4
YAu1ZPoQzAKYDhn6eQmleEHIUAQqHSVyGYGeUusAqs0Lcj7bmSnC5ctenDKMR+FA18H++usYX83c
V2siLs9WX1CnNldVzQWuQl9kjm4X+KpgOXEgq6oGPW3JjQQcd8rDGMPESDgzdAT4K4J48mF4SVFW
DRhGoDu2XbEGEg5iMmDCD6Tl8nBCMdxCe9vmYIMLrVhuebrCAIxI14UAEskhtHCsDeiDjEFGlKRp
mbPeVVrO4BypyRp0PE0ga6mUHbm6JT/WXfjXXeItpQ5q5G7KlWMJFJsLfIppJyx1c4fvPCJaoOO5
PdcLmPLrTUt9DtWMpcsGsakrGF/znou1xhyYu7UYDVkvy+8W6wi6ztEToSCb0YLULoE2bNG6ZM5J
1htvgcnWVWRQQJLxwbXNYFchS1qEh9FWskFfGLt+T5OnC35QYTPqG28ALkmhGPofe8m5+paUWTea
NfdmdgDQBehbubOFSDGgnUyubLgQ2V8qkkGD8A4bM/jonjbYoihBk11IodLjoYM6D4XyL7+FNZnP
mpVh58DkuCdsuQve7RTkzw56tmlEyk2KArMaMexnXH3FoXQT12r9Cf87t0XjEMAIdUhYfUwFBitV
GIjxhETLXnAflBobbZ52fBP+rb30Xmj+w6EdOOLv0EHWa0ZgoSRFl90uqKqDkk+A7wmpfwH9IEeo
3N810TxiHrR1YJfZgJBXTT7I0oGiE1ANIGQfAYlaBjrSEbvuOkIwP0t/wtySoQ5IpCyqaBM8A2Pw
0fHNhODHL1vlm+wL16flkPSkHRoiM8TjYqmKbRr3bCxaV9aijmftP75D8spAOLABxhHlg0HCld2O
yjTfmvXaAcijfiaR+aycVZEe6CFwUwKVndJvsebZibb8x8Vl11iWvwN2faLhhl6uW0oODwCCWc0D
xsImtUnlRnaTvbN056xnMSSf8f2XZ9yg2I4WTZ9ZqDeqzqbf8RTSBQ0LWSfOo0GPL4vWsZ4Hjlp4
4uTAVfDlpdphKY634SO2pwIW6GjGIujbKHlf6R2C4BizPESUIYNm2dBSNr2hX3OZQ2+ufSxNVAj6
bBOaWAXAe76G3SghYaXZd4tQo93HCpqEzm3uOu2naCa0Zyc6DoUvp2cub4S9AjuJHhumbm4WKhlC
7Jg+XwKNRyKV/N9IXvZwXBg6D0HTQgcVKa4B7iRpP1u17weKXU3nfLCzSHs96HszhYbehbv79Zte
Ten0yQgwkNiUeyU91PTCPMKx0HYyL2Z0c7icvZKCF5yTHLRVzJSG4zNOd8UULf8tVAUtvx2fJsIp
h8yZbsPIRWH/bv+b027YZKXKmMSEqj59rPWuFyM0JvRvVZFVD/hvEMDhTXyU6Zss3X5gjldh0ZbK
sAYJo+YzuiRrPXYiqau4Rwu2FPlQtZwR7zkcYCeXedZm875nES0Cen/AY+fLSEeXZqZVTavl32X6
C4zHoFHhM3qHrkGo2BfOzz49hTFGK7IA+9nlZW01fiWDRTYaXYihUoaRasswDnZN3OjltAgAcGxU
6fYUAAL4cX0RvrVY/yJVUID3ZJaMfmP+HdKxQrmEBcZKSgpg/dF2BvQhVAWWLE/03w5Ni7l2S2tX
G5nOByUi6hjo0VxDFsPkgWxeAWNsJ7ndbG2A86sO0nS2OErh+fgVSYrspb465Zy/B798buHNs60w
8lz3YCTmX+Xp4Y3qk2Z9riUCjp83/bRHnCDAGpoFUCyqb5eK8JdtiwKt8WEKAabpijNoh5xK/h6n
/97Y5VuVvhJAGqZIo/T3fPqZQJV1F+LXGCRm3y/+AdbJzmqj8FOMrtGb8CrP0KXH9kcO0qwSrGTv
PzQ5+efwDId9uxBZv0UJ/L4prZ5iuxIivceVfg2bTafSIIUnB/MaKYJDPKSUnfx1eYVv/WxxTSuO
96X1ydViSkusWpj1HvEJEBCoouAoZd/GDppCl9t2CVDIlzA+CjcPG37OpMZqROCFRnLR9qFonmqA
hYlvEj7WikMAyPzwvgAvYffaNfWpknoOKgLnRqlyUHxutZGPf7ez2wuo1wCjq2AEtqq6aXNM02Sw
wsXZkFciN0LVj6SdviW8gmdKvbeBbQ7GyLhO9NErh3pXMzDrMIGmmtsNM6fNhqoWGX5gnB3l8CV8
hPO2ZsHjvg+QdQUJlxvTCJa+fBAcP3g81SJhZ4QkJvugOnZe6oP87fLii5T7Lw9S0bYDofuWLlQs
UTM8ms9vKYFXx3WNroA1mFto2/FdVBbuG0tO86PKGsYh1lEiumhLHWxoLrvcadzNV4Yo0LBFDxQ6
gx7zAtvs+eGhZgWheKLJjSsBOjfRiG0vCwMPK6wo2wiMcdLNRTZBtPh7jTPCPUNGjCKld1m1vZci
x5xvB3zrktw6rPv4OdncQLsqBN6HJy6mxur8jbrZ/l8q9hqL6hJI24m7Dm7XkAHL+l01rONaQtA9
UOV0YJO4oEaRUKVn8MAiPEkY3isofPHDyPuWfAs8FUDXQ6eZlyG9whQiGQrLQGxJdLDcrdoBQE8e
ZtHW4Rq7usE80x2d2krMskuYflOQtamKj28tEez+hl++pCQZL/tv1hFVhKb8M7e6FodvFWsBNzOs
sFoKdtcVo8Tss6RitmK4Aq77QujcX2Tqvc49NLwfZQw8t+GQ0WbpwwMr8aKE2PaVVHHDrM/ZlsmG
ewnNZknbTavbfTeaLrQKWSRlJWZJFicCJPJncqB0fBx4BQvLWrETuCimMpHwPedFGusHjPgSVr1h
3J6WVOkCMbwNtGT4f/jeXwj4Mt0Y+xXH4EVcPjZ2Td2p7oF0PMpF3Mw4ouPitI/K1QV9t/J7vhh/
rUs849HnhwrBe8NN7k/dZT/OVIW2Gebs6W2+1vAjo32i7XZ4xHzeMy6ej7G0Goca7npDkE0q4psl
DDI3UYgdycBg5xZpa5t55kgKdLrHfMeeiyYEfM2JWESY6Z3eZk3ZEBmByl/kuc39csRAVYxWG02v
YNeb9+ftbjczQdusvnZtY3A0AxTpvws5NWlopsRNl0HbrKpKkbcjQ4l6nFTxv+olzJ6kCt8UrFlE
3wfyewjwUXsQDYG7gfZv/D/z8HGofK3nC7BodzrndQWl3yYvKbfOdLsxn9NeS7OetWjjvSqvhlIF
VRaImJUnWjKt5gIsf94SyWSpJwCGWOncAZvctDIHudn6zGJdm6YU4+ZH5xc2B3aTaQ2LY7uzNNMJ
0tuSnaIqcmaI8Zalp6FIRK10u7cwiEYxSnHU7gclnFvrwnErQvuc4iHouShkhHC7ks4jSP17E4DJ
XCr5JmuoRWzFYzqVhrvE5a5K81zM4M+HClU5friKH3LzyeeZ7S/0dU8FTja+KstARj2bqMGUgHp+
/jjD4oQYK5qZgAUIB0dzwiTcXbDG7Bb0SdmnfjbJXFnpgXLBUfhR6k9jNNJgx9pcbrLX6cCzJuqG
b5TtNVtSTQKty90b5BNpkF/xRHNMYZTfwlAG2hMTLlR9JVc0QwSg0q5AXs4OGHDw7dEvifbUB0tB
cQY1hAywpofS7wzM94JzQF/1fLZYgc/KRtJf0YhFSDMwo5L3S6BWh0dgwfaGAAs7lvRcgRJ828jS
gCVBdtFc8oMwRurWqvLqI1bm1wYM9jrFXEEdl1rJsJqL75I3d2TOUOtYLmENKW3+CRzPkuPNd0fG
q2jksZH9wdRw0f+fKdvjzTvH9yA/Rolx7COp0jZwx9o7r0EIS3kkchnTYS5F90EsumRfOrh/CI0H
VJuEKpo2Pih4Kk8Zcx63KiFAv+prsaW6UFeYkhbaYsVOdY+2FpG6fGGnWpab1nRlVWYf3ZdilXwh
GXnJtHnzS6Pa5G/v0hHcweDjgwjODwf5Ja+FAwqx5LqMYQUufJ8lsBorgYZB+nRhwGjf02ZDWjaG
DCV02jUPevcg/j1l5hWsVYQ/1pP+V/fHeFiZSJVuyVFeEDfKVrBcJjH2UYfwqaRdin5+FtvkWGbl
ik5T0HnufXvoG2MfO5DjWj+YfvHN4KIMhMl5sp0gzbFwzKy4Rxn0/2ScstEK9h6rzkVUnUvy1BcZ
oOkfzlyBYeLlKQPYIiLHy6d1kSWw/E3AVrVmCyatlvi/y8931jDlbm9/Co/1TBPKbItiM+HcoKCR
bU9FEBUoREwLotKZUbKFPCRih726zoh723WuiBkphWk16NQ+Jnp22mIE/DshD8eW/z+mBK7Qhn4p
0HuhD4qtjS/Au4jdpXhnGARidf5rBgU56XWwxnJCLfBqD2rlQx3JgCpZ9UhExs8+Dc/ORUovDwv8
RucQmWDCrqHyly+Xj/hXmRSkj4NZ/yITnYkC105iqTYDNJuGQc/xj0H3AOGU8/N5yYvWVhF9aiF8
BfZNGjlzVL6Fz4IqWxoveynw6zEwUEjAVYKa1Tgs11c9Y1GkrRXhRzpw0xNGxyj+MX6i6JVzbiEN
kSftqiqJopVnOhHZQTL6O/+I2HIILldo2XswDlXQqn24YcNhCnre59Vp6S64kvnUMnbNsdoxN7cQ
tl6uoxVZMRiX0XzWUZczrmTwOF6aZB4/sK/teMbIa92eEhFjTS5Sj3Hq+ZvQmZhPNd0MXCNAPPfo
DKcTWgN0/9lvo0FBPFUb3iC1tKKCib/AOPKQ7FmeLSNceDSUx4uUHRhfCGHX1B1z9/P3BQO90NFU
Emhyrx7KBMnhqWd/megCw33hEF3lNG7xN2nQ5j/y6SOKwvKyDMy4he2A64IhHWwYC2rrkIL57E8M
aJpzQdIACqDr77quLdE+gsC0nK1fLcgHwmiLYK8qV8EplKkOPqYhbiANV/yMYoIxiBpfLuqOXDRc
dsq/opFbgw2wYxy00mz7zQIrF4eidfFUstUpCnh2ooG84li/gldTZ26PGECv2hBaq1aHBsK8Lz3j
keuBeQ5C1tR/bUEBm2UJVBL4MzZZaSVF7/Zf5jZ4z+T2hh3zVwyzWknIjh7t3ALrehXuh+dsEo4p
6od5xFbBJlEiWNV/vATUoilpZRThF14FS90A+uocrJthT+1fqaxMOcru1z0jZBFmEGKsybEwJeVr
BeWkMe/Du2WAal1poGh121tlGMX6HHxIqo7RBDUOjYF8kppgun5+heOEQ1pBWEF7a/+sEVAMIJWA
tOH7ajM+ULmTEXraDE36YuRMaPhPF9HceDkIFQjUkyaUBzZQj83F1x8NTEWucfhBYDNmpRX5gRJ3
WrllpKOaxP5KcEa7uD7k8PK4u/IonYOnEHBG02ur9Doul6BnyufgCvcTMuDeYf/+8w6lgkCSjCa6
oeu40N6Mv0uvdWe6TGDqQCpzuRlQmYU56jmXO5CrGOTtHjii4ioP4Ic6vdXNd7lZ5AUAZDRynH9B
FK/phN5KLJpeoBjR37CsqvBAFEprr23qmD+UEDI4PT7a3nZNP7VvD9h/nLTiseBL/uvPKwm7zgM6
xfLaLrw+cfsy0jiRU2J1g7+FvZ+N5juslcX1ID3lwZorbVxuQ9Jg9xas/CGGTXN+21oRk/z6nLxt
uWd7ACa2H4Dr30ktNJS78xz/wrXR1Svdt0dGmfPHjtWtTw2eHB35IKPxa4KRVBmYPggQlGCt8XaL
/nnC4a9gFyqylNqNn/LFJ2O+LQvQZWn+ut3+DkFMLsht5DILlZ+hXiiCQVH6VKdGZeFbihbpnA9H
tz+6GxY+3CbEMFQpD/JRRKyoOxad6q99NwdMIFKUvMRXlkuC6D6dWsy0mdZy39IVUZY4ZmoMpswN
HoqQC8n6iOZ0aC7OYqC/+a2Ru/rJ+o+rgqFOH29HrOAur+EzfpE6JTFUYOJdSHZrhFGPqHtHIVnE
RRxM5j/XRKcQHtaPwerLAv2GbwLKOqrwYl9bcezOyXrTfKgP4Z8DC1rH4eFf4RAss4U4sX+HlcpD
0jIsHxDXV0Dw1G/oeNxAlx91xp5OMAg5t0q5Qs6wJ6mSX/76rXDYhWnxOAeWUVRqAJosBmB++E9K
3mbTwdgBi4vy2aL92hgW9K5bkNiivtDSh0dmTdHGpJ/Ht32Fz8Wm19B0wHuJ0d3+Uv6abR5UtFCl
aqelCKfrLa3B946/axZHVA1nyHdRLqn0jyTYt6yy16w200+h5TdY3Fqol83lSFejIrHeTgl5EAhj
9cOM8aGEHIKWV8hg92nHRt7xA5q41B7sSHbUJSdoBi5B3gMlhd99cSJVaxpuSrN09FCdzbj+mRBg
AaBd48SzkwWZFHVrWZxy8/Oogf/5VAE5WihppL86U+m0nfrqgdTKONkAfUOQTR7GrZ6O3aFDKBaL
mmA0Gm+b0Hn8MG9PjIHNbolyqTdKYIy4YkdebtunmytgFsvG8Hk8ZYMZZkzPoa8EwX2YooDnD+M2
UcqY37GSmqVGZP4VALkWy0AkBmd4gD5QcYk8DRn9YA0RtRYEmX3polscXUuOtnJOOUtrxWwWwdGc
FRpsmWzVda5vK0wSpGFZ78Hwti9A2gmvYZxvlHB2cgal8Rv2M8d2VUFj8ckOHnSFtrR9CYAE8tXP
CaoiO8qzGKPbNQjuGh48Tp5BRiGHuKNwE+4Ucxl15Ca5wpX4HetIfQevAqlw/+Vape5UIq3UdFu1
uY5MM+/MJCS6T285Uq7iU8N9IEU5SdJEdcJ0LYJM2z0JUtkWZOdNl/PljvRwM3A2RGfa+2t4rEhs
SSzuiw/f18U+LhBgRhINAjcSIfxwE73omunJMnQIlzpjejm8gi/EWPC+L8BZjIYwtLN8JdHmfkfv
kO+zFDKsDEMVAztgzdJRXtl169Q1vpTj0dSU5cq/tUMOCpBa1/FAQFvX83I63AM4rFUVcLfWM5j0
dlOn2Oizi6OC+68jkc5RgVe638gOefkN0qan+t0rWvXWFZxZNIoVRsd5dGNJodXOWVCDp6Kl6Q6l
sTAIxQMJ/hSbEzh8+7MFFU5CQ2VWFKVZOwPtsYsVzFgi7C8Y5PTtNADY8/tvkBhIY517OhpXKu53
1TlLqXE5yeZKmdOd8ITXH2jS7HEaIGtEagtMF0tllIFeb3EbxIo2fBSlchs5qw1XLeLiZsHeYW30
KXL6DUv94+XG751tmzWj848rzkOAkfhW6vLjXfx/p+YkePX58XIGpmBHO+Hoxst0deu3PzbAEH6M
G2QWCHMBT64/BjAGjVB1VH7x3ffEQ4ayYfQDli/ekZors3crUuFPYm0BVbPoQkyb3iiJeWWMQbcU
rr88JS3j/hKJY3UDCkZU4i2BoEDfbTt98IqL9J59PqrXZXdx3PKB8Dc49l8oQbKsjYOd8pBcHqUD
5z3mrpN8YTDyAImU8lLI934nAsckZLs+uXqchlm5GTXBaHFOmICjjR0yvu5syd2E0yxU4nN969kE
BTui2BMpq6ielIuTmqLBt5uesm/cLtvkBXq1KSVqgmQv0v2Bem1KAOzIA+BXNlcoCPqDks3/zLUr
u/amOfuoo5glu7aGHrKQ+faMWCanDqharooXGIg9gu7lZVbLLXuUJTkSeEykrpOaprBD5TqpUbym
Ds92Gt3B+7eCU15i93m88fuFVcKq4sFD1duEqLKeHjFQw69yNVtH+TR07krjeQWQkUSxTG0a+pkQ
68BGFgwF29RLo9SaEbUSaHB2n70suyHVEOQL7K1UOfxeEvb5eLN7NPgZiK+Qa0l57jnBRPuztBxL
dFAtlkv3AHYYQaXurDOWcuzTx1E6HSpxhzNtPxUpciBParmUw/EzQ26d5DEkC5ZLMJsijQ1me53C
1O0qonQv1jM6tbddsNMqzzc4eZtKPsEUSGgRmnZu6rOxOn2t0h7XBaia1/Zbix7gu26AfjZk0d3p
XJJm06tHCTvZ3vv5YS/9BKiT9a8sUH4yhsLaatZjQBBzRCIPGKizEgGmGR7Lo3K2t3c7TNRx0vBR
OvJIxE72SN3mFZY6/ibz2jggYCzPBTm5EjxEHpSqPdydJsTdW+NC5iqjlutTxJA5HwUaSwHPOVQo
/Gqv7QiCuCoW+WllgKjT8aOSk7uwF4lYAnPg0wch1nU3AyB5B39kgKIUjrR7sVGM/T6ysqbLpdw0
PMHwFzpgqOd2pRdaF2nMp32hsDqKD84LK9s4iakBOTrCQvL+HkYTBRf2YyAjzq6BczS0AbCnCAjq
eg6v4OnT6+NBkpuo3yeOiC7XWhTXFbj5xPSHSOWEMpGJzA+wpaU0TEM7cum9ZIxH78znQ2I0zFpB
ITQoOGtE7CpwbAQ1EweIXf5vz8heqenQpssIBgzkC013e6w7AfMM5BsMdbHJw2Q3eWaqMzN180wU
uCjr/5lSrKPohlQ2NHv4DKq7UsEjc+NVzos2uvvu3jZVTZFQtZbCJM1M/mK3qbxs0z2YRwtR0K9a
87MXNDv1Cz7YbicOyDp06mu7/qE/rs2OORTKKeYFxOk6OS6uLsYRjlYWUnPGy56pCfUtSztws/7I
O76+bs25HwCZ2cqOomWAKk09JVrL6pxGVWoxDTMGgyDsZt8yebg9nWbUyD8buutTIlbOEebM4OgS
7+MHV4FKYz6zBtaZIWi2gFr3qhhlRYsbpvelgmIYFVnNLe1oZibkExHf+WJgZz3t9ZliJEcKuZZS
NDrl4EjZVy36HgpQMOXMY74sLFAA9VfzeW1j582Qr/HXpX9dB1Dg5Z+9GVsL/GUvAxU8EyC1+AX3
Rl0QL/V/lKKYgxqWfAHAkJxRYDF5mQ8hbOGIXL7XFrSouJVe1WfM0ki6XCmEeU4H44F1UEjI9FsW
bBSHzCvU1vRFhwbsfv9/zN1fpZoLvfT2sqTyjLWIYjQwXYCvcoVDiVs5dR2Xooega0RjZbd/ub9K
s5X4/00dcF4OgFEtn28tptje9zdMtwH+a4P4aZJs5nGyCvLfldrAefVryUjkKsRvoMsNI7uzMjyG
uaVdheJJpjN5stCvJIrqTgmYxog3HFEVGZqv4zQuxZqh5VoS7I88+cmC5T1ooDUVZk/EP53jysuy
zFHWdz3FycOfhG1czy34ZoMRw9USTzDBHEtIF0KpWchkKmH1I4A4HmbjftjUiMcaqw6UvzQz+XLd
S1IIBbLIyNpItzF+4p2SyKapaly8KpY9qA3AAOwudV0MFuSTCihT0iv8fFSkh8EFoe958W2YOWaZ
xe35zjxMDBEVIFWJ+9OyRRbaytrUAvuJTuIsf8shOLuU5RDOle63Vd5UQDvAvL7euU+S6qGGjREI
HiaayUcJ6tqDw7uXhAjrwsHZw9toGrsazr0gnQmERCAk5Jh9vBzFtfattNCCXtxvNr8ktThSySAY
09uuWQAuR5OdsYUlFr/+xOTaMMJlWGfsoftJ6sYg18TQMnrWc0O7pj4JSUMqKT6zEX3eaqU5s3VQ
nDPkSKxqcCAeXrNiaGDishURM4W5ByANzKAM3RKgmuFJ4LhnNTRjZFBN8EQYEfYCbegWLyu6k/C+
5T4yfgmrt4cktU82JBwWf9Q4NN5YqEiEO7MrUEx36yoYdtQ2MIz390vXga2+T/UiMK18UYdxayYs
THOjc/fDxX8ZMbT9RkwJbr6xUYUyTqVbk9FL+l/bFw2EOvMwN+/mDdkoEfeS19vSm3IXECOCCEJI
68NXZX9gxLCnKrgdTK9VsnLPnFx3cbvETu0xGkNx+LvLxMM36ghtY9wG0B1aPT4rnYdbKkH31Jdx
UwLDYq0S8LPK4/XjCxOo05BtQ4jgWgPWETEXw5H6yj58rzyzDg6ugBdK7MHMx4kmImxOdbCnubjt
tfRiL+8IveyXQcfds3fCXfzc3+inAfIFrI4r0oZYIsFEPj+OsaOJ+icT8wdeLqiepYvyHRU+ZFsf
4l6EewyhGgmnYYs7nqu0KzBBoaGYHE5Gb/96FSFswwwWJnehUJKEedyLCWdQaXk8iY2OTWyDWmF9
Q2T78UCJeOlHyV2I1KFFitxYGWFGBMVYtxBcV/Af7UynuyihfVFOXmIb3VSB+VDDp31bqRzqNEDO
fadi5+8aTPKHClcP7V+1Ssbzjv6w9mPmMhg9DdGRaei+FkwLeHCe/J6Lcwqg0bsG8QVIZ4TRyBwA
5jIU80VsTgVvaHrUnN+lQg+13dynzVqSpnY6FhDtV70c28o9Pq6YsFzorhT9pBmOCVlgmzvzeGef
Yn4T885xc7inujN5bCsm2sgU5lYQtQJ5sflStuN2rTNAj76RWDg2+nKNS8kWXgD+a1KuaeT6LEJI
xx9wxcFuEB4JYDku1xsOTA2yUWpyS5Q9qk5y/ic3jSHJaV6a/Rt/1BWeitAhcbumIpGIA44DrjN1
VHGuZD4J2AKeO7jNwGXUmVLMBtQs323xb09jzFUkow3WChVAYzkNz3EIofK7qh+tnRLXujvWt4U4
Jo5cMWdOja2dqIZrPnalIJPNC/3MWsYES+CQAzqfr0a8PKuEV5vKs1nhuMFiu2qiJnRZkqYL4du+
icmSJ3XZMqcMBY59iJrKg+56XuOhnRxtSl3zL64NtUH8QpPqP6oAJeFVJlBl41XnDmta0hSJgeEY
9hbfJ2n5waOpdZ+I12fqSwbZC+lpRkwbsY3PuIjsZCt6AYmId68rlnsAC3mlFm+FqHD8h6p+d0IS
NqnKVGpHcFlIIz4eTyo2TqEUOHw3oitr1sjsJO+OYUWomrvQwXRJE6oUBmC8p4GfRRQx2MeW0hpt
yN6rFnJiTtjDHlPLxnU4JlFv9famPNgTWosKiwpJSKgski/SBt/oEC9QobuOBTLmBq63zIV79zim
d1BexqmlSMZncB1Axc591ow2ojCYQK+Gd80MmrRoalcVs0tiDcPJ1xw1vPIR/Ot1qdC8S8YTygBf
yG5vPpv1ge6sFCM5opw9QE3tFRsHSa+ch3BbprLe1RHnD/Inhic4+GcF9dxbf6Ak4wAvXlndvSmN
Hgrq8GlKUCnsSzEBiWTRIQoHuTg6MS3/sc5pp6qne3/WOHtGvSev8ESZt0b6DVXLnlvwNnOuFhCP
q1sfqFq5IsbLQXlGnVvdJTiGyBtIcLIl1zZyOtySgTaQ/tlW/sUckHYJjJdA5VuQeTK2YwYxCzGQ
4TPB5IsUPBNcaie5p9iLTWul7g+nvU8hzELPhFMnpP4EMVC9IgC+YWgJge2P0rVEMTu8CCwdl7Es
yFfkLJ7UBBuuqo4ap3g+ncoYkSq3aLsI5I5I7v98aE3LG9oJAuTTQUtBfppXRjBd33IF2BCThaPu
0LX4o/y+/yiQ0S8L7+WDZMTdFqyoqJDbJ+c+UWY2btuVovjyixDEZwIIL86bT+yXFwtx729/2rir
nLcgDfo2FejQ+QaJ3q6m+9YdHk2hqng2eMtWrvdjJi8LPN49UYOTZSlxXMzUvpRM4s6KwoR/ePJN
xPbBooU8HSeelI/HEBZk0ILdPsZ+vTjYSVwU7d9qzBOSfxxrpgrV+W87RyEOGXZImzaEuGVDF+1Z
6XC4EkGtfHeUakBgTNMiqkOmubTrw+YvrVm9FqV/fO00jlrIslhFZFAmfRsl+gHnb4xbLJ3ZK7Ex
YBpt44gNaQVcBWJPli/najMR7SqH1z/Mrh3xol8eTIifrgO5RC6Z9mn+UtjYPupJFeHJQqm+ZEKV
+jMWzn7Qq5oAO13/Ea5svjdA14lhKYUbtL33EF5ISrzl8ESfmMwa09jiSszyWcpJgtU/XUed27PN
XlEtivoOWjiG0xR6c3AwuL7bw0Is9yOiXcgkKxlbfA2BsCs8COxbTXTtfBJQjUwKMBflrGRiX/Wu
iGlnapETHZniAah8+sHX984QumZAeszEQ5w3z+WuPFqOxXyhtfvd4+rDIqB4KttJgVWy7jeRBVMc
z9sc7oui3bpujpEuhTY3dY82bjeKeP2jh32B7ZI89navlugXEC9CPgoDEleb6jpPygLUX19F9gAz
AhPugM9m2NvBL1oQr0itqfleqwgWEYBXfN/iyR3dKWbR0Ovyo/ydNheGX5Xye+ie3HXlntRy41aj
EojM2qH26Ciwew39asDD3fT+Ly1HghrgrVx8wIqU4eJxnchGExawWQr8hRLG6wJXTYZ8Y6lB7qFR
f3kNAr6Rd5n/UsCbB4GDHTYrVaCgtEM5M/QpYE0yJ5idhvHwd+ySVQQ8TdfdHgEm69bCI66+HolB
XuQecKRQE9qBV+LcsOaKB41j4GwDA+NzHq4OChhFStGy2b+EKbcd4oNocNDpM/DCFafv9ISIlcHv
L4h5/GkgQWYSGMfPwBe3esI6IS490isa6a4eqTYuwPvYoEF6sdWEAHsdbh5d/oafEeg7KiFCqplU
AMUwh/pxTiO/YYSLO3upV4fIYcX81GJWG69EP+TeT0RL9Q1WwKenxcXDpeq6ng/fUPEYnQ9lRw1v
sC0ds4xWidCoqhyGBWtPWXkVMj5XaJZXU0xQQ5vv76qeX1ZKsN+lADXXfnPuirgEl0H3mTi57oLJ
ceLH9IY5fX+ZrkUyRKQf8N9T2XPH7QangbBIP68H8wMTJsgZYKj4Xx+0jPkDcQYVs/0MsrluabX8
spAG17pd7/zneHGWk/oB8CRgvdvYPCZU+XVFetHGl9s2/DskqEhXy+N9OLx5rvgM3Crq8I6Al5vW
v1bsmlog1wJRZQ3nONF+n0B9K0PD4+x4MFiHbdLX5k2NpIpuAo42nEBjeTgzI4J5Kk5bNQdMRy2H
sZGYwMG8mRMNKcF37WXzoADAwy2aak9wNxLTV4ACz1RXXKdsf73VH1YvGTt3XOTXltVRd5Wt/7Kg
9Za+2pkdGBTeC3vkArooAheMNgAzHipJhi6Ocuuh+9Pi96U9rx15DLlqGdY0XZHLsfiXIFH0X2gn
mTm5Evya5e6IUEL9QTU3ZvH6bxmzfvNzo+xFpI/rFGZSFitWxi5BJkCcUYd0NMnHUfT8z+2bRU0Y
MVZaOG8P33QlqjQ995uu6RX2AaN+DM5b3aSyWFbSl4brwkQ3ACQnBn1dU2MVOCiTuAAmzayhaOwP
4d7/sUw15cRMuYAlA/MUL+vwPsirx+lCsLa8XGW7KvpY1GCmnGCC7c58cEkIoppORXmodxitfYGB
dp304tvYawfnVhmoLAYa4j7z6RaMoupuznQeS+OGmtmRpmC9r1SQ3LW6G/me/taOi25NiLo7xPR5
vGyf8oevf22+wIhoh434WF+ESgY1NUST+DlJ8Zl6Pwz8MVXd9jQjGKYeT2vq82PmK92HhbgG+WkG
aiK/wrX1T8BqM+s5qYK2sxTK9sVw2tJWfezTc1gOQ2QYQ/B6JcGcJWCzKRDOEivFAX1lFL1z76hZ
M4wdjdEssx6xVGVgubcc4b3py6BJXp1lHXZsBM8tQR8R/RK3Kx8S0P2zty/f3n1ckcF86uPZahRy
7dch6R0CfLTbuUZpywynIbhbUD0ZyuUW7aMTHLKPPaSqJy4IR5Om26sTx59SOBtn+2ZPf97VcIms
6J2FV8gdJxt5i9ud7uTDz0Hj5HYJdqyKE8jE47zXSh7cvhpQt4p6A8LIP4yrgGreZ8w7MM6fQ5SV
eC4I48oIgGCGYCKMYVmZPEygdcwxzzZQSEdZaJ0ywdqoncyL2y/TIctX3Wjc3oYjfHb3PlkY08KX
eIu9NhTI8cRWnp4DmefrSpjWnTvY3nolNge9OHICgbZZd5FOqDFGE7yRk7EqXw3BdI8eHpY5EJXp
W7L8Gqck2TbNbbzQ3Pq3nFMgUskSdNHCXz2+WAvKzRH4IqgAsKxCUKIIP+x67VnrzmerseM3B/O1
sTThzoa80w1KabO7aKY5MNglIaXdCcvJtXNA2ohM+NBzKR0nO+dZaTsnAWsIKGfuIM4EIpkmt+9O
BWprtw1jCX/mGDNiSn03GYAdUjwlzI9qNxmZDrpXfhvyhQ96lvLyZsPVqjSDyeBCk94W29h/6s+y
8fCG/tLaUWRkyc7HLjNJx4N4ivFPKNN4ltB4YnAqNX60VFLMWZbPcb+pwxKIt2cRYgZBsyJZIdcs
52/pu06dj5OaPHV6lFNPqHkJSz6dbvg2pJLzreXwwJc7ec5pGrkgy1Zv2jcNDGPqyjrKzD6hkEBm
uT56tGj5CIkTwwZNvT1OHTC/CPbKwVwKwi6WgbwLJxXL6tpGT02yKlH/+2fAj05V8FQCycrrcOSw
7FRAc54EN3Cq0Y6eHH30JihYN3bsoDOWnX5i324x3BBCrIslai0wTvQcsPsSm/Jz9rnN8+LOiDO7
ZhrE4N+HClAl8qJ/YhgCK2tkbkOHne68fSNnu+jLGQxKTIQeGDr/isJvh0mRjUuDP+n/glAkDGMC
r96BECco3H6Y/UvB9YLqYJVayTP8FJ06rz/2cqfBlm3iHqrm/7onII/vNSED727vUiingvyORKsx
204cuYyv6iQ6aBZhDhRAX0BPUIz9QG1HL0ugA08Tvs+DDoQiXfceHZVGc20O4Qcw1FDDD13ZC99E
3EAiVr/1W+Cnbw7fNl+mHPXI7jKyj7wan3GUheuub+c+x1YBtPahDQ61aWC4kk6bZRwxmTzdFZrz
BBtpUw0JVY1Z5eF3bccUvb/Tt+h0wKCMyQ95eHm8D9NrFEknVxh4VXP3rVS6Hi/9soB1WA0bU4lB
3EErea6tWPonKHhIR69RMMxzuuCEEF7isNpVtep40Ev1XeIjMP+h2U/ikN6606oBm5tmFTJx+CH4
6i2hz+KdEMx5yAPAlhieLVT47mcP+/uWdi89Zwy6D3ut+PwrjP6OI72Oi+0ba+NrzLqA8hpwEm9S
HOZi/T7eCKI6syM0RqZZbZvccLN3qAu0IOz7n4tumQ+tDlniC2ImU1BgYWXeDXl1Y7C0HEOEeuHk
lvY2Zv5vSviZ4c+y4RKuliLtgfP1D78P0C/odtUbQsy8v1IOYTqbG/FexytjY57eKZuMVXwB71hj
/7GXxpEE/Euu7+eG0gwraSmViFd958n5CAov8sLRkx+rckKaCb4MIno0AJ/Ke/7bn4gjZ7K/n7Va
IGE8jnsuj8Cg12qyYsqyBOSyfLlnXX+qDD0vW6C76Jk0BR516n/VZe3BahjCtCzbGvaGou7Th4yB
ZQet4sqoSSV5ScA2eHJwxLnbWS9Dko6MFFKR52xi0Z7Q85nw6kOZ7kN5txr6XLdOGtOTLlElvisZ
R8sB9NwBthUoUl2HLsrKXYD2xPXhidiXfpykDx6hymUIdr/JvMn1WOlB7nPKiaU8clSfW3fqbTDc
9yDmIzNWeJXJaMQHtDmRBsWKxqk93/SXcRrY+mMSSdP1wVTPp6hUBiqIbgndrVPZwGiE4SCVQsP+
ow9GdJ3E0MrA1zTQCIe1icSvY+pWUOg6eKw88hleqp8NzgMS5lWMx8gtKvE8dRLubsp+WgadHCCL
g84wXqs38Tcn7g1slt5aD6FkZ7QD7OGPdn+HOuUUi6UnIpVHyEnX2dUSKCDoXoa1qDfcrWrpCvA2
KKKbV81kKgmt+/MZjGRNsCpQKDZVWX0w6dHCzQ7Sp8pBKIp289mHvDF/eWtU/RYOyhAmn3MNFG3d
sZSAsPpC2MlW1KWVmNAdwIz97uBvTwIcuhLu66mkmklT+GQnib9HAYhigov+bJXNCWgs6bvPx7cI
CV7zysh1gDp/QhdIjN0C5Gyvp6aGD0tAvS7te5yUIeXnyM57kzPmOO0ayPlnowvIqlCcsLXgcNP9
4121MF6QQ3D0Qo8nCGD9oXlBJ0JZNwQZhpjsC3bTSGnUQSEg9Pub4ZS3DFDJYGrlEOYfqQkbh/PE
8sOB0nAzpkDrOuiQgk2BovD8JFUABtMM8PfNMFBz6X3JQCZmQMBkcSbU1W8Yf7okBk3l/4BGMpky
3/C/q4+bQF5HzfKc4oIof05JaT537AjeQ/nY+8HovQwi69XAPGFh0R1k1wzWzakreLYWgLuC18WW
k+rH0mHcVHNGQu+mIi0qw12vyfjB6U/L/4FoyTFZp7mVYQZkbg9RDR4cc78BIOCXBNKRU9qN+/5p
q10VzPpkGaxBkQsdnyUIvG9p50dg6CoY28Y4glE9NkWqIjUizJmpewNtTuvh75LmzI6mVIOxWFRE
TzSR6SMNEn9+4hVwhb6tRloFN/uRm9/ktKQIdA83t+TaStIxYR88AnnOi0wf4peEP4z0zBP66/Ts
eF6A16Lt3msR9n0MbksxGhwLvfBlLyP47LHnq5x/D85S/GG3+ahBEF4z1FlUIvT7FK0MY3uQfHUw
pThGML7aZpKYhDjq+N+ORPa1iZ3NRere1YDgyTr7caja6++nZLz9WzjZki72/pJEjnhhinaoOZKJ
xcksLwrr1P8TXIvZiTXaJwY/kbVyQxGPyPbyi+PpfWv2E3bK++jKC6E/Mhm4VRRmUYeCC+YwxDVs
CdZ/Bz97+J6p8/YKVeoSzhfht5HEOTmxZj3S+X4JeAvAoZDOgq1Lj40NLfRwH5lMcQ3hy2yXwgWp
sSTc2EQbklu80uJEMwLi+pMc76byHawY6laqZSCXtpLOzzRVEcJTagJuwmJFHvy55tod3P9u8ggZ
6MYC0UuUtUcJ1ACk+2Pg+O2vx2WntRwmCG9bnk7qslILbPwRnvse0vHJk78nHk8jPS7dT4iCdvOC
jvK53+yNAxqarr/GHjMhREIQKCz5G2GNkFqthbDIFIXlfXLQhQ3KYzM2W0qbXPeukOl5xigA7plD
x5W/i2yalAR2XNjUMrXsDqpyag+vryiyYHoyAGPubI5LDrSoGhe8XFs8etMp8oNS+hUOIORM3MYO
AwOVZki8VV6Xc2Oa7HHDjEMgvzLZ6mSWrXb/ueVSSN1e4RLjEoah77wr6YqcdsIiIWu3oeIdboOO
B4/N8UzG+m+erVBk5LgckDnL7S9G/2SkATmJ8Ufb/I1AVR2A2sB09uW1TIHqNOXkAybUhOIHWyuD
EFtT2aSx9swaopAcj2FijW1sDh2rwcLNZUIpcSq02z5yTgTpk9NjgRwAVxcjmedyuF+3m0vgmKWE
L8f4I3BldPPaPhEl4HprErZ0siC8SNvVqwNgnO0f29SNE5JTsJRlFZt2v9D9Y55W5A/vzrR9WUYm
dN1sxOD9JKAtYi3EMpffvMPXVlF8ddnv53kDrUs+ApzlAz/YmIfBPdvDIMelg+l92j8AvnsPy2Jd
GodCrR2QZPidTispiJ7WruTVNfmTYnuhhr7nRdg7yPLY0SbgDdhxmhUOwChb9ugRvaQsEn1sluUZ
6fMz4ulLIj/UW+ZyhdRrXMulzbB1i96vReNQSs2DIogrLupay4rSxbIUW0j2oUeu1shf/8vAH8a3
5R26Ld51TyKJpYzkrT0DcRTbpQ09FLY4eIzNCGrxH02MPjlLOlo/yuzquZxSO/lwAcpsFXm2vV97
yVtrmdCZwoZEGjz6K54qQL0M09DlQbCbzXi+07RsWSEfnUhqhpsEG5lA1M7rkmD8faB8H7x3RN75
6Aqez6vEl7FzAknxBGzegHg2YYV2x+6sbzcLd5RWOAdpoGepjhtYPdrppWi77dfUjfdoDajC0x6E
Xjn8JeD7JekMxQ4dCHrEi62IsWKrbpbHRRG86YABBa+sQl0Iydg+F1Zm8RPQs9u7BEp1dsO1zGFH
BQL14Y3ZdRKo9r2kBY6q878Nk7w5E1GjJkFzqctqqUWs5uS2rxijtKG3t4h99Ftt/Jswdm4jhYg0
i9ovzYV4UyVYzEw1bnTVZF6Zs0PUg2zPrMgXmDFXVggnOQ7SUeDNkJsx/tcTpL2KyY9greoFLuHj
RRd/2hP8UG7wuhwVmXkvhnSniBgIiyOUJKiXmid44E5MSAFkcJy3MXGLxYNKEuaJWI/P//Irq1u5
5fW4olnMsSidHLn0jW+HQtTEYUgZjIxJE0PQovxFz1SWCvDcqqBUYFtlDq4gF72iRkswRDobQ3in
hSUh5ImCOZaajNnUVsScd5ivQKb9ZU1rjRBWMMiwikTEwd2npV78u260R/+nfwomY7AC5SpgnbXA
+Tft9itbxVPmWJf9V7PJphMH2GIB0usNSwm4m7Qhga0J+N/IvOGOh8uQZLWH+ZIq+yxVVx6SFLR3
EM16+61n5zJ4nGCrHeyE10Owf7Cx91G3iBb80w05Q49/zwvjaaLluYqmOOavZnK63fPkpr6eNbPC
Xqt+gNXZpzLVDepnO+D/TuX8ue31HDsuRr16ghPpIuaTjLGMd0BcDk/A4bbFdzgX97HNe4fFIF3R
ldnP5kWW5wgysxj4+9wWfSQijBiCASmrlqL0JStK6yuSdcIX56KcVIPET0y57iTdhqPp7uuQa+tP
v5DiVn7ZkMDDk2uPTaNcg1Wpg38p/hLSofVcRzRca811yOUJLa9yBPtpqedlC6XQyyuoMgMjjskF
eTWsg/BSLe9Np36cD/OfD4R7UhAtGR21VqRykw6oooEY9+F1ZRBjrn7aIXDvaEA3oHfSjJybKsB1
1CHu8/tx3RS0QNLR3MRHXo8lh6WYi4eRirJ9fSDa2CJx17oNSBlxRGDhipQ/tlT0tApy1kUZ0998
AYYC7O23wIv05Aq9+8MpTQKcC22X1C3/0BEWPrNqDUeD3FEA9vY4Fi2uEFIJkKVB7hmp0qxNtTYR
58jEyC0SDxcelSvvBuqaGxTbyDufq0xGLUitJr/YdHIc62S9IkpwJBzrmbgsXt9bIW7NyBLNMoIz
83rT+Z0f3spI3PmiEvKTs+XG6OkaP+XzwXApQ597oxymyBsszUokmRpgX+P/1HbrfGDUNup2ZfRT
JnEF4ckG4sDYE4B7KsWyno0qxQ4Yn0SHes3vSKr3+s5t/7lXo9mL/sX6nYAJF88DqG17O27mUDSK
k4kQqwSzvoT0AUGDvC8h/6wH8wtzWVvdHzOxDhZPBjZv+czaNXIMXT0gYegAEXeO/WIf1H3oflrb
W2XrHQoREBBSu6/wgsUJNi3eeWf+29dC4/reT1+3tw4rHhvHxVZkLq/C35oFXFgTcsX5QW4ug+un
cZmPS0aU4Q+TI9NqS1ZgPUlGdJBHXcd4h3YWWH6T/Dc3KAYh185rvsWZDl669+zl4u2PyjpDAJaL
gjwr33nxxaRJigZFQpqJYrpl3Mx8cMaE7Qid6eN74GiPO/S6zINJzNZBppqMKsdZuM9p9wZIO2iF
Z7e8f/fQ41+Vr1nRwALuYdgVZPNUR8kiyBdKLWREBmxprdT/e37RYqx9i8fNjwl+CrVlbzOF9vns
3keRfz+niG3oNn58O2KKhM3W36MAVX+L7GmwzCb6ECkk+KGQehRF/o5qWeRkVUTL2PpL5JHbDzUe
ArLXsh6rrhjaXHMHx4FEVaHsjYN+DAZ42K7PXAkgO0lSOr/QTN5IANhdBdU01NpY1BdiyjEqsaZJ
GK1fsKd5BVb4Ml5zyxGq8IQfo6ESUqA2tPmarh36lyaHj49ukuXiAtP9FGhkhRiemZCJ7nhvlrOu
lkqCAIZXwzi7UqkFjojAqSMjE7bWygaP4OuAn+TzbLoDlWWHVphbWE1ZJFC3t+NmNLpYGMUv0O/B
ooF3oIhT2sYj88OJDTfQsuj/7KP5Iw/JKJ5KEUFBDQzTnnaR+o0sn6Zyu3Zm+NKPpkI4ODWhulIl
so+/WXXILgD+/Tk+Z3UaIadbp3vx3LO24nun8iM6WaJSbq3EAxR2UqDtZNfoQ2QAseumTioYDdOk
ozUcgY1G3g3l3iSUQYX3XT5fmhqTDQr+juEKaK7uLVWX0pJ97KBp5ab4Ux7TvilcmpmmLszQDM04
1R796wkZk44dKN5JDu29QB7+C/u8rzwx5+DUVeTXj6z1svB9/utrAESkD1sSuSGm1aUIWr3W45ty
0XECu5PccTWiWCQpMY22+ydaf4FtqCvF7fjOCsflypGNh/TM+Yx2ygCkzZaTPnQywxyaAsgsqSU/
zE7mY+Gfp/ChpWC8kCOBpr4E7QXR8U5tFcAo/dcnxM7xBpRcAjAN6QuTnC1YGLe9dt4vPuFGt5W8
QscMshzaW5b/YU9y5LR4eKNAkWU7HcmiVM/y2Z04VXEKQn3gk0hsnL9fKbCjFfSby3+Pi4djazRn
1E2TKnYarCwDCBGyB6IaaR6eP5hE0RPP0g7vi5Jm9St7CofnV0Hvseg7cwZqvyW4uwh2Wiget4f8
z9l4AiD8L5/Dn1SHzzYzmqQU2rnEb4lUrd46am72SX/s0uCvMmu4lrLNP+PFObMlYfssmFY4ZCPy
34lhwIYj4A60tMGvHRhnCYCDV5lm+S2R1pQuIWqYqPghU4lFhFJ71Z1KBUFmQWxIZOGSNKGs3rEi
7h3xeVz2g31TtOU0UvEBNlR8iZaSLmySD+7OOtyKxKz66YU2P0ZOV3wBpaQVkbpEWMcJXe28NqB8
Gwq3uDyDUJH6/jZk0+fFzCkorZl7NHxNPx61R7X5MZA+vg82TYe2GzrdJHJAjIXHMFfVeGMju7bu
vAgvc9qj1XQRHlj0y2u5HVi8oegHFfP93GQqAtMwAnzzM/S5w1G6dzL4VN8/LnRTPcDyiQOMRV0e
66ysfa/jPaurkDFpv5udX4g059WHgpsN5eU9l1iqbY9rLNNmfZxID0fKOjWAZ37dkHEh0ly0PhwH
AOlh0jDkxCBKTF5v9YTgul1iJnqDUUR+r5a2gIpIFGkc45DmAgaf6errBNwCpchpytrNRfEKTSU+
nd0LIgXOQeQZjRP647g8bDV8qT35IqSMs9BOhSckeSuCRXi9llWD/pmhvblfCpaTGRWsWb3L8Ki5
Ctj/mrG1FQV+fagFApcz788C7k9BnWYe214AByL53Cm5e7R6FHtxr0z6sNyXR29y/lEYgKEbLQNu
LOd+BZskCME3REO3sMNoIDnq78cibVB/39vkOD5RPSUApBiE+ZT3JNtulfBr2SYZnKg3m2nVDcxs
Dfj5tyloyxgTmk3UE+zWEbtbihydwpJKg2OGmZiSDzPOj+yBN5p3kX6FPwshKhKglgZQBy+xHAtx
7NWKM4AuPVAOujttbe3aBYscLsnJRoi9N6HRQlHf+vX0UV3hfKoNW7eXwpGM5dTRz/7himiHhpaz
NzuJ9pmafQ5GMRHFA+PKZDTz9+Bpaky2+xBOkdbhRUBmkUeAdxZAPGJ4Ao/ogmwDc1gJzjhs5DtG
/Um2WRpDXqBB7d1/L4ZnOIHoPi6ENyCvZwVcpk3HEfPtzxso4XM3gLHlOZvjVXoqCzsxYsH1exvV
aWyMmVHPWGVjwZRqF1VyYQRhlBbbYSBCkHpkIUD/sUiNZQr0Ve5muTYmyJzZ1BNikEFfY1EPnDIa
EOvE7pF9bF9IRL4uKEVk0TEU+AQdWq7WJupjMjZwidAuP3teC0LAWFmvVHWjx2IVhnhXhRyEeRyW
kAM6JURNOi3WDjjSox6WMy6pibbSpHq0vqWIB1y0IFxbVraiUnJV+hoC9mfo8YhTZ/kvjWdcvppN
2NgZZRNhJKNljJOj9zzw2sGEYnwRAueJzokeMz9/SzFGzNIsBc1hkxpoU4nptS8pH8wzxdx1xo8s
CuYqz27mdf/h5qIfbgfd4E5tqeZSyyrugaWaV7fZCjfSfxRLrJOKDV+bwK8sWm/sOsQ0V1vn17LM
lNuEyAh4WLcAbg5pzCTQXUfO+DsLJ+sMJ+xSUdDs3h+7TyjTJsMYSKZ/7/YPy5GiPGnDxO1OMP8w
36YXReL7oiZheLjobsYYG7MypbKdx/i4ZTzi640QbyAkA7/rCxTHA9Y6hHNkpD9KW53PmOs1ngG/
REQlNhwGNIp1gBx4lNTmyeAQA2RQ3BD7hct/zuBYWExRF0bIVsBHUU87qAkJt77dWCseQ1xiIRgw
QepGn8ov6BoUAH/CG/HajdlN6wTBx0cCSvTp/MWw+hH0n3ALEB0+yVV7/nnetnXkMAqa9FbsL5Z4
GZRDIU9otfj+aCSDKic6dT7FgeSTkWqw0VSZhrQvesB9epT9p8pN/4zNX5qrfHrmuicaBaW6ZuWI
Hd2jGM/wY4SCf7w1krVMT1KfCRGX8jlOc1vVZGZ5T0jBbyTRvmJqEQldEg5kpFx8bYysHcIvTPXr
7+PE7pwMIZ/keqIS05TFh0yB4VWVlmchCgd2cjaua8BtqDfUwutM9wTyvbPVKqaE5KzyppKvKNKv
rT0GJGjPhti0x3X+lTKNBe2e60D5RfD8MKHjyGxDSBwvN877I1rIzM+NXx2nwbu6P4SRjehFeO0H
MWRE0KictX2hntD19Kdekq8BD+n9u5WvkbpkFy3Ks+4t38DADAYsAug9BPn1FzFeoEVJCRzxE8mS
LcxLq172FeUMRODDP79lTYtnnJ11Xn1LHTtVlGpGWEUczfRT7xgjpdV0L/1qfLCddsHsogry84kR
HwbqQg9z7mdjKXDfm/bRGSEEbNvj2+SgUJJyNKJfDj9U+N2kYYJLtPYi2+87iHIayZ0QRqoGYnf2
R9/X2bGLX3k4ROE0y4Zo88KPeagHOHqGCLg1h+MI+O3zxuRj3Ttc6urWMzXiZ8RJGjSKumdxpDe9
V8FmTGn1EFSht4RMCjaqERFYGW7HK0UU8kQC0BLuX2j75Tk/IP1vH2Muo3w2v5l24VAj7cBKicjf
Fw0pGT8eOAyHbVq0y6dAQe2kPNycfb0arZa1OjtoHaWs+oRmoZIhRDy8xfuDUoty2fdsaDPeD/jq
BOE75w9aVmqador41gUkeZJ+YsQWyPmfbOYem9zKS8TaY79EkuMU7T7vMd0+xTXMXAQdJPbeL9wo
C7Yp1QAycT/P8SmmD53LOeNPL7XHqTLIshYwfMCrnuHhMsno6QHrO2YG9r0Lj1BszR2GvwTe3fhQ
olSx8ftbKMIVXoymJgXCiPIQ0ugBfOmXS1lmEZq+Ayd4n3YZEUpLTxMPKrxbIYFvIYDrYDAB/W2C
G+vGDT1iKQrksV6zoVPPdPN0wYFcnwnoOsGwsSO84FqUvnYpwjnPo5kvuua9EyUT+rlNBGcAepKv
ItEpjWOkxx1kc2n84U97tn+pU/nA/9ZhP7VSpR6HKi5ubfyQIYQb6PqHyHYGVDaejEZj0FYe6woh
HmN+Jt4pdaENv7286SC1KXagpVBx9YqmaBRpGVcR3iv70+1U9oWKz7ummBZ3Z0Hjpxs9DuAnC7/k
f98qZWPrbGBKxovE481gGMns+OMo3pVAsuT3eyEAdWDumcF4AyMwTd9OJNMbziA+qB32s/Lp4TjU
dyjI3MEGZF0KXwXbUHx580PP4ypssUfNfi2Dl7J66gr6ZafStw2R0n4XoFulZM4eXIpAAfKb2BzZ
b3R9PPBcHuQofOK8bFV8Imp2xenRt6uXYLs/Jd0hoUdRfGgqsVgjamZz0bsADFLzboY729BzZtLI
UpBWAabvOoCLmeeeyJnKtBInyIOc1Us70/7+SFhRrM+LGMOb4EfCE3oyJZq5h/TxkFZ5vPTjU9EC
kdyHRWdVwFqsJKJODwcKf74i7COZArbnbr1puWYGFGZjwEtS7fKV8Vqq0cumgiodc/oVKG1BUVEj
wLGyNhUR9QN8Ift7THiNlyTdeki9+K2kbiouIfaX3sY4Q3QScsU+5iPYwGSyJwCHFPUhXel3Fu+7
h/VzobFS1jD8aOX1KrkzPrj25FPMvtF+EUWsPm9vx6mo8uum+TatPLCvCEDe8bgPDEB+vgESgEey
u+z8MVP9Zf+tQcufjkn92or+KlnvY2mDyb2HSpggzUXju4nziexDYtrGY6q+qa9ZkLrY9ZZd+X8M
V8Sg65BNhKHoqPDWTy7nbkyvcO1x/PzmTZFUOjQ7etxa+0Fo6iPMN006irRfQjz3GxxB+9Rrlbot
Q9un3smlvLT8fJhgxYArG3b7fY+SqXiROab9bEp+NXGHU63mbmTurSW+NxonX9yhUWpd+G8crA4N
6Lqzow1CGyrL9YJY4A9yHhWVRiKE5GMi3sk9iyRUOL7jPYscKAg29PF9kzsyU8hkxKfmrfdQLUP5
ZKa5QiGMIgVubTbuiVWQDKe0X5oYENr0K56e2cc9NvQfn/ihwq98bNaJYX8FQMQ477QZW4Ruj27O
prZI526Q9E1YDpzH9U4sG4we6niJGTTNrWMzprQuoB8jd8WP5h5JIr4ILde+ENyaxjm9vjoMgXMw
BN+Smms5Bo/oePn4Q7C5ZRIu4D8Xi+JM3l5Opq7ihoz/hEs7daOwrcZMLqBvaNl8nbpW43KisTTn
1Ilw6sMuRjOSpHDoLp8cg5931cVNCNkFqlopCrwp5hG7a62Fn3pzvlSyZ4gx3+gS410t2NcGLIa0
N8mfBRS0PLPs9jAI0BT6TasuGRtvRpLIDE+cja/vkSIIL9RWoMluJ5kr4TeFOIZ/TOnyiNcTBHjl
DO7Nth9hSWk9SpWAIuBhnaRrFRT9KoAG+3LXhr52qzrWAaGxiJLqjwN1ZbFv0IRUgmeR7sjzxy9u
gGpEw7mi8Ji96jFv0roumR6CMrWssh2DzFCkwmjNOKe++5vCVpB2FE0XptZchI3l2ROP1F6J/ZcO
hForKZDEKyOHn5qEUYgiFhVfQdIc6vhcPFhkE+SyDwCsY+zRKCtyumAmGUkrHt2KGH9PRXABZu6A
EGKKvQU6m4vxEXrMeAVrY7M0LCv8z2aychbHB4CZPVfruN36AEf0vOwKj7oRA3+vCuX2OZwlDUhy
SgFILQRL1MOZ4E6qnyItl5A1KWColuVTXFgIndJ3QQXA8DeffeM+RmY8UhX+eNkJBn0Q1Q1rPaZ4
6HMR/WhzTbeTr3Z2evzSBccgRc4BBWtmhkjVyHFf0jjDCnBbuQOmhe3PmddkjAL1Sf9EXLen+9UK
x4U/LkdDiWju1AuqVQ/NyTFpvd0/b93WAIH92VJa53SUlC3Ijl6Od0/jLEU3hPpREmwHYnnu5kQU
S5k/qoDQcXPmxADlz2/1BPev/tYAacO4YhrxkIBoi2+Y0/XDqgfnvIeZzgyhYrxB4f6tlCankewa
GqmbTxM4P7dcZEx3AVy1lQk75zFfQX8vU5q9L1UVVBJpt8ffZREsncQ5k34+Y3e9LhoDG8rIYSJv
doVyzfo4KHrmIbfEtioKpPj6q5yN/cyJmzy0mOKu/xFdPx2XrIbYkp9G0pSeR07c49HAI4vV587z
qYYt6+MxdqMOoHbCgG9r84NkiGAsNPE7+DgkmZyUUkhgIORQzCazmCECrYzopZ/4kjIKVGPHNxUl
SUhX+gN76wcZXUgzH785o795t5N7kC4F0SsLUdUY3Y35FOZk5XpZvn3bwtv7KgpdjgFC6iKEsUAv
lDyWwR6ovsFuIW1zZhxj4+vl2qXvHUI1bd1MO3IPFfUDa525EqTMVPSeT4n6dGDf/FEI+PxM1a7/
W2txc3lsO2FpWyRR5jdIQILjtqIbXsQ6uj1aQX38W8NKEReyqCo3pDifMqUD7u6vXJ6xFH3EJb2I
ASgN85QaZ2AfO9ajJBrqDb/SDtwjnBpmUP/DWPsuuwmp0ryy8FubnvMpQmg5CNzyFs18M1supkLh
byQiOgVrr6lsxO243xZ0cksflQtstC+/GO5a44Fr/R9WBeH7fCLQkGkiUoLP8sQWRMdLTNqidfRE
ucBGLf/ecilEVlVgDssj93UT/aXJjRlaqiQf8TkTeoxJaeTanYOh0jOt1n9hDfCEol+v6oMHb7O/
AxrmvhZq9oRHX9yXNhdKWe+CwXEUlobvqhJn3+bT5oisW270ZcX5+janKx+QchHYEUeVKmzCtpPH
iJDLKghQ2uI61R8Q9SAWCikPpmi7f1+fIlWgMkyEcI7IOBC0acQeYCFB/wgo6hOxI06PxFEVnWWD
CAwrIP7pcHEDnQdM4yOHw+unIWTIGCl00ov1C3Sm9tWQJnrwDlDX8oE5+8IafKlqdMe9+v//m3yW
QGB2bBnf+sDVfKg2RD1Ahy7b6bltgSEr6WCIja9Z8Ciy/Ebl0f4+IFyqmdyh8qxU1WvAWho/f3TO
Mki1PZvAbHvG0q3j4rgTx2eH+l85ESrGrF+ob/BLg8WYq2u5qTooc2T2z6+tEKSbtD5M6CYSWxJo
UGcnz4goxA1YA+I+z2qCG5wOBJuDXl+8FsVAFKBAOwyd417WgYxMWmfpTbf55AibvWQIT7AjGBa3
PTVGUe55F5wZmG+hFM+DdNBqreTzb0cUOI5rngyOHj0OiXokL6YxNILqmMFSdoPN7NX+vboOZUiU
4IJkAmgkVyIu9Q8rCFv8jgKHmQ38NC3SreoXA34q/QE2Bv3JUgWimTqcqFRknblqSKjHUR9FjgDq
P5Ouj9Fm2EbAhr/G4LBXznw/C5vM7ClKOMAyyHkxs5lJqzXMSOHNNKN4QHiwiwBVstqrLwJC+Wmg
0Yf0/rZ9vi62yLaWSpWWkvD3cw64ThriNIo6uyNluV4oWPnC3OwlDpgORodzWN8jhBqsv2pWiEXA
dVMh84dmZ7KFLigLVN4gv5a6u+CFgZwpJ0vqNECNu/RqVcAi6RThI+3P27Guc73av2mHVvdI4cs5
KTow6OfhXUWpIG5FLMrLyCFRGsub+GAPDFLaxcwIXpH9KK7/jcdn4qt7qvzxZY2k2nvO85euxuOn
QRL6l/cV2aHUtD7TnxKzOvxmyy609b315JLyvjUYJOSyplDmpND91n8Ezsr1jW6N90S1lK9AL89h
Fg/AFCyIgyvnbtfUOjQrUbMMGPet9O0jfP0ZjnVg/NSc6akYPtWQ9Sc6f95/ZvrbxxivnAoQSzA7
Ge4ksgLk62icIffh0q9a7Eo0auik/GPk7X/3rmprIyc4hDBtvv79pJTbmysT3+SQ26ZO9pSavrsK
cTgOBRp6XYO7WCLf6DZjdFGufXhLeb69p3O75r1kl+iP5bqMO8ZjHdk4RPJv37+Cgy42hxu5upjC
18EEWDg4RxozMw0G5zHGsFWjlFYHyyeiHWACO/ZrHHNP6lUFbGDwR7BJRAjblOxZkRc52Mhsw2EJ
ZkGQqh5voiCcYDAkhXfg3tOwsXYfkS0nOT19uHuXX4pKG3I1s5xRmH6oPgyvYX8gjPnvGInnprZ1
id4tJaShzGe0AxJnT+cjG2XLpANxGxlkLt7KkeONBfnJ3ksG/9cnxLGqf9YnOF8L8B5OQCZhVkgq
OoibMoAdFE2bGEkFr2RuB3EGt718k/dspuV4xBUUovYpOdsIdqJsuiiTRcshRZVJVmS7majzYDlw
rJIffBSDzPHDlYuFfWQt6P9KOgu2YSOCf8g4r1zVQHn9dWZVLCUgztlN5H23NKiLCR4WFEdgbxFL
IWDRWNAS6iViri7CXiVUT90r1OU+RmmWJOjmzhvkyLhaIDfuQ69EHG5VogsV7zF9lppsb7/MQDja
Q1HzfR8JHYnNiiV/eh5CV4/yEDRimt23vif6qK4KtKXEiDlA4yXEjfKqyX6qTJVT1RAAyN3I81Qv
ke6EK9MA9xWPhm2qTx4jXDg/xMTRK2PdoucvxZl1UQqEfnMIKt2S7SFgAo+kq0rPxy3grsPBaqBa
LzxSN+laeuFWAg17NRVwi4aApP0jjFVjb9wGtE2NbNuIO7K6KQxuL6tbxFB2Zg1kdBx4lUs1GNK5
O9nvkYK92lrus2EZO2uavHQ7GXpgvYo4YwxH8G8Sv+Aq/6z5hpEdCwFmm91DK1vuakYHlR14NiUc
0cOulNm76wODhZwxfII0etncEc88tXkxEQXzIQv2+k1VEAgDmwVMUdnRjVdddM3jpFQ/srb1hmtq
WwpCfiq9iV2u6AmE8BNCYtyCBL6cGDPH48XgRcXoLvH8J3Jl/mr54pNG1xju2mMCXiVso2rPw3pm
GOytvJ+ZCwlmcMr04m7hnTT7ylD3IMDQx3j3IfoLF+shLunBuBkHpVEdhKbV0oXFLqbP47+o08VG
ij646KIhQ3kZHRLDd/YcMcWBW/v4Kq85zK7NAXR8P0/iIfx+zhWIQjFE+s8S1c2HVnS8I1u48Smq
nhzDP4r//GzX5JJrMJsDXLPJkuQbVcje1+FFTqHdL7n4B3s/Hy8HgevGC9aWwvmF8p4rW5kQVX3W
te7uNDUYkDURKOZDrReTbQTB14J7aJuKedw/WomwWPNYoCArWwVZ3NaFW3DxY0oDTV8wUEErK1Zx
mEgp8l88wdruNUU05CxOXIFI3Pii/Ml+aZMcAZ2I6ZnKNbSoNbf+XkzhrK4WR8NSkpT5RLyXPeUw
0edajcmLJ9DEJ44LImBOTxntu+ur0nwWL9yyHUpk9au6imZxbeol08YRJk1HeFaQ8Ny7dBlab/m2
OKy8ZaxogF5vIBRiZ5rsp3HBKk5w2rPnVw+bhfbJeWQxxMU1fgTbwvMc4IfAtHjKBPYN2FVPFz25
wGvzvdO9ui2w/ePi1HhJWE+suJH08NKAX8iVA9cBNSPmDjpm2/RkSfc4fV5aLINEWpu/GmT7i55W
L/gmgwfS+esb4+4rV0OlECyKvJCC1FhUjf1G4ic8MkVLAFUyLdFMG0g/jeAEaG+OGlZaC2oUO71g
VgXaNGjB/iTDj7L3R0wSbiTmFbHa79RyfMWHkurKVaHmzJcdnYAycc2sQbC1e1sV8bZaN5u3s55c
V89t4IuaeM2LASEgw56PsUlx8DkWDYstUtqkq1b0MLBS+6LtSuuAc+JEL7Op5HflTo/JqfeGKF/v
xRVr0huT8V4YY2cB1s2mjeZv/y8PxSuN1Fb+nw3WM+X9RueV7AHuJV/93CrVmOjoxKuJzhCfucG1
SxgNbfoBNhOXNrsZW/902e/7HDUuIlGHCMNsXYLmX+9KXafLF45HnUJPqmdyTZyVwm0fwAzGXUeV
aIlGFjpwfScHVIHbthEDAk9PveaOIb3Y8T5QBG8c5UldIz/iZ+J86IykArb3pspr/HggaJNpzwap
tt8NtWLhUQwtAhom8xSsAgs3clrtOVxRS556pt6BBrX/X/i0/3AsyMQL8KudN9hnDg0PHrX2yAGl
hJIlr6fFi3ms3oOEThX1hpuIlUOwcHuw/of8OY/AJkCHTknNdU7O/ExD4toL4c3iKL5DacQ2qBlo
fjp7cieJKvhQhKHlMQLVJccmoLtyEdQMI/jISHC7GDctLgyWlRDcbiH6CP6hKyY83lg4tJuQzeU+
BWYCODm1jNLfrWDVtZNoWjmefc0zudnhLKbPKsSo6OlZSL2rgD26DcP2ielqgo/lsx/TWRTh8869
nxd9J988/g/7qWU5jPD893mZCR3u8WDfuy78oneVcVuGhuAgNui/yt1EfNOfIyiJKoXD06XIsXiJ
W1jt/K/PVq3NOCe+offcJpLSfuRYGIh0JX4d7SDLx7BYL+kHIGt++jLjl+CbZezi2pUdN4tL0bcs
BvyrMkAQg9eC0M+I7TlSKgypTp2eLwj8+XNqlFw1ytm9H3qiWdMcGYfyr+Wdhq1ASBBNgd+2wrU2
X88c+2FeuIvOap2HH46xx7CWB8YLO8yxJ7BkvqeF7jX42ogFDi94ez28T7QbGPkbfYAlPxNk2uvQ
9XnMBr2L3yINy0BF01zX3P5/96Rq0NtciDXbzaS2W7uKzILke41xrTgdIAuS1HcUUjU6RUqXdqQG
duQhPBiy0q6ET/YBCWLtXZy3DL87IHqDc+WqQIyob4C3WEFabgagRq3tLcKzWF0tJoHsWCqv88Wy
cpYKsvKccxkp9JkS/iZcQK/AwJCQGJOlf6GKADipmINkX+DDwcSsb6lvyxVIgLhbBdoAqspFqwwY
R6dar+74CW8KbNdU+RerqjlsnmOuLqMowuyEG72fJD9HmZEHEcJKSxn9B1oKF5x4qkXDDymG+AVn
+9FeEwWHVk76vMRXrfhdCKUBPHPb2rM8IRqlHlp9C0G5YCtP3pCReErD24pjuGUwLjTOqaFMXg6e
xhtqG6FBrTPd19ji198mVsQ8T2xBAS886601I2jBnw882XTBO1raRidIQPlpHvjOi4Oc0Y6yyPi8
0Mo2YMtUR8V7cBN04jy1U8TgothFZH+dQOgx23N4TXU0rDGjFi4ZrQ6j8nH7eSAtQtV2Ye/Mvlb9
4WfmT6g5DQ8f9S1g0b/fBb1T0R9UWZi9pc3RV3UIExRQJGOboM3Q7EmFf8+japOMnpxP0KXDrbnR
PxqjFaSfmav7f0kbIbwuQ5wMxRXC/aM2bZ8C9/N29mdpQNeGvyD0BKN6nS7te6je6BVC05sq/Vdd
4RkA/TFMxUx5YH2bZQ5pDq/3XCXmrObzVsQPwkF+TNOLTb8eolFnlJVpYvP9q/sYn4SuiBBwwB7U
YW6/druHdmdbEPxZtMCMtGSCL3Wljj/TkGmspYDJZEO2zv1rBLdgRbAKU0eltzjivCGuWrRsATJO
+avH3HZdh6AlgbnSeF//u3PhISxrM3TjbJHzRVw1EYQG/D1wvBu5WFLp2oOGxVJzhiJYQ0cORVhf
6lUTvKwf43JpqzW5+K8piUZcbWsatZlkc7bwM6Hlbj/FjnuAi2j8DZ6AMIRjIqDeaJzi40PkNlS7
ZsdPLsRgTDxsEFKA3tt4QDSjqvm1wcYreUXvO8jUuvwMMnhf6MyA29+4+c14R5xtaopXT6Dqw8/3
MQ6CIEzdWL0yNZQZoDwY0Fgj4n9wNnWxpPTK5NeGU/Nt2ONSiwn0/9upNu9EtsqNSjEuGWgTSd72
1S5kOq9zRG7mntvFpRVby4hRIvzN+EHYrCVLWwf6ky2hiBh6lzyxw4SR4BGlFseb4yZpWTplj2OM
uh8lr4FQ8D5CoFMfZ0uo2tdkpMqs2jVCjeoArlSIwwSAcnWuPNJI7bZIOhuSY4uTD4bjhP+eu55Z
G0rZdhvODzSXbpQ8aPrInOMungdENeSFuWvF1a4Sbde1ck91jbK1Z+vrvVIqo2e9XvuHhZGVKZW/
GjwRMfEcW3GuP89lB6giVjfW6JoMjVr86zrrl4mcfKS/HK+eNQCRBLk4Pe21M235d+vNXXWzIM6D
iL4eYl3YGL7TKUMqgbRYdFWubdcBcvfZTFTe5BLyJ7MTfqZteqZ6VzQ/9a2g5lkJVVL1E3/qQLnY
GHvzE6x335b1TAqmK7w8Sl2XU5XoeVnfz5OEXVuTGRwi7J6Ge592Migf/zg5Zsbs+kcYP6QZVdtU
vmQjKAry8YSX2YZaSweN2RFGKzJ1WVyYO/IQxTv+WZxeZMD7iN3LDdKS69cVTKd2Aq33S6PiAZBc
dUMOc/8RiQzZLUqKJuOTmOK9UmGybbQmA540SDgIz5Mb7tqZ/qcXMWILOjKwkgIyBGYkAHLjh17s
Ey9dI8xFrt3ipmNd0xHhTm42HuwiauzCjzG9JS+MpN9mGdscoRhYEr+pgKzwrhygi9gSh6lX8ze1
S5CA5kHgV1y2J8uPnftLT7d80sKiC0K74gSfjq5WVZ9BJEx6HNUS48xjQMCEpPRsDPo3tKmQStm9
l/8yeTqLitEe4YE5Oc5PM5jIkbzoxY8ullDuTdpkEAuynx1oaharPFuauwSJ+sgoztkrubjPTJkK
ISVEQwlbjsuLf70cFSias6AoSS8oDNOwjhGl69iMPwJg5j2nC1XnhYR9iEzS7GfVJZYdmyn5T82g
7LIrtZvs3+OuztyUZ7soeFH+Zcce5xaYf62SxBrd2Zo6WmXr3wQ4AmqAPo2MCyn9zGDYnDYDSqNm
XtxAP3AeWxbpriTYz+Lk8sGZrRrcc2HBBkgnU78jU3NEMt0QmkYBh2Bc2As3d849NVv9IJ2h80g6
CH27K3zDwN4v0BFdS50cLAVGRUKBkHFrdXGWkAbo3ns98GjWiMcJCUgTpsKkty4DxFfAyxkQvYul
P075uqPHMEcE8o1e/8GHkxwdMZKwTbZWzqhMOXf5ke3r5abBmwi8DdOaTM7H5KhfRA1llS+1QjvA
2yFXnqkqvcL4Xu3wPfJP8b+w6ZdFkxh9rjlvL6TVtT5Wr5SW0dzLyAclpIfpk9dol5Vwacd9/I0a
DUFiFdjX6nACgtYB4e75NQLTUrz5IRQapGtjEpF6b49rEpqyq0DS5RWx7vuEmsIcshXLZDGRK/eU
1n6NlT7kOqs1IO4sMKww3BTxZIrSxp3eQGU0eFkUTvBvKHFVHKfCalug0nTrkCr3lBJrUGOcNXOB
ag+f7sDIYAzJg7LvhlyrXsqxauNrjdO1UK91WlG722g9+9cHiKX+ILsZJjCYUQGRBMMgkX7KH+OY
v50rWeBYFI1eJyK5fQexV3Lygcpj/W2Cuww4c7E/D08vU6VoODyQBIN40l+Q2fjvbRNamXq+5Y0s
yTRP3himhHwSQ9kaIZ5TNzVCMIxl+lYpZIROF51u34KaWM/S7T5pUqAHlOz5k82K+ZOhzA668S9v
uPDhrBimHzH9jfl4NqDsLB9IcrR/2vpOT9qSc+Uo/pUupEB6dicwVA/DHqbzEDYNb/s7/tYfgnzr
CZFCzzehau3xOtYidPb1jJ9OQLgguDvaCxI90eA9ByA+K74CTuq71wGKb8Tj/V7LrlVJ4flJs4t1
OlZalJQ+4qxw8rp8mCvFRYEMXBFbNy6Gk5yzzR72TQnzMRNa4tUenGUYG9d5Y4d+rmKLiC4UD/lK
JOlbbglJHJRQgnLM0vXQp+d7FHO20xlqoFqAyBOlCDXO1XFKNzN8wS51HyqGkSZk7FgX9V7g7shT
DwYPwMZtM1J88l4OS3cxd5wyAY071NuF9gUo1CyRGAXnYZDNu9T9/iCKhU7WI5kc6KX0aVex6HUq
DLw3QojqyhTTlJY7VT6INqgl6nWyre417ULGANTiuAHxlVmwa3AipQ4+uIG6SjnBPgpE8nwk4Rsn
CVQGMGXC0tDezLwKRm1fomuwhEYToL07Fm3tzaUgTWxAZdO3SqzKTx/fKUJYs6slH3Zl69gup6ep
IUIEuUY3IwasWDq/cbOAr/bxEiAcHNIg0mO2Bke0RCtLO4fjSk/g37CDr80stKaREug5darQ0MhP
kE+Yae9rnYCWX+dMcDZVOOLE8mZKYdxdxzrQk2r5J3JzsjhJ/a1c9VhbADrSUPI8hC2+P35bIQ5d
jSPTZqerkUXKvh0gPXMbzwPmEoa+hWk5vZBz0jR4Txy26DBUoLw94R2w9RDfzq6cZamvqH2daf2v
vMFogiHZR+3x1f2MIh8zPzAHpvdPgPfqXvKTbRwHp8lfH/PHsgUG9Rs76QwL8rMwqRq7eZzFDQPg
CCPdzOuL5HojA9vHs205TJw2P8r1t4pMpHMOojrJiajAS8tOk8kDTZsUZifz0Xi09dYKS2FWkAOQ
PqflBqekEmwhBv7ffzW7FJdXAfuWxyCu5v9Olw9LE/1bSG96fUqIm/iQ2+aa3gYSBULoE2eA4K2z
+aVTJYvg4uKER6b2vJztGdqiGlRcNsY39mi5RjIsdghyD5WmqR+YBLh9DI68W0TX1IZ/en4MXyIY
jD2jdVGOqEOIAq7/9u2X0dtsAlMaTXn9qbTTsx0e+/p3UDIWsbY9ZrSKouQdMZi8HCgcsn3cusAn
5pI4Df5vuQkP1skekEklg2qRZtgQ1/wGnUAHI90chujj+wOnCvr4dMPHY2T4I5eA3yacZz/3rJ8c
ZlwrUUt/kmmgJfkGobLqXaXARyS2m1sfJFMxCDc2/nNy843NgBUcwLBVx6tYUaRRtgQd1b37HalR
eYsFy6e6EFqysOsakKWIqhHgTncAHqLuRxvlaKApkrtjsGiAxQIIseh+OwKG71CzhYoquVpv5W3j
OHh13WDr9McU3t1qjmFM+4PJFIHGMmvr4IbANlmOJE/V9rnL/psBGQ0qTVEAefr6O6q4Gw3n5UVk
7H2teIslO53NlsEZSFgTo4dKfRiVxzhEUIj6cKd8oxdd+GxZV4Shm5AhGjQXSPtxXCZawu1iiWyB
sXacTIGBeJFprD8b3ztBUa9fbVt1y2z3AuBqqyF5mm7z6zdEBIaFr7y6q9c+lyMyIO5r1ZZlERKa
SB9s7S8aOBmfBzYZKYZzF5kDFMgELf5kfAqEEuJxk3wVHqIzkGcP1ZfdGCrtbcc7ifQ7dfzvl0QE
c4fzA+OTCZJ01vCQIudhol9RrLkZgCPjJRgFYtNSQf0stVF38QczXw/9Pvdmw1wyg3NTdHE5Ii8y
u96fHyBk8IuIKspocXmKNvIyAOs5LyBVUeUJE5WEf/MMr1FHcmmXmXCKjQHcSN5CIdgAyn1G/YiW
JzWFCHpQfiZ/ehp4PA57ZQB8Xqe3yCjIowbUCqFdkdmQHS3AHxx/LA0dCk/hYMUQ+hX68+E2PP14
ShxBgfW+2qpdxLo2Lz97SPdIiSCP93+qHVXSE364/P30QuFpGAjQ5bljtl0OGXffz6AEpf2C/g3m
mRAT1JoEbFmKeLlyMVPafUZpf28x63wYgklFQ8cxlg/ROU2s8JkjDpxZWRWp/Y1T63U33kkTi7sY
cibo+B/FeEwjUv4hnvSqTfHZR2B0+E/OPBQhDzanhg1axgjtPKLNo2a0898n+6p7fPN8isXV0+Us
YvQtXipNmjrTljGHkayew75mUztDIKcLVhtCGfKfcxXETpyPQHrilzT74EGhASEHdVOY/VshYpwr
tkmg3yfl8nUxxWgefgZifFPTW+rgffn5wC2gAlGzp87OBQ9CLtZ6CPFmiX1XSaDjG685LPJChGn7
sJFbKc321RS15t32GPW0ByrkwO8Fekp+pGQvTKJuxING/Bf5M5UVGLcAM9dL0cGOffXmuAAoO1ez
gwKEfCaqm6UsSQwJ8OpW4XBkwUpGjdKF8mc47ieIkzNs24/Gi+iooFZ0P+Y0A+FvNKcw+M/29tvn
ibcjJAzYyZiT2ESmnzwO+D+wHgOsreqxwQpT2cyoIh6a/ItE0TX0e4am0wSdMCGf4NCbrE1y7WhP
Ai0wR637Q7c7ftQqV/T1atcaA9Vn3clgTDtqkFo8FPaUH4o8K2SJULIJZIHSnAJCfPdQZUKSRsOy
BETQjhMeeDm9zgoHKNMZSkqCL8ROciATSPlz00yHVGZFyI6/EYZsotHpgiqiQqkEZ/YnPVHuXegy
j65lQJk6Q8KQSWPcVXTzbTfnc/wwUYJmHqNHSjZAgviIHt48h2qgX9q7WIo/fqF2j+rAEAxXt/0a
ohTXMvrF/Gm7fMwQHude5yDqr5kaPiNPQqjfkmj4y1vawUZ/ecJhzzhmhbbn4kFZvhlEQWOrob1g
A0EB4PlxXot2glyjAOaRv9473b54teEWwk/z0lLiBEm0xgJrfUtGpovsXwxUpx82eBnhhfrWkAxL
wWiKfZejh3hEqh9zxSBrM9gDyGo/TLl2d4csmgz0o5JWPIdqzNF7JIbasJoEjr2Ifdqu6zh+iny6
N8vjF7NP/R6rT9mECc3XvRbdMp/CDosvb4xAyCv9UUmpSCcyAoR5RorYAZudKtWkwqCnAuADfZG5
yNQxI6Avq3LC+RIE4G+lCWXMF5xKnzIeviXBIPPcYuTn4FSb/2/iUhb5GhfFjcyWmyKN97idWeWx
0kTtsNxA3m6WwjSHFfFeia7d1qfy4X28Zl1uJ3zDoAwmCDbLlV4GsgXzZXJEHvtaObolTmc2I81n
plF2RbncG03yVrwlPBslI1A2+f6w2ZKU9WMvos8UnAaVoOcZj+ZbFbKHbHSJGZWl6HY1gehXcJa4
PXoG9d/vVdndG/+ZEAA55LtzKeCjZvbugwYh04/eQM3hJvsW/5z8x8pNl1EIxdz2UntqZSe4auC3
VvefS2p5x3DARJ7em2MpPzoeEONcNjl/6RofrcwlTAXxWVWqP1Qz9yfkua/Z9QJVZjlUBilkOMBw
+dRGhL4VxuE1rc0VlBGIoua3pEq68VViU6NDlcoAhsih6xvOX98rCEOx3g8Ih4J2UF+xUCV8j49K
VNCk7pGyEaAmWi21cR56fRHXVCLFh9Y7WmbnxBk3vUU4qnYVc9bW7ttumt4ExI9e83hDWgUGutr0
kyepFN7H84pvWSgUH+HBTLu2rIS2vqWrzFi/t93XdH0+aHg0Ff9Js5t4+8Ys7SmCXPIkyxHnhmFb
dtGBI9wPq62MZsaWo3ltinVtH4LuaqfwzHjp+FJdzk3lcFDNHAWzCl0wv/sP9tKqSQQv74GFWga8
0fWwv0RVDT7LF65NPGJfDwjrBdztSl7JRev9iNYlLS3e1TN5RsOytKJ00OywvOtJcdgWXtdAYpPq
5yJPu9LYBv+egMKYxA89K3jMgJtqKsSsfhVKEG0ykndKR2HEs5z/An/WxYXMEVryyrK/MTM5ixyb
HAf2q8gRsRe9y0nSj24QFf001glAhAypxt8wxG1B5LInaD4Hr6fW1QOMk0a0u0ooovLjRxxadjvT
etCGJnkPnmDMHjAQjlT5+tM387GkaIfwARcLUn3jIKtdtk62c5LiG0aQ/0MHnkOo6JI7kLRAuGnE
PxBBmw5dSveCBnbPKVBBo8+UsHxLYrvKdbTpFMcvmKycE8FTxI2jM/qLW2Edguk9Ev/74qu8Cb1d
PW56+p7EnNxz+SNrqMeDwQnJVz1roZDCTaqyyY6tk+QwNjDZvIFIfUYgsk78Cs0O4DL+q5kiY6jj
P8Gg05geKmWB+u+Has5j2S4rQODSWUxdyLvY40q26Zv/uFXXlJOfPqNgtRbonxUS2efhgrR9W4k8
4d1JjhEltv1Yo7jqtnuwkdx9UJjTv1yWT5/Q1AUFOrGdvcyIYr5n/xpmbm7pjDekVqO1Qdl7ghV7
ydsFXRkIssLYdyY8tq6qRMWAwfDGFdJXk08rV+NMzVqxuQE7Y2y037+y0kkff4rB9OsK+kT/u3EB
3KbFGxc62AdsvJTy0yOMK0PA7rnts5ipjER6uKGv4Kqe/Q2rPxc3SVz6AqHWCTX2kcR6ws/QdHhJ
XUDCcAwxAnu19IhbutlXxgxWQ/cUR/PkQxiVJFEtCrTTHSTw9/mCpOWLwqhzL/q4tDarzaXWr4aF
hDMhUte+5Il9BdqV5tryNJFBR8Uvuc1i4eHGqH41Pn//3/DhZORPiWaRNIyusVTJB7YKK4Ridw5v
/aUXsAppoaMdbh+Nt1oUyxLjN89MgrEpqEVUG36kY/hE+PqUHprDSZBxRhShURYobyJPcIfR10jL
uznwBhoR55WozULLvIxz8RrfxOuMytw9z1R36RCOzVO5BNTfi/OJf1/Sj9tj7b84NqPh+kM3l5gz
sjBpfNPXf7corBBQrYgXlgLwno3l/EDkt1h/8ayfbIcZwSJJmS7hqA3NpQp9E+zx0n9OOQWnsce4
wjew3SXMpCc7n20bvwfbqUbElX6JBUa6hx/fXPslXmfrgq//NAsU5nd6R6fZOeQmkqQfivNiqzmW
pdiMUkPZSW4nA/Nk6ySVlUZn+Ywp0yrcnGR8oGY3Gsag6Fdeg82NJLLtioOSKxfTUJPO06jYsl+d
eTxVxGpZfDk7iu3xbCticR51W/dt7TjdxyCyn1y88DdRw6fAwgZbnv/4C3lhndNC1aKqJJwPsNoO
/ZS06qwXET98uK0cXaR6FAk5pYNjFsHex0WpDgF2h34rBhz6f8bl+TWlmNNOzNPWMR867Gvd/YnA
PyUC9ep8i7cVmJjBWpuhzFgIZXHY8T6ES1S/4H76P5DVxN6Eg339s/1vL+PFS8Ib+H5+G69UakJ9
EbAwEM3vHEMZtpwEpr4M6UTkyNcEfWHY8j0C7ODL0jMoUwQQyaADloA6+LtKmZhfee/JQODNgOxt
8gWTX47hAJm1Seb+9Hl9/HYl1chDJbgBosfyOjqnIV7mMCcHOtgyuKRea532qCq/EUzRmIdNZmL7
acjZEYTAYZANzv2y75kdPKsQgU0AJ05pQzOod+iS0aO+rPBihnLGeNh6p0XutGHGhl2az2If1dq3
EKRGm/gGlOopPVFWQpib3gZdplwLkXDGDj+nAZ6D8RSZWqRO4mXdPEajZUdu08Cac8rszW74PatP
ZFdm+rVWM+XhKmW9XSyWJ/IPKJ8zwqjIuoXn9WiCc6Tt9SqZhqch8h8Iek7WAq8TJdPrNNzac07d
Y0KzItLjhB0OF5EV/Ok/TKCXPpZyGl2LYFwqiZ2phrtkX7UYyT327e3cw0AcTrcplhWvQLNLOXdP
hFedv32riFRUdx1UHHIPoRbzPYe+D1T3RgVI7BGhysTHtV4rtklBm3aWE6jFX+kv3eLKIkin9NZB
si2obZG8BFGFMVuWmGgCaw8VoRY8Fi02u094FUaggPNjWWJ5wc3fo3wQp4rjA36CCyYro3x79nZQ
Q6N3mnFlimeqhoECF4xg5CEuHcsMaUp0Nv27C8f4AnMJwlhVNgDGsJIUWeXjdRwQ6XOkBmZCcBuo
0++Y/kOshFYoB+MyJcVkLnavT88vL4nF3u0zAN5ILNt48LOTWDDjk6EUINC3KLQGN2ubpFHClnOQ
Og3eVS4ekqAoPCNMHmIfaWlhopyjeZtqgwSG1za5XQ93dhfd03Nmjoaio6mVLUPLF1nxvF2zD4VK
cecSivZr9nL6Jl2yGPmoNiVQ+4aQQZh6q89rzWEkyWcOZFAZAbXfMuiWLfodzFzipdk5utYVne9K
LKPOzo1q1c7RNaHx388JCXe2rgRUPEq0TIWZFrlafGZiLKr1/bhaek6ljWtSrGbT89AcTOTdUZ7j
0acqAKrpp33Q7FmpBhzw8X2iU9DgAa14qRITbkeg27BhoTDOmg1PsOz/bIqbPCCVxPqT0Xnmr6LU
0qhVqBQ+HWp9jMws/M/zEd1yJkLn692uMOYLr+BQDZB1fkA4nUBlIq2I6aKjX4RuVb1cnLSNNUg2
0IdNynJ4DKI68spmJoKH76yppSZHFtEBA3q3nSGF1vVDzfxai2kba9i2dBo27tBsXx4Ix5lUrziF
cGQ90k5AanSEh9YDyog9/8lPb0t9l2J6ifo5EPzYIWI9zUcL/bJIegVpHtauabZqYS2s8sB2NW5m
nw+nWmWRE/i7pbJozV1bohVT66rt9MR+QRYrw8VzVJBaHMjs8zctcU2DqqhYA94c4UwcrESf/wNu
YOmsmcNnWhGIVKTga4cDZIC1jGipe2J7MScQjnxNRWzRqkE/QVMIdtLUJdKHH6yJHTXiH0dEWu3w
T50t9D2MR3PWpIe2sHfvJIEQDr9GYLIPAzyw/l7rnaJ4OmKciy8dtHfCRz1ZN/ShEVEx4CmHnzbx
cGKzIJ1qtQGYcGv1/IEpsq9P05InmJ8DJLXhmsBo0XU6dl2av98NFxNUS+NXZRsu6IcgfFg7jihY
/Gj5YjlxygsO3m+bDn68tgl1YbqIo84j8uh8nob2PLtFpYoLxreQFpyNtPPuZTMJjc7M2nNzr5Ou
hUVH3PUBERxt/AlTkknaYGYz4tyywRYTwxIRKP9yXwb2Uva/H36OKzImffVbXxmp3zpSL4bjAEA7
38AvT2gY8yROmcoAfJtBekiLJxNbX10GlPe3ZYxhmDHq7g2gq4dZCruPesFaALUcOD75BwzRVfPM
HSj6BfvQFh/TIMmtBTFF6e96vHy026MzCiN049Vnqoe7+UQWSjp9LPs4OO80nu16ivVBrbigvDsP
aXflkVRjyzZ0zA6lu5I3pWcxkZNpo96FYDgxfsoq9Kwkgja11vBWDFQSDhdhX4Uky7iiwOYP4vjn
ShxooYl3P70SxptrRhTE3eQ0rRmvsP7JXpDB4O6ri5EvjhfCupz21iy/mVt7BA69pcTsjuPik/5c
TNyai/Zh3Kg6mX/TuRZueVuyKjGeOeNigtmUhkl00QrEwWRiZFgvL3PfY2cTyW0xfvfJviXvDDCT
NvmH5nikA3vyAYbmwlQLf5zdAG9cXw0Lmh6QdlDlt4h0yVbwGojdxm2we8ZOhHkbU+NWxGcPJPiL
spTtVNfcWU0Fv5+mdayvQsklW3aylQzQhgo2XckWR1arUAzLnKvZQfqKRZukws5gG6cjHvXPr1VY
XZnQcHJ163AvjNO9zm5SF2Mz7qq0vYV0EdPSWuBNQDbtLIR4NbP7wGtnlyY/Tx2/+7zQtm05RvTq
AG83Z8xJ7KT3usywniLEOKQ3vRAinYszgzCVY8jTMq5XEJ09oXJzZ06vIXspYD7ZQhhNRMOflOnn
w48L9tUp6I6pEV7obggrdefF3phiU52obXWs+7W99lQFnT1aHCADEqha9uDPneIlxYY0CaNv5eep
byHdwNhkJOmV3E+0wRhPmNiazQ+BwLto2vJyf9jLRuQv+4d2hdZpAQadPgK6kxuvB0uVxPR0sc8q
DjnfpKKnyKtV2zg29gptYu6dCScPYjTu+OUX+RnPa3MIpzcUedcm+sApCB1Q7hQfvoZ31IUmNaV9
GozXudaXuLA48pcQT/KyJh1b02yJ4/OWsvojdop8qlSrDKKJmjQJx8GDdOXqbtZUEBxF1Va959b0
v4QrQLSGiXiyY2qdfc91d96YK2s0GLRQxTgCrTLr2iW+dox56GFhHPZav0w/dYPLCjIu2kgZWXhA
7c17wVdAbAlXOSrDUCP5uYGeKTYYq7E/975qB8Fs5BayndlqU2igk/me5K4Kybm3m6flBAkwyKBX
fAQRsJdkqksGH4BZ4+4bHwzB9oh2SzDQPAZVyeTu/IxdkVWmJ3Oeu98CunXFY7u3And9AZU2dH+C
jG6JzDC5tYMxfbg46utB0AB3HpFK8jFj6p53w0TYKlvIZ6VEoCGrYG7bKV0AquUt6TPA9INAnl4b
03Ba9WFOpgTiLt7rTdkBJjkE+p2LHWxfQLoFfIdH3tHN2JX2PxTWAI6v5D2kj/whSAPr9nzpEwdz
ATTXOhmLaHDuto1Qm2t4DNutSd7Ql3WXAKYMs5lNep8RF4q42OLnTbUuzp+QWSeZ8auNYTuqx83n
0lsq1xLsUHuT+HJ8SP1zG0PT1pb76NqX/QnP3vxFUy+9SlbgTdCGLpQOrSgaXDHJI5kywvXeNISY
Gov1DNTW1E4M6gGoj/pnJ3Ot8y7fiYQqleUfh6NNjKufbhaSLcR+yo0Tv8On9huy44rY9RbM/iOJ
fhLy8jQ+rfZGLc6A+Eid0DSOZlAvzPb6f/X0NS/efWQohRE+dh6F3BsNfkaqHgHI6EsKmjNT+xSh
JaxbSCXhOtJU9y39pXrKQqKO8HEnN4PXuiKDjfDaXbIET+2EDIpdOMgB/J4ZGt8j4wHr/B0zM3Xy
5CXV5OI2LTaFIO6zZHt8oGs+7wNIgNhnrx3NwXc9TZdgO1fV6mUPN8QjlGP1maUUqJhlmNIuVHFH
uB5s0rENFO6TK5cVbDEknLgJfKpXZ4VvY2vboRzTCtMW9hUgQskdRb70zU7rvlzXJH5IYyC534ln
pFVDKfNmsiyVjsAuhJIeYBT6VhI0eWfbCXszTnzaNKePfmlA1opCi3fo5G+nfyzmSBitVCLg0o1c
iE+qb6uzr05hyHaprU3GKecBCYw/uYNNov1AVSWZhre3Scvvb3sypu9ryjUfDGM2M72oHV2Sx6XC
3WBkvA+9fdj3CO0wgVXSsHcXtWSW2V7rYZsrIY/hnNpu5uB1dg6Ar1upk6W1b3qEgtE9StYWv1AJ
cGqxdXo4eMJcMeZQM354R/V6MkO/KuQjqo7DO3wNa2pieoM4e/hx7gw9KGlDJNso1h09vY0PQI7G
90hTwIL0qC4auMmW8jNbA86lov1NbAznCZkwWY84dv7o+0Am7mtmIcm7JB7vQ/o1AnrrbhQaPJP4
DrsWZ/VNXnUIaKQ26mdJ24CS4lVIlz3IpAyARw6LTNk9Iu5Dj+O0XtkOuULCTKPwOkD2epaD2DYa
Sx+C8KJvUul64qzseEaY6kFvDPrlLsDGhonw5bf/BKDof9I7crAt5AnXolKyaHLPHyFWnY2VH2a/
q0jrBjl8T7+qWejSbH9gjjxWBnSE22t2Zul9FK6E3XBaU93g5OzrTOTU1pVB1qdNPkuzQSo4/T4K
IDHF6lnncpsnDpXYpTc5BWm0XLFZjmupUInzOtiu5F/2EwBylV3pFuFwvb8tX9/BZf3uAOjbKH8o
ZfOaONRLri3SAD4GFobIcSRMfKzw5QqlI7t24j2BZivnEwm8OzCyG5bHZiyS3dhWeMeAzjPUpXnX
mAkoTJNCBQNzn/e5lRZtbyP94lxgav6H0v4roQG2sp8qAs3ulL/scYI0JKsMSDcX4x2gIIga1VQ8
JSh58DQv84PQabUWea7rJA+8NaxQKFLdKBajsHzaGEEBOw1zGJtYKbo2oifEzep12EFhxhS5jpiz
d7mkrn1Uv3nCzFg2bhCZzINiQ7iHJ0JIVZrfoiweYE7npvEO0xTbE4zK3AE94VC6gqF59vterii0
+KUw0Xh44AQ8Wd33+BHcfSC4EhGBvlza6jGnTanmeJbmKFqVCJQqVhZd/nvAiyxSUmBmBIAGOURv
1Qf1SU9RSpJI3TG2oly2y87VeJi4wDnwfvkzPapkXjZida8Nct/1OEOe2qH8vphPuLjBz3DdxO9s
HA954lq6Didnl0QOVlFq1Hi0vcMTdHGCFzDBFFXFvizmG+/HOU85XPCpVhMr5EPafJQIJlXdgon/
YaQEDeVm0Uo3FxE3ACwPAZGVRV3y80kA7sUu6q0z1A8AfH8IDwSuFiPDE1dj5nwUeC7uwqO6kTjR
bJXAHLbhUZtKn1U0f1MFXg9Rl7wlEkf+tDRvMXPGQ1P5e+EKcqB8YBorJ6f4tRK7drN8fku3ReZa
dvku1OhxaNrpqzQFNXmszvi69NK75TVJXuzraVkeL2MIbiMPgZ/8zkaJMjS6z1jtA1BKoh1lS+Vj
dOzsFZmP16JCxPxhxpF3USZ9eQuv0FWXvayXm8k2u6wATF9V7FrS/xNErFrAAa1mjNK8mDWW8Vx+
WGVwZcx68qfsGDJwfUGuEGLx1ShxYIQUMbMZkFSHesme9ZVoscyd4gWDnU1JXy1PAKUNP4EkiG3p
oybvN6tJayZb/D1WfED/YYx6lqZwRwwMREL9IxHcj+T38Dlp35SQMQDSQe+4SH820gXmkWtpRrkx
dPEvvx+Z8kWpsPcOjScBkqnlxAIbZHCBL/yBIumRfA5GW2UsEafG84Vgzk+tehPwtTon3g5ztgCW
voAiwx3PnwITXz/of74YQYezvA/h2/w7YIYXyTx86TGhdrshe6m45cwxY1Bvz47jHbzvetVIPKlB
GxEWEDvXW7tt5Xnh5eJetE+WdFD/Z/3Iq1fM+DTvzvcD6db39SIfUxRy2FPawJRXWAVnRkkEGnR8
imV58zpGR8SE9+xxPiaGqA/SkhfWYt9fyP/WbtAMXcma71pdJ/8srYSX7lZsfVOE03yHk660VH71
1tWeFqxiWbcEEoWaZsvCVZfeeRlzEEaKH97eqqmkkqqee551nJr+tKdHJwqIECU3Un9O113BZrz+
eMBxHPGznBuptnePqwyptGY3DMxglYarYs+bzlq76mRgMqd0lBah0a8K5DYE0coqCUw9u55RTF/m
1He+nPrOlt0VfvM3clUfMDcOzpHp5dozG/ufqzQpYRYyUV0UNxR89v+15U88Pp1smsuru5Ds7q0s
Gk2KP4Sehcr8I73Eu6gVMeCscaaLX0/vCzqz8Z7TQAs4MrRBVCniu8FpuCya23fcT7x0DnVUbLJr
Ely7mA3RJoLFa8Ryu2q04liRpP+9EpJ0Yg1jl3wEqnpm36i7qFgbwj04MVjghQiFmhoOMZkes7LL
7Et7HOAfGOclt+cAyow3JxFaUwPDbFrEZOzVDo/c7DuLE9hNHd09VGzqf8gvOslkiYqkE7VCTBhn
vHtN/55xZrfa7ZzhsveioxUWI365s6Tcs51SSKh6n35unMnjt/8nOwo+noxUDa9ymO4AYK/LoMG2
RQ+FcSaDOl98YTC34uOzoO+ZmEAD3sECtSwpJsYnhuPeloQdwa82tIW+GS0O5hF/MFITmjq6DAr8
/ReMtwoXSIwsk2Iz7S6vdaumAlynyE5marL6mIDWQaesbhh6PcJguoQhPpg2OV6JPxA5NhwsQACQ
gyje5tWBANn18YTxFCGHSjR/KJrD8jx3y//bUGDS0t7yWL6KwwocC9T32wnQHjjWgR91JvU/VXdL
8aAyja6Em9+TgQdhBrYOMmDyu0Htqj12Pl96BV2vbMlstIXJIAHo4W4yT0xfYTAHUwIRovskpO5R
Duf0nq7y0KCFIgglSp85Yo1I2SlB4UuClSBspsk0xaanv8DeXejzrlYj1orpnf0Fjq9xNHFbp6N8
vFxzV3Vo4nJ+QBoc6ZoWySIaZLa9MnunRdGYX389ED1C3ycY1WEgN2MRFiXsymfIR0Vf64hr5drQ
Lb5u0GZBJo4DBB4+Mdwdb3uQ38F11Ic0bEGZPFVtg0lkD9Gl79qHAelzyIbuSIQmbzNh50EDedWY
GkWNPKA88OE+k+coxGTVEvopX633hZqXEF+D6pQdOYyrrZJu5kJ13sZ1uDqOIKYyg8zSbS3PCnhg
v1OGagTfLL0APlF5inuvem7MqU2hGrC7OYC9jHejlnBHXuIHT4RWUENu5oTnfCL1npuEXYi80BcQ
0dc+vlymlByQ+gGOICeYss5HJ7XbJCJXpFT1bQZoVzjQ/8VtK5PpFQiqtHJkLXk1R1W12BMVNFsa
MuMhV9/W2LJVbQ1B9bKXOfVL37N/p5oHatb6ojwfdHL2L1JPc7k7vmxjnfmUfKJEHcLOIXRWwbL4
Spi8TEHUYtCfmedYryhaMhLxl1m5/TgwyJGO2i86K2gdwbRQoQMJakbkxuOFtqL2MnbYB4gSJDZ/
7o5Cun4XmQmBcV97SUpaYD4OsKFRrW7HQsepwwfrgYHUSOIVANIWapi74/iwg7on22myd7QkcbyM
kRdVxSm8vnto9WN81FgwDv6ZTIhX41Hf1XqKn5+zSXJ18z5oi08WBKqO+qEW2KDfYc+p+FR/XlDa
jh1sePBPfDXzCwPRDYgRCbUaEW2fFODe4SRrwxiG9oqN4fC5rYQifny072Qgf2+N/kLwqP2qCRPM
KI1AzoDIosfHk26utcwq/v9tnjrcsdXrid6tG6zeHNXnoeIg94Z/N6Wgwj1WiVpiUYubWGBbBd/Z
7fqaC4tv2BVK5lfepEJjubg3DI4dm8TcRCVbV+HauqR0J1Az0NbakKVqyVC2RwJxXruIIEEUGeJF
2Y/vNH5NUsoLDAUxV8F7TZ3/dANYxwRLSJCqHWlWM/zxhuXlmY4b7uSl+SQnOIiN1DqMqgCxZAbL
ePGojtCeAxqh/QAoAKBZLRjo7EbZ3T63jefSE6y5P9fF+WPPMN/zjPXnr+gWI57oXyV6OQCLHtwl
i0V/M2NV4UFf8j+qxFiMa9IWCjmfypRkDyZhkkFzXPcBvv8EeRhsicNlGMEu2sD+ESWim4mKXVae
RNsMhu64qDmPUvt7ZhqcEQYoLqBK6us3KuVrDXoH9ylri4boim/JxW39g7PwLYf4pN9+/FFiJhQy
2EGVkp6agUSvJwSDn6jJTbbwNCG5Cx4EuQrdtlZm5OouIfUZ9IS2u4jtAr+uU3sCG2M0rZcIba3o
0MpZrryKRZ2qpSHb17vC193N42MykBzJj61DDKfmGIH3tOus/La31MTytQX+ws/SFQVxEzYzdFQr
Ldjnlw97+GNvh2P3oQbX1z7XV9F9gA8VD38zYZYoYPBO1WNFHaX6BW9mBkoMEjT3EB7AZQNYBRMP
i+PdM416UmdnnW9pmmerf4c/H8vlrsAfS5bWcPQgbYFsFKsyiCp64gB8otReC+oZ8rG3/mWkVSbZ
21N2jPFhGoH8vKtI1FkXu6C5JCiWlXRSiQexmRp/lFu2AymOQd7TvrAvXJ90ENdfJzEibbpV1H3/
x9I6sRmwQ9EX0ug1BhHXoAE8nwpRGonv0hk/QHeG19ZsC9lgAFkeuIY7lE4LHhRHEV/xxm3+FHLG
/gnx/FNYn9x+GN9M1Sc8h0MFvTit/S+//rOku+ogXEgmU3UVIVCuC9CPMqEgqMkPqV0cPX5lG0Nt
Ge10dnWzcIaxYuJf/GIPP9D3tiVV62Ejl9ykbPT7H9cOL2cXsKetu6AuuFGDjyVZI75O0t1sVqud
BO22ijFrml8RbS6fVpDYTo10zSxfJuwuMx5TNYD1RvLHPvmtJ6OmYqMJDldoi8r5nqoRy9O79m+y
IzXcDwcDfNdFwfcM0yescfQoGARaX4AOvhFWBM7p3rfIX/9LVZY1471aq69idc5lrI85J47BxMLh
kWsIl1zpSZQjAfvVKFubM4osjp2zDkqbb/ECHuc2fKK07o65Bi544rgg4q27MxEWy0RWZHrQipWO
/sDOqwVkWk37Vutxpjo0OkcD99rN9plSSEaPpFKSCXPnqW+pniS6y4SSxdjT6iazK/ZR2leo3SIb
oFiGT/P/2Grzxxm5nVfLA1RtlRbtpksGm0YeTMayYQi7TliqTnvBOQgI4gPxuSfuu5ARQqi2Jeea
9J2AupvtQgXVnv9HR2aegNuEjmmbpyLBzlfX8wWllgvNuMyUH+igzN5z2lXCwRDytH1kS+lGvRj/
3k1sYcA/P38AJjSl/SSmeXaxtbHyq3T1iSowxPEEgLT9uWXD9VAcQJ2GPxlSSXPhG7npWIuL/0gn
tG96arzsPSjIZZDWVTocBeguYXW7l2jFCEhW/svYFXjDUlJIFFRF6cgbjrABztOmgA98jaFoLLIz
1HlfwRbeGe/geWY7zysPzHhEMwCAgfmxkSUqujyBAf53jfT9MOVvpYJtsdszFEJJyVtuoW3Cs+u2
o9djrbOtb6JugEi9qtwyAz1ndluifitYieNb+5CAVbUXCVs36C69EVITOd/QGzx8bf+AiBNtLYtw
98QVrxw5VlEQT7PNTrwrEfKUs0UykGr/4mpPkZ4gHDvBQSSwmBvAHXY/4UTjEBSJmq+SRZFjQQfG
gFZopRsoxoTx79EoT5LSrS2Xa7bra+VAbzFa2dL5NuO4NAD+aaBRElEkHzJzzmyXanynOZlJR7ud
Bj3s8zn1DqTDyEHbOa8DJhQApeAGEtliQeKbIjZoflhjJAYa8AIraPOVyc9sYfxuFkjqsH9aIOou
3f875ZksdSb5h2YsMO9fiqhQUv4/BT0TW3e9FmJb0JuLy1ipJYxQIm0jKlhRM9dLHw1AYATfNQH9
E9ya4hFtVwB+OYbrZfQHdYikjAiIn/VXq5iiAfoC0eajKNtTQ7GF3KD0BopF01iyaIBgcl/f3NYR
TNh4i3OUh8CGi7AEmHFclFPGtJNYaHJuoP5BJxX1OygiLREdsv3l5s2SAhB3+wRYlpI/yJIXzFXu
4Y/UOgGpTJfDI5pmqV62twmrViwhCJpR/wcPWVqAAM64UQwI273076GP7dCffkLGciuYiZSPG5co
bs2c6JfPJ0iXFpwS8Mjo4MzuARL8DncXnH0fVw64LLz/5YNzCYZ6KOJb7oOjYJ94ocuoaH3s/cGr
ToY4rEulxnsW8+nn1BoOXm+rhK7Uv8v7FDu6KKtx6MgN0Bhnkw7kUOOZBWwh0tyFwBqbsEFpqBUz
judx+xKLy6KgR6Ku6uEFVgySYEuF/XIaqpizRF4ESuF9aQfpMwGnGbaRF3+Ke/XVk2oYsG0V19cu
Um2NGPE7Es0wAYgdMyQPDpDNLgKWmJZJyA/zepvdO3I435zEV1qkptEmG9a14ks4aREvzMrWdLhj
WOmNFmtbgBqdDLMVSZ3v4x8HphM1NzbujBe2x810lod3SX1dcSCOMtgqz49WPiR8swzNGk5AKXfQ
3/SgMbVb5MFvKxHrixLpe6oB0fMvOMBbCdhMhbgk6sdpyrsAqfBOkVd1vqCoEx8SqLNO4Z7C8i1t
ZHHkBSqlckar4cTxhUrhk57qFipDybQx+BIYQ+NsOBuZ08xPrGu5KAKaKytsGv26F+GemyJZIYm9
/E4SNq68s+yqEHdeqsJptB9RYv1XZHXdu8tQT3rsWZGRyqnfEIaj1Fg/iI98j+NouYxFL7hDEyoJ
Jjqgn5SjIaaEkiB3+iqlUOcRXYgBzmBTYz4d+skLSZ8J2cneebB56iQDS4e0Fyq3Gr+Yd7O8Sxrb
1/NDvDMOi8RdAhiiVHiSslXobFMO1aBl8p2TkUceti6dHzTgu5lcH49vbiE1xgMdADjW9FjjPfug
QhGOk6Iy3VWYnu5ylNfsf1WPeA9e0Hv34x5MdzaQVHg0Pgrdx2ZKW5jp+SjY7AWSinID4OJj/iWO
s9jYMnWSvCwaIv2OT/HBshndLnQoiX9BA8eVi38+FeTKsmZF+idTgt9lqX2dXJaPG557UJm9zRXm
ogyMz/pPo6CdfDcnltuDW2+5ikslLizZim+LNuMp7FUP/fp8ck+w7ybBhbiruX+VmLn2h9mI37S/
0MjhmFsE6YVzOVGCCmb+ULv9sSwO0J9ndzq4GZ6tukPQMdKlbbkzmUalGqmHTCXxOV30+Ln3Sm7A
SdrxEvdPBMQygTbcrrRQ5yyuChc5TG5MKq6lPRVEmk1hGsEXrXrbEpY21pXfJiyinURhJDdCp9FY
zW5+OaKVHeBpc0YfG2bSU+370B59GXDQeLFEQ4I7tkxjcxgPQvLEc2Qce4+sHpXSsPeWTI4EjhfI
LO87eeEtNy9BUOcPuLG2aZVrdWp6evAaLeCQ5gRZUXg9eLuym3luRxPU9zJuF+8wi2INZXviGv8Y
C270N7TIHTQn8W4f+TjMr7kC+WXkWyVBo2CgMfkwUku2VeBeMD9cBtT7cWdXUMulsZw++Ks9FO8+
nb86BtOEYloP6Jb74ZlZ/yQssKm9gfFd4f5+tKSrgPntBc18SxMuy3g690yTB8W81U9NOJhOXhr4
0lAzIRjD1rEgukP/L09JmdYWKkYKRCmvfG+IHsA7j9EUqRLRGnpC8baWzCTWCUNRW4Fr2K7vZs1H
hEWVD/nNHZvbCl6z7LlCC0ZFR3ZnfEBd2v+BxKgdurN2JnhXfqk68xonZq3HCKxiEDaABMhTv/LU
H3VJTthuTtwG4WxPiyWNA87ShYAqhrGb6X7EGEA1FRYCxDnlEHwZCIkKfRxq3su+vnCZ2JBuCZke
UsFyZK7muxSKg6jRV4EMzU6eexDn7Ze8ENJHJn8sbX4OZBwka5/Rccv24Gl7MXVFwtmoi2ujJOs4
aQlyW4qE+9Ucn/9sdKdvC+5f+m/puUxBCPhbwk79TSCBRo6pRkbGlbt3NYdXAbge9xKvUsC9SAhj
NJuWoIL3ua5ERW54eTT9qxKgH5hLjkNT8uM6DkiXCubgSKo49a41OoEnynJxuan19tL19YtjKMZo
XAccaYQKyH4WxBgPt5n2SLRD2q5cE1qTqREH5pW6g7kJhyZHKF17tGJqhpuH0j2Dxz5dszNT8qMw
XIY3ufvy5Bhgq7g8jScViCTB4siXdHGYinOgNBxmwBB+MlgI11e58oGTlIppb1tp753wIOiTzY4I
JucvNrmiurp8PrsJCIQO3fvZMqt4Ynjh7L+a0Tmna0XI8jVIkJWLD04QTzSqu5lBJqpHqzAZBpO5
bmwaFFSN4oNYaZLwzZQ3vewn6jLmkez5wFeGk92IbgJ52uJTaN1MtywRbYS5Qp7UQJxuIZHQDfAI
KYQrWh5LPdU3z+7SCYl2UeOCIo4PRU+1pIFdaFoATkqf029lPF5xOjlzZ2dkqnNPpIe+QuiWavCd
KK0od7BrbxPCVdDZcDbCnwCepwJtNDmx1r88z10hCpHjLfl39R2174Jc++4bMXnETVvW+GKqz2cW
tXfg70ttMJJ4YMMhhgICiQGY2Ro0eM/EdtWJhkUe+dTaM2TBeJDazliKnf6v05CfxC1UCYzfxqO0
sJxU5P1PpCxiW1TgFpSEfwVbA168AiZRmz2Dn+JG7J4qcg/BwcgO1QrovDi5g/q0X7HJDIw4xvX6
24e8KBiiz7Z7b951jm3Pmcmja7NK77+08e/930M8nuE06XLi55uGBuNHe7EntlSfyEjFJLq76Ggg
WKt2pbROxftVuEwcCTsqTC85FRQdMC1Y/dXc6PB4VGI5Y+I1HoFkqzjHYslCiq1cX75nRev86vm/
NQymLT6pWg0BWcHykGGwSMH1sctVzjZ35RFkLHTPtNMnngJuP8XsFE4w5hYIVRTZUApRN8bLcnSl
+QOmOqqi34ZgPjFHriWKbq5bKYymUudMvDggfuj4Qj4OAO0MjJrZoRwUb7ym4yNR/yJFXGojZb60
PfNhVR22yzQT6AkvsJea+f8wuU6PqfAiJyzYsueVujd6h/JRcbYwR1h+l/THOElitjJy7uPDEg/s
6+EwdnBBRykCDSzurYSevOkWCZyX3ZWFuKKrm4b3WfoefdCHn/T47UbCwXK6gMZdTLx7eQWkVWUe
3aslD/bCaS6/M3WmT4pNTAvv5GlnqgHJXRhEIUpMBdcatOI+3Y3rhWbxyGmTcSAC5enrXr8EajYN
NnaOpTK2JN5WAkkuhUeRwoE558M5zWW4Ub9AqxdRb6LaIZ22OfgyEesNwCBbzbjtAoJCYTmi+Bfq
ss/lbw58CYTL8UMGBo8NlvaZeS+A8dUrUcudLIwzX774lkzc4hodQb1tgoxdiBQ/A9nuUQw8YSez
DF3ZYDEBHllooHeWQF8sFOj4hAMwRDGMe0XePTyKLsnazSRRNFgb5kvali0jBnhK3jxIgk1E966U
w34alL/rmqu6vWcHZ/ehg8woUQbII36Bw6eoA47sB/Hl1nio8hiOD/tI6Eu6Zol68VMsu/Z8+Mir
2CF6Ktu0Q6VtiFahvKD3VAHeyabB6nN+vnSj4vmIvLH2IFpY0xBsoExhGj9ty0c5MNPTB9BZx1It
tcAIxBlVJR74ZConTlANEtz2+Y5IxT+mCykRl5VGCAGFU1FG44EOPXspf9Ki4l8THS8a1tzVbfx2
pMOKfqsDtKmnJkQ3QAmU49UVvLimGqEm7J808ydb8VLYP11kaxKEGdrhll8AthF5ZX4oImbpbjAb
vWQ3jqCb5ifn9wPkqfq2/2FIbQvRdwpx5ghKfQTm0pxN0eB0FPSC7aUha/tmxKWoBsPF1MRjLjvJ
7thLjZYZp1ykZea+pic+G63UXqeTFoXhwHl+v5H0oKTEkV1wP7OAWAN0rCr9B5spHbemL9K+TNNy
gZYee/ELQjOMvFiAowCo61xHBevFT3aXVKQUVWHrKGTdVGkpPwAvdFl/8duFPy727r0bXYmRKvgM
kdO6/P8zX/4c//oZRH0kLpiWIH10ybB3lqWBjfnKMUZw1/2nbG3eRsJf0CiljBQBIGB3OSMrTYTr
xq8BgawxZod8dBx5NaDBVpTm9V/dUAjM/obUHSb76GzRY1YykdbUh8Kz+/B3u6Oj+BfjbdSJH0gv
RTrJJYV2350zrViDEKxfLUU8YA75fbGphkzl0ZUNZi8dyIhD8k0ePRTO/l7/mWeR0XlX9rUV0EgQ
jSfr2nBTRmi0kwJDsp6Y0paYaZgaHozVM6eW2SbUpeGTpT4KZrXvYoF5QIUTmNOOkWZJ3G4cl1TV
+zqXFSRDmq3qc7bOBG9QUONFvWt7LKI1skYj8WMKckMWPbqehm1PcOsnKa7bLLrvJNfbN5umPmxR
778rxXI4Rxo+DLNjnYtR2Q0akbt0l2lrA2+63xqi58aAHx+LtURfko3UfJPvEoU9wMviJmmTvOlu
x9EKYALpwMdrEbtiRCLfpxVd7QxInLoAPhzZYglCLvJpxxiQBhDXe6W1p4TZH8v78Wp4QnN+LkiZ
AeA7Dbs+mq8pY2CDe3SAqSQG7YCUfqq3kjRvcPqTNcD4JnIEjngxd8DYx0oebgsD5ZAvOSAqAOgE
m5c8JiIoO4pxlZfL+47qMxYaApQMxza264LYxcwE5C0BFaxkTSaUgw0TM3TDNBYSQ8BIHtLH0fAT
jIvanRSvAkiSAfJZ80PFQPZmd9YWHM4wMKlPhI4bBbN2GmYdbQ+/dd9h4QfKfLUyawlMlcvUuAgR
QB5NYDN9Q0Ub25CWNJ1qEFvyFUJ4TMjgSi9mgvnI8qmIeR59W4qb+uJaZzs6SF0f37RCQbbCAnWQ
zFmG7ppp1AWH29GPa488YFGDcIriqWa5d6OMgcTSOMlPmc6/deDrDe6+T0wRTfL75ooq1oGrrp39
GZs/L4PTG7rgpMsrLXPSYVAi4nasURKAE7RsLwfEZxwNrcTjnHNlTTRKjZSEDsbSPiH3xOrqPXbQ
W1bgygcE0fl+5FBPdeL0Q7MxqKg/ayFZYhQaNEm6rVqrTe1XRYLwuF8X6lyvUAIxjeieKKUPDTXD
jKvkpCUb1KMU3ja3FJ/lxl+OIHx4LavL1x42feygHELZxqqbZ9dvibhTFkXZHsf70kl/UTDf1FqG
r4njfLHgWH0vKxlrDOo4nBFxiatJS5DN6y3+kDzGXsNzyiEQO5jh5cP5jl3ug/ks3OwshtuLjUrv
mKohDJaIIKunXNU9xU7O2y3qyuled3aShDwq7ExfVyqIk+EWKmqpA0n2alnZAbIlBcZnBx2Wq1Q/
3IPUcyh0r78CewPMbcgKqnpatzlIprbAkZFD4iY9e9/GBLohOdrbCrkpFHRAoZLjhHeNaTYdoOpz
6iARbB7ARizvn1omWLbIphQfq/hcLKkMZrIRNe7YKI9hbFUIeEPDlod+JCZP2g3d1cPjnqIXf2Ms
/6rsQtz83LfTWhaf6NiW7x7BEmPtftvU2ejXnCebHxbLn7PKZtbBMgloNQBV9RtDUsjKFoeHOFwZ
neE4TeKUhc6gpARiMf+nw3nPNRWl/Q6uHsioLQFfQ2Bk1YNAeVtO8JLcN0F2Vm6jiFeJYGWGV/A+
LfZgvAOn9uXS55P8PHqPHOsHZKtZKZFO7x6mFaz7lngY4+NTQ5gx1kyzRu2MAqCBE+L4APjKOrg8
mMOGFbznadgTn32KIuBPX8gGWZHE0Qj0PHjlXKZCzO0VMeyMnMFHhrg388tEVEe4ibtP/tP95NLm
WbeGql2TeX3XTNsZtkWx1EdkykrxIiczhgY+SjPcx4O368J6n/axGHDVtoBYrRhfae/bA53HZuEw
+vb5Swo9pltjiHDPFYvFhqdpILUbajGXoWMJmWPAyzyuDUC6z3j8Fb8m3r9X0ljD8zPO/YzeUmWy
JE8q2oA81FzSMomNe38nqDasw5tYUCz8dBKvkGtWRwSAJfOhy+ZQyJ61CnlVsHOQYnw53MlCZFrs
5n/auNk6B3oVsWxvif4Fxi/n8g7RAlzZ+cTldaTVDJzGoqUmP39H0RujRtbZoEX68oI9yqkGq9w0
6O8YdUE1UnRla76DEFHhhobY7/LfYI9Xe459j6EefukwHfNIR76UPphf4cNt/jEgU2UvK4T3fr/x
feHIsXA5OFGiAccXPF8+LXEnPRh7teVQTr29qX2VF/Rgli60NLEBtzfJlFTt+7n38nUL3VDAHW6Z
yFK4j5zr3R3G2G0bEuyYQANd9XSOAtVS1X5LenCaMxSOMHUfkLT3hLcEClcFnYVqoH88zvkQ4HJx
GfUGHztnuMyszR7UPyOY/xUj+h2vul+9TXdL/v6fZqzkOf6uRCOPLkOn8Jbei5GqtWmwOSIzQSbJ
p6kVl4PDV6bwdAut3THgc+bCShTufnoPEfXfYtbcsivX80dXD03Wyhgo2rHOTewhs5SbODeP161c
hhMHemjkWJveBxRA+cFL6HPiM+JfCkzb6OlPUWCaoD4uGSDmEGjGb/4ozur6j9i7S0RKRReczFKI
ybLp+u8bkCfwR+a8XxDZ+Y70QwuDQRf9x4+AOCl1jc7zFlsLiaRCfrwA87WwCNHEil92e2TCjRBT
9DDUKbGHMzRAbRLp6/fh3Qm1hKW4qNmhuNjG5M2FC054tK0F/G3+FeEqM0yVlpQzc0ZmISBQjfWD
K+YbOgoGT/IssbVq1YDNchyRKO4bYaMR8RfsrhJdfoBAsGlGa7LFwjHQ5eAHnnbBG9/Q1ZMEkNQ4
N8jiXNntt0RkKoNmJj3xwiwSjAOk1B9LwOaDGH0uvCmG05EzWHt8YNMZ7pIeIwTSrp/ZhuZi8WWe
oMAckpJhrD8ctdXD0x2eWCayZ0VbQ2ka70J7gy5FpfBVj7EcWphagFj9pRYfYacDYP+R33oa4xpb
cgY4bFzLyrD5euhP0bC6wG6ygxzEbahbVixnm4uBpUca8fowPlZ2cZCjDzp9Dv8x+3AMjFsP+kV4
tRJsJRG6tUY+00Y2LdMyoOzr0TZwUpP+bG8jrqowlE7Zv0C2/TuqZNF6zl3AamHmsJ/4wNO/Atrv
tWKRxz/GGqjMcvofiVFqQO0srA+ydn63RIndrZvFe7CVK9fD9Z38TyYr21db7iSdbQmG++VqM91D
5xCeQcF0wFPjwQkvuRDaTwPUzwBvh0FfoIm2FOxJTT28ZKNzsukz5HFtlakn251y8W7ZcENCLg+F
rHxnIdloH7FEshO90f4EMOVVqGeMqdFp1qINDvUjhnU9BPkizlSeEZExe4YrBJUFQPezAXwwxBuV
c+ePfUfIeSYuOXXS0I6IV981Yb3AlPCJGoA9c82rP9kyRvgQe1aP+Zx62iNKjRchPHns99xKYFu1
mz4m4z0XTwkiNGvz+Nh1JwEv8b0zDS53X52RPCCvJAjftJDIqdLbPfXQ8VUrJewJjjODnjFYPA0W
fAAQzVlVu8o5wBpxAiRVYSO6IhzhAX2shGhU0wz+ml2z67s4WlXfXUFUDOxzim3jWJwwbA6jVp3s
Vp2OxBQdkzl0jW0FkVdLcXjK78lIIVM6w1w7eKtagzr6s/DTuEFcHrPPybotu/Usaw/HM7bbgot0
lEeJxR1x8oh8z6rlkDco/eUY+0EhLs5w8MaljXLdmCw14OG0jHNSaR4PkNievEBegUp7fuKuWm1w
dBwvPe6b7ez7g2H8PvFIgu8AVmV/VL8MFdtmGjV7YqVcrOXcUoSXml7ix5qJPkLCV2L6s6ir7bfD
cholmotUHrjwfuOhvNf1BPCW2rwD00D4jYhSt+EAaSpEwrV38SuT4e3f0kzuchBUOoMnMo15BSrn
JYURDBqCL0SU9kh2jAhdVrdzNCsQ9fJDcIgLSvlxD5aimXW0Y806W3SW/Z5kv1QHgUN8eZKiyqPw
DvmGpgh9jGHxkQTWrOT06EHWZ/6yZ9xhb+Lc6uxsZeo94SHvgsiUsGj+UPjkCYyKqcbJFcVhXSHj
9feKxws3qW4keshIL6b8irfdpexbA+1O23FYw9RCHEiwws454YoZeLoGF5gl229Yb743ZWgb2Mb+
z/HwC703jFQa0Niib6stIUCiiL4xbHVOORk6XSEuD1ZglJTXNpb4D/fP3oK00HbCms1B3u9NyekF
hBMMrFLci7mFkzP0SG/i50RXBk6kwo6qOaGlA6osJD4R6IgTB5JLKlrL/nzEzU6Pl2/aPVAbkWbP
UBsBkVEMXkqMGQbDhU8R67LrBQI6Wo5R7S5bwDZg/VUROIlwA3pUkdy6llDgIXkOo8DMEmrNhtBG
2u66t/wKyjGFd54d0/oe4KI4LvPRRafsuM7YMbqcQfvTrg6j0qP6+fGoQuA2PsTiAhpAuf2shCKi
z87G86JAz3chGLRAfe5+zY2xBhr1SjRa2QR4Q/RVWR8EW3E7jJCLWZkXykQ9kx/EwvqXd8gt/ad/
ATY7pXNQmiZxxQ5M73CtMzFeO0Gnh1znhhSPlFyyVrUdjJl6glDydQC77vmDm26ZRF39Z1hZp8Bo
Deab23Q86jStgM/y/AsLKhPbaTpcvJKFIwv1KDUaT7yzLv0lg+bvozoOHUfQl3LRfUMDGuWxsOO8
/HDd7gTGy+JeUw6z70bw2Gvq4eDKlnCwWC4Hr5SXMqP8DZ6SiMjAXtUbN2V5RGBZE1kftSe9Jlb/
xzSfkKW72DgdukrtoXUuwRONBUeYAQMXDMw092l3QPXFiu/JgW/qE6zCObJdLlwqk3RTIi/0mO2u
DbMfzAsBYQbo3j/a/RDJL3yH4WG0m9hJONzZbxvPKK98/Uefneoi11FXVnqRiE4VEa1UNJfuk88p
G0XYSGW7T4UG7LzD76mD5pHbudbsWeYnYugZKO0fTvA6jFykUq9+nBW3ylg1D2S55gc042hlrCkn
61FWwJ+8w//YxdLsb/UDz1SJLWfwrBY3KkA19xtje2nUdL3lXR8PawaYg6OVJMu1OM+wivR4QgwF
9Hzjqqd+ojxtYvkLw+u1jthYEx5hh9BBot10bNtJ46xJ45bS87wL92LmRAOMUkVc2c8CxgrXAogx
GTZ1b85nuwga9F+0uVIRD2tVHOSEFaYexTGv2dWOphcnPeCHB2MB3lbfKKou55ADpmHDFRKZ65gb
Y3XbqKiR7PCYnvAFbujVjN5YzFXLqKhiZFgDiz+0U6zSm6XhCr65/mFhJyNcPPAuVlh46dSlpADe
vrs7SWz+v/JUDE7kkzJSc6gPAPOYewgIJYbFZ9g4S7h9sJNVj99mFbR1AQwn3nFBjdqHA0I95EKU
BNv5U8vZG7hubhvYGtEfSh3PjTwIgRnnVT27rietRmIJFKpoS6mdt3Hq/nn5kZtBHrl4JWiQGmcM
yIQT9HOHVVDaLzjVX+yRyRdVag6CJE36cJWhAVRbT/DqWK6ONnbnNxDqqAvbRhxXbR6/racFdPC/
zAk7VB7iE8loEbAYbzf1OKYQhXWAyBNR68fxLm6QraD3/Ilo62mrEiYgbvyreYWGMjDfefEhLgZx
r+61Hrper4Ow745hr3LmNAy/mqJdmDaar9nEzU0o60SLqo+m1SHQnFVjy5fbMZCjh4YVmNJ1hDEq
f6dfpos2xnmyKfh7i+8hol8xB6p8eslEiTfFwkS2dHNiD2ZnI6REG0UFiOp4t2mBBqyV7/mbHu86
GhQXHP8krA8SSzTE4EyDb9sfpCJSBX1JXB9dUs6wo+5H0ANBNXwl5Zr8eEgAhDCs2o8FbiXyWSn6
6imtyICHsjmrhUiwBKFAuFoFh5nnN82rMbWSLdtXiJjaipCs1e6wsg83Nc1EFl2Z2O38zR9z/9U6
GSDu9AsRwfyxNvd2QFhmbYS0LctVD0zKdHwnksHJ+4ITTENIvdk9wX6OxuQuHnL/Su4AiuxgtnZe
JSkzoi618UumyL91+GXodmm0E34ggc8M4591hL0kxilBgiwrKlYQi342B8tW6L2x2RRlfNT4RWSr
I/Q96wwrumeVEv9UcBs7iCi1PV/WRSlfmG5/LOjuGQWFVPUep0Bk+m9huEeQZ/ikf9zQBnAz3eWs
xcQN707cIW0CArfD3Lr/TIeVQdCxFrCrNdmDqk52L0681PsiEoxh5oPfiPG4MdY/YMHK1Q/m2MA2
W9s+w7aiqFvRV0FlReWReIq04iLBEOdChQ8bTDhjkNRg4xmJXYU0MtHlSF71rvN/HPBinvdPAha3
SyeHxDr1xvUpAli/P7vKYVmJ7jNGvKRWy+CBdlVz/WDkrB32EmrzU+LhGtqeVlZxofrS0wKg3c9Q
Dcvxuot5aochBtGxtqUVlyTLWnahqfSSeIT/RqttqrMjfxz4q2Zd9jDgamtJi6xEd9wLV0Lt3jbx
kDE3vVDmmljCHxLtrYgHdFgDFoZtV4ARX1DiYgKp6DnIjrUEtciMF7xPxBKQc7HqppLnhKrgjA2P
HiXJtLzvtGfJAsHUR7RvHJkuVg9NnLlUeir+AMi9Lkgdu8lPCXHewUfE/K2gK2NnG6j28kMN1c8u
3nwDs8VqeK9gQeE26W9cMN12/qdKPEkaNdwlTZ9Av6J09WnVBMbC9DcgqM6kke0GW1Qu4WXtBK1V
rrMcSt1WGT03J95DTtOoXIiln/io5x0h0FWT3BCBKNWGKkfejvF30jM8QS0uhX/MLgwzHajOx03+
goSUD/bsSA+1+OINftikRJH0yHVDbYmQrlFHQE3jf4W2GWw4z+jLIFw0rggPTkTNQoFKTpNCiSq+
mPDEhDhSXM+oXheXramTT1oJI/MyZrMFQuhkjb1B2dUy1rN/4e36LGZZUSemrpJ67NT6YcqcdHk0
7XO+cw7GOTPkKBW9WlMNYYyKt5ao6+crhWWUhOAtQib92aM55bRewgbqqCyF+u/uyHCswxvIbVr0
t4hNYPrzrp6utv4DXJoeBC2Nu0uGRpu834mTQp2x1iEtEgwvJkU8m5fXSLbBfX0a4jfsCBr5Wq4c
CT4g/YGWb4fB9OxumZHMlvFUmqsZNMMD7wgrqc59p5hDLW9lyks5xQEYFpvSPle1kRlrnswegU6C
HUTqF9FpxRnl1e8wgURplGzy9Xu+SSqENhJ2ILXyS/xaZJoMURzGZkexRwgkGxAB3AkvpMzkD18c
lBFHBWYIZhELZRxXwFdGev3cZQIXDhbwDsHxrYV3x0KDqR37RemQZSVsU+WTTtaSgSh477ku7kXC
yh3lgBcFbxMAkR2iii7cD++dMY07TBFrtITJtKDAz0wjkQZlCzm3GW+IpK1K024Sxjz7+ggyU8Sl
7uBllaUDw1OglN9xp07JiGGl9y/KS/cXdIIpHm+DVJKN3xjwXGYr02L68IK/AwP4GDQZ3ZAsANwC
TI19ONaL4Kvu5azp7HKs0WhJja6reFPPqCvczq4OiaicuWmnQpdXUyMeigeEfVhCF9yZt70Sd9Dr
khD99It+NW+5cA8Qy1KcYettAfP2X0g0M9/9rAw0ZTHAtNbrNq+KHmYpObm19qOCRNBaAmgH4ccK
oCj85gqLX6SWLo2tzZuC5u1frVLen8jTqBJuNB5UDGdcpAD2GgijEgHktD3fn295pm0KcN/OVAO9
ocOcJofLmV5wK/jrcGxZZZJczHKc9t1BvGmE9cGFlVRFBZHXTm9lN5uHLveRhdaOAotE/62j9kQn
YuEfylRMTY72TN0GJtC09jZW+LpZrKK9S3XvdpaYnU1h04Cx7CjLeWXDNRcIX/+ebKrpUBz/isYx
pkOxkuWJ2OnyMdFIcLF+1mGg4HsU/sxUkjR+BmayLfkqswkcuN7EgRCwaThCsK5zn6oPPY99X220
+KbNHswmy5+GuHFpgUiCeSAbUwOGUeSeYHRWyZe4DMbEr1MHMDzdnzI+aU7LMmSzwE5jwqJXUhcA
ascBc1ecFrryjj+xkeJZz65iciRD7h7AGAfmz5bDQJYknvH10jUuprLd1KnU+Zg1uqHP7JaKJavp
JSB1CFv/EtWtv9ggiIublzhwn7WcvxOPmHmSxeVdnHA6I1cDI2Pk6QqcE8SmKqzJ+WOYABANpUV6
DsX6jhQNk2stTglQjqxgUVHdxOTBoyfvNMGfgARghRysJV/8IyogXrbPyKxp3pG/aVy+oLfFKywZ
r8wvVH6jIqEk5CC0igDK/JBrk5mAwO4FywiVFIdyz48rN5ngUl7syRzAUW3FgfA8uC4SzCkzFLSP
Gaiut8yWrvJpbWxnaxev0Io5VRhZwp8CwvDlNEb4FF8MEtZRR9RSyV6WLVXTDeOHU62mNiRcamK/
Gzum8v6JDSZZQGUBq31GER4XbgY33xJXU++a2svencx0IeO4x5Lg7CKS1JlkCIvPnATJLqewuyJx
96mSUJ6djqiQ7kZpczOZe5+PSFKXbDpRN3zunrjJgV8PUB1/xh1LU6yZE2SijTrrvwsiDYqQntGH
x5AS7icKOBKxuUPxQA2xoMnSNPrgC5kfkOuLmnWRdhWSu4ZrUvwkNBZ+JaLIZas5/WSs4H1mOgAD
2Eyt3YiRoMzBCcO8oKyFQelU/VTnL0v07RdknPNZ5B+SUQP8Na6vNHN7hgMY8K6FbOVhLK1MQ8RP
ob+4ZvwCVZJQE+4Mj5kPdb82MjtM+19NNTK2Zduh1HO0snUHi+mUtJdX0ckBTAOxMr8/TXoNxs2p
t8sftel4PCpfix21qa9Il7P86+hO8+5ZHbqw2Ct7zqTGh88kX97Bq1ReWIp0x7wOLjKMRjtNW0Wg
zp4M+03p0DNCkuMml9AsJYuhbtMxxnJwXHUd49aLYeOXBL46g/a8pHJLVxAojqAmlZdK1whnW24H
XfzYfUNloXu4VqSkSNs+hA11q4bAZ24CN+v8N1RrrWQRGQXS/nWLbFLEOilQ8E3ok7SS+tVcMx8f
BBXUHpFhdbBnQNiB8N7trL+yii3Cd+BrxgV2MFndKTJeuGuPuuV0D1lD+gcY745hi9TrMLxPUMJ/
eFWqgS/T6RG1lEfTz034wbaXQqEakUH83D7qePYB/akm2Po8AfqH8rt6KQpl7AK1xT1nosSKN+ZI
EhGWDDky6ASEsfH6x6DcDcuv/pvtW7d/sESHzW1bcqR1TEo+l/+Ixq+SxPTe/mj/aG3ueZstwop/
Q54eihjLBD+xw0Y9F6HYRujfv6yt7doWpJ0qmUlNFb6xlyLPTidzcygW7HU8QbaSn+YtgtMAP8lr
WHgQjoZ/9+faw0eWl8NJLPsXQ9IEMv4Je3dFQyRhsxwl7mEfz9hp2aoyyKF/KTMutMiiNYgu5tP0
HBJJ/8GBV1wAuxRzP6ixoKUC9rfKcIqj/8qy9aEbKSKeaqXPpBYdRGlto3iWSxeqe80W5BuNUcqj
yTSBEMpwCE6tXVnarP8E1ZzeKqYCttsswNWsmrOqo5rYWvoh7srMdG4PJO5RlE1kreN9Yb/9gxWi
qca25pj/F5fvEnBRzn/Bn8XiaewQ2ikDVVowzC0PvJfUP/bIRnAowlHv1WPh4Amvup+0QY5Yb4cJ
PF8iRkYixRgkTsB5XwobBrDJGpRITwPW5GLN5npb9CPO0OZgGxJFUCyoWVLXeCieUHh9rXx2mpkw
wOUcK0u8Z0LXUU/HRtv64nKKUMzjJlZFS3kTubJ4G4pA3J3W7JBmtd0j64F23CfHmrEXwYyHTTGM
OxkNVnNq78E6IcN8y5uBLnO6n3YEk4kLDYHtQ7w+iMRkO6ttM5GyUm9WBR8Z+XE3pv6pSflqYEeN
JveWgVtp3JkcjDt0CHwlTcW35osVo22LeIwNvoH+KaIr1eDNE/JMiXedcsjhjCoGM/SJTPy3K5m3
9ePLymlwdKF3v/3J5JxyPkXWrW3cEcTDQHDV8usiklin2VqGMpTt1VranHB8+PYgAN7nSF+u+s+l
Fs+RajUZE/+VSetHNxz9xkSUqrNV8pOh+d1W2/JEuXqgTohtxDe7nEUp8IXscHPz4orTLzwi5I1h
6A3E0bTwlGQJcQeNYQq62DCb1Xzf+C9eF9KD93mzsLurB/zIhDUz3xYZ2gmXulye7fL9NmQE0yTj
l5d5VwcyVRM5PFWbZ7vDAtguAU/5M4+68wzGWnx6bDwEMrOdJgZr9uQ7xZcqpgjTpabjzcPraLec
SRvSh4DPZLL57Vl5peWP0VLWnT3XRC7+duHJpHZiMPEiZznpxI3npUS8Lg3Qm9WjUWGNcERQ7VHu
VCqwlo7fUmwehS8OaQNA3SmUQsTn7sdiXZKpSLyGNLcJViiDn8xfPQhQ66cmVHZYKsdXCtqAhLUQ
QS6TKqtwx4axNksUMzGY24Dlm4edJ69IJewcewF1wkcdOMTCRupoKxvGjjznv6y1GxW8kbx4vo9q
rK/XRixaXCXw226DXwKHJk0O6xFX8IqW/QpET4C9BjlA4HqZRxmf2x22+giTVL1Mt2uP7AkUqeXK
jHKL7pq/r9wdz6GeJaF/t0qo1ZHsuwPepXYc7YCM6fUydLzAKQIUR9PHPObU9j6jdJRfSFE/ndbm
k6lqtTfF35/NqqkqJn/3ptVQfc551W2KYNEm0LBDMU1efxPi34Z+aLWlhylaYa9ZR2JsvCE7wcg5
xVIGK6OUlF50K3LgzkbKJOXYQ+ho4nxt8UjGbNvY8940VChRZ7h2RT4m/HY7V+74c7Z4L7b1oFZc
JVaf4fZZoixJLd/VQGGHyax+PMJVlviK2jJV62VjA+AsCKQuXXWJChir43csZRq1hcg9kK5RzkAb
GDb2HFPxjMlGuXfWr7uep2MLK6R7Cut0ZlIlWGgy5HcaVGagUMHuePAdOsIMpJXPCxy0G7L9/Bna
PRanXmofs8zLCadRP2YcBaf2jQxs1StcAhYfeNNYeG9YYUyCW3GVhOAlvhSgRk7DhqSIwjrtMdgr
CQEMSYVwb+97NRnkVRzot4sgFu8d6I3DWEHYjUhrFh9IPnU5gwX/pe2kPICCi5c6SBMrqn+7/uc9
XLXiiF2cPfw6o5PF0BvYDuj7uFEaaiJTJZIBhSrk1AHBGbsFuZIX7HHOBe5BWwT2ji3tKdNhjC3i
WxlT7za9mwvrg/SufLfEjaKtH9muXePPojXcmKUfUJIHgpHjmIsD7llY9y5hzFwZ3BG0RLPLQ1Rx
5FjX90uHYCbNz4aE5uB5lio6zDiO95y9nnL52OmzpDQQoodZosEtREwDN/CPqn3w8xDI4WQ/oFXC
Mx+1+j4nOcOLUS+hIK3mLU4l5VSRhweKa9C9jdYjrQQEEVLgZjhWBqh8b7n4aaavTFKwXWh1EOzx
D+aHm2oFC4cgSASqZITDSpjRejlNMkl8MajlxcwajejlMGZmn19SntcaXttdoVDBCtC1yE3vJR9v
K7m1iBXWD0HfcvJf2OjSmEiQ5tkX61anzYRwR77OEOpdC8yoWtepikVuIIXVCE2dSifRtgDvVD0B
9G7T85fisrA5iAweZxlKgps+rO9U0WypGxgGhGGq6JGNrJ14PpkFgm4AfjtGotmQKBDza7CDlGLM
eTvAzsuvae5axGPid9MYkodx/YDChzAxyGSMCWmaFrrWuMu4ZYiNqAN981S/p+UOve7KSu4c5TM2
cOCdRto4vFiMbJlR/aIDOazi2wAs85PnFiZ3JtD2SQRxrrh9CN4/aY3mYzksYtu/uhOFc66VpKbb
pstKOJvbo1k6ynWIEdHohXY1CI+4h4HGaEAb/Yb0fROqltbMSXDop2SZPWR48Bzg6a7UmxD0Jm2/
ujhRm7JG+VsgfBK6kH86kyWCTPWgygwEn3ewDbweKopm5cQw48Jw4BLuzKyzWU0OdRRqD3qQmHbx
fVzDTuYsV2XVDqb2vctlbaRCVFnypa0ojPWOCS2bqYjPO+1YhgL1KIArsPry/iIpJnFgOX4p/URp
F066dtRRpjwqD11sVlYwQlbi4vuFGouFUFBDbMxaZEBRsT0UJ2j8A1BR3niZxt3Kk3au99pjNVlo
94hbnnSECwd3hgMU+KAfztff+Q/zhCpt6x8CPhmP9Ks1ZB0EU6vApeVEqqlGArYl7dFOLQCk6GDJ
DIWLwapyzNzq1jKOTuNOnmEEmEV4ltcNv6fd8MIaK8lJl5KoIWdUJ+6jS8rYGxIg4n8nxhcqzEcx
7xTVSViBryu9Y9E4oYF4xame4+N4ohJgplT8W3/7cXldxIGu82k0zZQb/A/pGTdRS9HAWkY1icox
Pl3Ej7oNWMjpj+aJgKOx+ebIMBW4xOeMgKylBlfqKLR5CLuu2uwy31A9oDBHk0nTsO+DS8u89N+8
NM0fwArxiA5LSy/2O8xFCfC3RHDySjFy7KszZ/3sqrbMPJVrCBwF0ed26bQXkIRs3cVfSKR/ggjn
0CNx0sK3kl/k0VQ7JE0KRz4z9JlLljSb/SCTJwauAbuDIQQwYzGgUsVhOh9TKqrP+7OzkplH38Hn
aZDDmjcwvDAmcG2MPhG84yvln8aUt0Xg4RF3+SOrwTEXCmbqA/q3kUJmRMYHp6b5AWfNb/W9swP8
mJpB/RkEJC3bGPu17LIffU1aI6uKNwUPsbM0lJbU1pSunglOvEas3G+ce1Z3tDlFPXYial/AT3gl
rUpLg5emmR0M7eh3IyJxO467rLIixFKMellU5aoFF7t9evxzPmsQE3fRfwHoZN9YOJOuITKWGicU
24PRwYXvep1LK5xFfhzYNza1/6wWVTXpgyPRMumxPa1/CjCAXewHgMm/vCVud5ojhedGCt0etirG
2SFyMJjEw4G+RIfty1onDwJOygmuA8hVh5ysVYe09FBnEIiNMKNwB4DZpa/XV+If/txIxTMhnUUu
GTGZ6G7/vmVB5INZ2x1ZFtieINhj5bkiqVTNM2ZCnQlVv77Ivd5L65gjBE3Sxa5HPpkZp//D2lOX
Y1fR6M8s1Se5Joo8rsEgWB6SX+KaBISJrgxcvXaUmFxvooOS22w3N9m3osvNB1NiQpF5p9qLYNXf
HLxrGG6HHDFDbDrDcyt70a37T4pfiydEJK/GxugxSH/D7eKZxLR0fhniBOeVN6JKhSs40270QHIz
UzOIeCoj7zbmvIGyzkN2tGI4k24K24fQWM+9RRyg0NKMqAS/Pl3y119hHpYkYn8P+bkeeAQuBskR
8qJWaOrcXaZY70P1aauI/1izEpEWl4tzwHZHSZpVEegkjOm8TPLVuMfLZ5sU8ub1v2BhOKDcjJ4b
lGshz1PjgarQoAFL6F9W9AwcotjFcYGcrcdN5MrZbR+DPlSxryzrIEW8QgnViWrtXn14JKqdgy6A
3cduVOVfUuPHIHY/cSQ0WuHOfYysigalLuUmq/8cBR0m3dgU972aLiNC35XaHz6YSs1fHlMaWb7a
mwGOYp8xqcsEcz+lr4X++0tEpCrn2hLq3HHVsmNrVdKgbfTTpwKndbo1MhfaDtkhBDvGXcJHoUlm
9RN59i/ZkxPVW+i2q7qAD5baXYczjUAlkBuKh6pG4vKuf+uznOvZTMItJyfnqwxZGvvAq+Ffxjno
xQCt4HH/NvkrG9F7mBDHLjgRnTGxM2jyJ3LFXMblljr3NL4IOngXXucNIp2Xh3UQx7Hkm6Yxo4Uc
Xlrcc7X+g5clOD6rMTUVYU0tTYIA4ldi0gCLaxOwWLLuZhlHugSy01Vb/xZ2CNWB4PmB98RawEd0
+4ZsB7M70Q8J5rdiMHB0SL2rP5ivayVoX4KOvfalt5akMhTkV3XpsMVYG/y0C89CgYEWdaXDIV8u
lfBvHNBnqFPHZBHjFfBd25aDKVd1Kz+Xe6GeZw8mxRMeSUKNUGiyR6A8T81m3/suZSuceJdV8y5G
aeAs3UxuYGRTC65CQnlVCnh56EaXISie9MmO3CRxMiJTD/dqM2lfzt70GayoK7ye9YwV/dIYHx01
6AOridkdvAGgN56e5sGhNBFi5h3NxsPvgMl1s2vA/FclgemBZBNazuUAyR4Q9eyV70DY2ySvcV8w
//jkCqlbQkaV0DzGYxIGW0UcOBclLFkaM7nLx0Juj/dNU8hRpJ4RzChq6GHBF+CNu0lwXiRFsGo0
EvBZBNzj5jI7hYCiOome7vmz25miyvtYntdPQhJBHbL6NbIRTj+4rlDL5oQVrlbH/Yto+S8XZwVT
B6+8kUrFLp50fuRRUx6U26eRH5B4gWgZEVj+8Mp+c5erfjXLFSVgu7vFJO3a/ibaxOCb1CHmF9a1
wuvzZ18hC/1zWPDU2dkyYFCnt17rkhjEhyQOolgQm2SJSHvjZ+w8zr43aau736K+HB48JHIZNf+N
wVpy5bs+Tfc8VoxL3hGVvn1nu6q/4pz76XvWI7Q+ttmzB2aAqFRPtQQcBPdz1d0v/mSBJctuLxCr
mQRcL3OyCE+WIMND5nz8yZ8WJvKI+Eqt8470NEf5Ul+kbX5NAruQsoNwAMX3olrrvv/+k7nuMfpF
S5N7qazmigRq77yNSdDebUQpz922rtmtChHdoZ1+Z9tmCeNvuY94iFoqCWycYM7sfi7J7oaWchpL
W3PA2tTGlgYuiWUaZVGIw49EN1WVyWtSlAlnPcQ3+7v7DevQj26s7n7wYj3r0jAluDl8NCvzVtLu
/Db6mePCUcI803NTPgdCauFdGDylRnuDP6Nq0ClQfO9ptbfoijbeSJdNRX+yR2w9qjnUI8qs7Z6s
BAi/scfdsPXrUhW1Ad0Ezu3OUNgU51u+ciOI5765SzR5MS6hJc0lvGTXfh+BCiNzXEkwwBByROT3
5BOwOZUPd0mMoNLASg03QJRISkkrQJt41235gjfvagv2OtVdVnhFOnYKVCmw09octqPjbvVNwJDA
9uAx+CWZ1uFCV3II+E20QV8enRw9XrvTycGkcopQkisajgrpG6r9fVFOkYTxKiZNXTSYno2U3w52
1rPRn0Fb8NAdxSbCtkXkhRYNmz5hbmEpswdZOKj/lodoKwcR5HddJ+oKJBFnG0SmyxUGNoo19JaH
1Fk/PliaQjuf99FZUZaR/ZhseccGSbB5RZ2s2L/F/2YI1hEyL5mMfw8NFrYVu4s2N9lzepx46tes
g5p3PueRU+rkExh5knhXp8IX8VQPzWu2WmYXUWZwlkdUBxpPn6MbP4Bgk3SGh3b81Qy1LfoYIJtW
70fIxkkDLw/TmJTI5l9OU2oJIlYhyjB3q4lzUvpDcVMt16W5y3OrSq79/o0F6jMZiiwj2YZimq24
H2qqOwsE149XUfge9BZgA5bd8IPlGPAWrMNM2Za3vFFT2vWWkN9sshxH095oGy3TXmitAFEzUk3k
14a2BOWWqBKokpQhvHDPU+hundwtR6gKIVhrYGJIxbI/XSX8zvp3mdDlHrq1CmdbfLlNwHL5wAzH
Gvy6CMoIUyp51ljOjNCZxhursJYmuli1zzQYrUHA+AjIjU655vASMla6P4xF0Qd2M6R68YuNNggw
pWgDLzIx57OQMTlpK1zp/CfEnPJIfX3riiRdlUcbxTo+DN4BhTLFD98EofCOsmU9LqNRu1X3aFl3
bJF4t6Sp3ccOXOeWnKTXtap/+9OIz4056V5/tfDdYTHqlmlGrBlQ3eejonGPH0IyoSNZkUucrRHH
xhhNZj4W8soi4VpPbvkHyAouEubc1JMvx3Av5+FHVSFSmHHgoV0qsp3nDloCQ31Nw+3mq31n5+jd
F5xBh/hP0IewZvONOkjSuMTxxQFw/zXH/CaaenY4ySqwHGX69lJI1rib9957xOdyWlWjZnbhMHko
wJx5/WCMTjbYubV4w8pGj6yGObVpVEotmpDWqOF8Gyi+r7wpxlm+CmJb3Bo1/gYXZDDSYUotZvj+
JfauXDCk/66XeBN10Wi0jmJLG/XvhI4kLdAw6+gnQdSzo1ausxg3zfHbpdGNMtGgb+Zm/ZpSELSB
9GIRyD8+FcBy7JLlrtcoGxLLI3vuckskG++c6M69YqPx1baVQHGdKLWigD3KORisxJA2j5zcCy/9
tz4qMXvwKE7UGJnJ8Rcd1OznS29+/7dG078oSIWR4O9pZbbrH8Su+/6YgKa6oa5Ayy7tm7I3xTRz
PpX1zDlB7Hb4zQiMQR+swm/XJ/8NLyNl4odmhaPBq3j4YH3FljcjjsXLbB2QFrLqyhReFJZG/ZVp
v1xLdSSJU7471Nafi6EFqExOpLl/N52b/NSvB/u1ktCjjPR9K0WwwojeErY0YerjL7Yvk4CFSVhv
AphDZ0r50Wo8+Rlhgf9WULFxl83xEPvVlp3asTBSI+sVNYziWaTpkeNymmQfDkdp1y3w7MZySuGk
NLcuRNhekGACvTQGC1Sto5lDD3uljzJJqTAthiLrUJTe72iudnbeMCTGqo4NiEAsL6m7S22J32ts
UwEs83C00VdefHv0F1afWzmtNVxlqWqK1yiiJHOsw7sS3ng5qTsMOU8hmGJOLQ0vlAc4xkvp8xu8
f8x1CRfk7IvMcIboFMtY2sPJxyK4FC45zH6G29qKGFN9cangITQKPaZOvlkJ2BuUElFEm81I8ox0
IvD/r4+omLa9Hs+yijjF1PZFkjxp4NDSAQOldgNAAX1b22VYTly34sfoohCrcvSoFZ00gsIc5crM
1BTdZqxmcyLIuGACJihK7rD5005os/Rf8beSW9VGZxFsh836THpyKdk0Hz8bp6HKh2Is2UDTY131
h/NMSfcj58dLBaMDX/qpZUUCcvtsQeXeleOtwc26yYadUTp+M5UR1DPKtGO/IKvptO3H7BTyBH4f
mY9oM9hbQ/W1OY/ysBO7bnTXWXlVQKU5dODWiHfqdATlOscyoklF5OyMgWC2zBLFmBLCboSv86qP
Rq9ZfMAkrAsCw+gXgfhN0ongSGqOBQqoCwDgQ7VrZ25x8R/BzamjlfRuO4kna6sy07b/qh7s70Sn
JOL6ob9JNepOKYFDvESKPEUXyNhwU2+1msLwVseutevJpN4Tmrbv/89iHPKcfKFNV53QwWVmMMYG
nGsdQH5UKL/h0iVyaYAs1WqAS/TYRCidm2syam9F900m5ZcfDJGPDOwM6g9WWjQoK4THPUrPSahW
frwspdXbS/WZgMd7WNP3eZQsY3hbG3qrAATLT8mv/3yStE9TVzXIWtztue1iOEwMqnUNpQ5bMwWY
N4fGRWFzK2AuCjtx415WH/AwhQv4LBI0sYKTkut1LQfAttdScIcFN8iQslU+nrUlibeXsSkyPuJ4
whPb+XyH3+akiBF7NKKOqj5uD0F7QQDMbNsX7wpUfxhpXpSQ26/HmkHLZFJtEmqW6b5Z2LzsF7hU
ZA9nAg0PVliFgwhW5eeoX3COw0QywsPlbOnVCHzIW3QxNNz7tC4CRm2rDSWBNlRYq3Jnmo2V2Gr9
g/L5dlr7AlSgfyv2q6zywpCVxcTFWFWAa0H9n6/NPAd7xdMCihbXyp1n9PzpDEu4X6/fK5GeReLY
JYqXfFSshebJRFxAvALH6EJ8etE6GimlhBHs4GheDCofaOU27f+nPxC+NgITrGgTd6ixbyjtODfW
Ttf3r/voRlIXP2neRSLgXgFbScrmFXlsfW/EuWNzX7nXYNmR16LB1RmMqtQ9WvM9yBuzlS9e0p6c
dMknYsH8AKoBO1rzuZYUMLLmFgG/ZrIj0KLxtVthdLdpZhwlmr956MrqdVJSi3ZWJXutbW9Xx2uH
nOVKNeu5kRP1fNKUkX8/VNTHp4F8A5Jabk85qti4m6UU0Rul1+SqJyhgoKvGbeeGDPry0qatITc5
Ulph1ffPyBxuH9Wm9Z/WNb3xy2jAwgAUMUUGc0coCc2iUJWRuFwG+5RQ5Uyj6IU4wQs7FnxfHCEU
eZqV8l6M4OdXtpApn53s/M3DdBpCpNzNAGDtMUjSHPDeGyVq6qekJ+iXmdzgrrV7t4Hgyn118bAe
yXR3uAlLX6sdsFJh/sUqNfuAg3g85wHmZIQvKdeI5PIsTXrT4ELEm5RrvoTKJNrH7huKQe1QgYFY
fZUggGEv14ydCvrDMVSgoCiat2Df9VC/c/W8rm+r8Sp3jgWBUe93rGCgiGPU/Et+wqzoOINzJ2F9
I1mlvesMc0k4K0atCHSBTJCZq0+tfRlT1bMW+44HT2mTYeeN8JdNrOshN5rBOP1m294peS9ZMSs6
8Vjs1vFKhOlm7bEC8El1ymPOR5kHD9ENFiaqN+CB7iJEt1loY3tBNuE3l9Gb+ZQDchMVdXXYhzZU
6NorrxVrIL6RCwBzpwqMZXqdFHtR7l2ITjxpfBjjzxJclxvY3TuW7h93WeIzHJ4zmudBR8LEHs8E
2zJ/ue+kRBY8gggvLx3RAZKzCidqe6FNyHbFXi0HNoqFxHSHRVAGetXDahKPC0jyXbZB9LTdwZy+
YYE5MQ6mw4RP9tTGGw92gjgRItzQsT5d35Q8ikmqLZ8ZtdzPeBJCFKs/oE6VO3NSZG9WKQ6tgTN8
6xbadrW+DOXQKqQ2zBlxfiRGdCFZ4mNQKq7afqzKTjWn7p/gs4xFD7BBApL6NAAMLT+I97S1zRlT
aB7f2zEtAw9KqEV4VoXeVLy7DQQVyZ53AJHCe+PXDPbVSGRC7sisfSjL8XUaSSTQhtg4K7Wq+Y/U
K/3YKkOqwQC4xRZ6NVgEB4tsQTh9xnRthIDG0j22MkLlNeZCmnRv7Lsfd7aM0GUAcyX/oP5XW5C0
lW7P8rGRlAohyKyk0t98v+Bp7+cIASvR41vAq18Vf6mjMG1bIcyPx6NFKtXG3iPLLz7UuO0btmZQ
G1YUgf7GaW5nC9HONaTbVmu96t32IShxtDnb8FpmJqNQI3pYGtWp7Z56vwwm0AxuuSP3EKnKjHhh
QKCfnl/VaqRp3UOj083ByzeWWhzOH95pyyLYUZUfMZNZk92g5Cn/UVzfnpaVLDg+D/FzlL0pmgAm
Zl4x1eAIZx9whHgh1fhiQZgvMfQGK5Wf/n+IRmkE1P7aMLLAWbB5snjQvOGDBy/JKxaQ9g6F3Pwo
GSZLyFeNZ8Aen3NDVfx0/qpIVfXip2IypfCP9MBDcPbpPoYGlbvbAQVjRLhTIdMnb6KW8arZvwdm
t4aKx47MOQnLRRrP7uHf1gLBIaP0iDdCsD+WQwZXBt0DPYGnMN0jiFCEgcLvaHlwTXqDSL8m4W+N
DluQoVXrciuaYbfJQbEraGtCPWL0J7uN4JwJ5xQZ796H/wLlqt9WD4sFaNJ5qCz2EirhnNd6TTAD
csv3Nlrad8TMW2abqH7vLa48qgIwemeEPdVophs7o5fEiHPRqqOlMh7GmB25pZwWW2VRbFY4tTmr
d7EFS079Zm4NNxvUF8V5B2Th1Z2HAuvAxn4vmX3lSHRS2qeeH66gsgwWLfxVOYaju7bAMf0KDTUV
M095dtyXxpzh9IQSgxqa//QJ78R75/c0nzEGuDlEmcoJwm2ig/7iNU8VBlHMESxDB/u3AQkirk7J
TqFSHjhvVQzXde+F48CkwygTGa2GDezu8+LoMqo107oWHTK9kZeQTX5GZxV5l0ECPM8Lwtvyzr27
1QAKJpcsUoG9CxfCmsUeC4Z7pcD4e2I/73Ye2MjP7cxR/lKqVI0/DZbZTMR73nnBE3knB3dp849O
Ol0C4qHyw0DB5YzZPd43s7QRTtBxJNyTd8t0++Uo3yH54U89uNZ9b5P2sMIJ8QqLKNCnzMW8YRtJ
yoT2mmrm6+wPqhWCJe1BT5bN2RpHsdCExIKGHm3m+x8LO/Nvk2ff7R94rDOeDLHNs9gFNfCs1ikZ
VwGHVkhuL2//osLBQWX6ED8jqOXjnIBMq1xRDnzeUwjhxJrtehPdAjlFrLZMd/JEY3lz3PmkwOzq
Rtia3JFs+saq8b0RklrFaqaX5Eq/AYeqixAfByY7P3YxdQZA8/x047MpIkiW/FNoB1kTx1A0ReA7
xAoHhi16PG+kRR29Ri/nKR1tyQt925LuIzrVKjpkuV+cJ1LvqPAkuvWf7mRvskZuXYMce/vLXXZt
/eY2qhkI6A8XqLo/bG/dA2GnrfMv8rqtyjlhmD8wkiiSjyrsYQ+5N70kBHZbwSgAbXdQdotDLUi9
KF4oVo5p4tlzI7yvUEK+mk+xa7hWiGtWlhIMce9plLB1NtumI1v5dTzLep8FXEughhigVL7ffd46
L8EDu22+ZrrkkDErkhor4aGHiBNX/IkG9cItCkhKYVZkCP797a9xfOlChEjeAMwKtUtcxPtABKQO
lIzZrqOGYROkjq/UdEavbqCmE02ZuRIJelK3Ka0t8OWfxT6Jw7FuMweJvW+Lpb5XxFVcmv55380S
ULY0hkW10ZlKiHegjT/XysrE1VBc0YBeexwYXjm8WeS0hlOvbV6jRnWskHBEt+4O3t6tHVd4mZj3
NhtYM59mlihNQRP3h+Pycl81wELmfcnWeHcePcQgdKtYxdtMGTJ5x16Ga0zP1i1kNA3BN60m9joL
dH3nLFBp1ZUuVH3QjRHFaOHotUl4Bn5KC++KbZ4IZt2rTZhSufKVt0EO/LdDkMrj0uuLPYspJgHn
dmbMuVirXnE3ljuB0lmxYt1XWn7UEl66Lw2bydKeVuHAQO9c7ke46LUkjGEdNldcZ5QIVIWWc0Yx
+ouDa6vj7bOjUBqKUr7LT66E9VkE5+imm33H/kW7Ttg++TQ7FmxBBN6T03U9z/5TlGl0lzTcPzht
gwbbEbK0q9KUBxGwyVZyE7QIk4jt/nnY8S+s2N3eWSfoIku+sWbfvEXW0Wgoy0XYcGXL9nzmuVEf
mjsShImtVeRRVlvCQR/xxpwoZ5/W9/V5mZJW/s9bylaErk+nELB8J7K/eYKFLK1yPFI+wkwYivoc
6eqeSgGyU7DP6dPXvbDe2bfVWkNG3xs9kIsdSgugIx+fZn18c6w9qBPG9+dkJFUQq8rgSe7TzsTC
RLuWSzwBEk7NtL7JV+zfWNIAeXX/nJmhv61mZBbFvrhyeVhC9L0MJ1INl9AwGKpPQwqCfSz9PkuT
2ift7vofTNr0/TaHLHE2j6AGZr6/yFGV6Em8abAZ/+8IU6tnEMsz3PKT0uQm/C4JfWwKWyfdpySU
ETJb6lDHqbXwe3/qdQsFvuiP0plOcEofH50VZpLlPfT2tca4rcndJI7pi4RPKynUTMP1hNdM2PAW
KWns90YpJtryuqkjCY42zAwTR0erqvCgUJdtYZvMISvPaPHUYfxkjX0w7sWbyApwS/QrBydLrOGH
ELnR1ygN0Np527SaZrbh5fTeDO5/8rxv/gnxL3YSvLQoRPkg6sEgcTLuxe8mKJGN0U8cidGitO9Z
JjakBwPxZjFaB4qEDeJB31eb3hHl9RWA4TZXzM048W/TH1kk/lKL8NQe7YhF2e7CWR1htodiMjZp
8VR0YmlHQwpqCzkn6r98il0at0+ttlyARgDfXP4tSkQ3BbFBV6jOspoWpJvaIPA01XZ0HDgrKNsP
Hpq61/kOGr8kWQZrBhtni2IBAi0dsyt2wWGsCkGp1IPb8RUelovk9yJEUGXNODFdNBpWyED0EKqP
mDO2fszHlqTModuBxAAD5maoN90XN/kNcoajJM5Qo/mwcgz7cTtYAIssqqB3nvQe+Zi3fQmEkHFM
juCqOLDr6vasZylWCnJE+3Nl3G6RosEKLcDLMuEmpKJRYk1dcnJ5j+7xv5DjyjDEnjUWuPDNC1O+
7GjNMRL+LTTE24+Y5+5Gd7wHwFCmYNkq9V8AAzN7RBpTCcgeGLnR6Zg+G5LbLFp+ATFRv1n0wijZ
O4qzF3xfTFMDHOpnGWrVfE/y5tOFFqvcQB6YoDBudmJtIeYnH5REHFgEkiW3lb8e3kQCgQJQ0Haa
SnaksikID7ZURpKPayY8J+BLon5jr72wc15baKwK4ZPdKJksn1GDgtn+m8qxu0XsCtAuvJtXSQpW
NS/Pw3X0p0WkVp3OnSxH9U9eGaDhYzMbtejgkaYkXckoGCqDfImHNtux6b51X3q6QKCAtfuk371u
zPSHKrecDeP+LQh15WEnOp+JiG3x8NSdIJ8jRGRdnu8Cf0+XHm45hyIPdHwbA34Q1IQ1HAqSVGRS
DLPQG7bARcY6PCmCsRdCW7bKMrWQK7hMeEt/0xq8zAvKjPGotphKWmWF+nCn57jDnipsMu5IaiKL
lgfUkTqU0Apjs5QFucty0EmeSI6GCjj5F2ZxX6AFGnC7ughPfPI33Ps+vuaoBggBSuJW2kECwrTr
6fKqfa8ZyPc8GA/W+Hd3oMRRMJ9xkGhiBi1aL0JpOZqmb6jez94OugUPTXryRh2d5gfm5K6YUvAA
2sCSvUpnb1inWzSC56td8Yai4jRCh3+ka0KI7iQFtwJryvaln2jzAdEq4zTcagxhDST8KZ5VRQci
MS88gbx438lm/7rp7RQe0t8STu2KrSn5jet0yeGHPbcmd25LrObEjXVWNAdVjfWAjJtp5WyQ00Ud
m8AJorvcnLaU/rB9LX7eNAO+egLabaWzIaCMW89OQVvTHVBTwrRalJZb6a6yG6BqA0dC6HGjFWyD
QkljLQVJZzUnEi/y/nDg66kMsS7YBHW6iTOAnN2d0lIJbgcOBgpj6EDUzvgGL3rkO9rgVCgzfeJl
qaWhlnNYX52Pnet/CxMdxTlGKuxn9V2QMu/N1c+bsbSjeXXTiTKEuUTkVCNYd52IojYSN4Qh5n/X
Ccc5rfKf/qRTFncE5AvXOUSY7vJKJQEuokILf8O6EqfbzKEZhhVC0uuaWN0nS8/QKliRSLjkPCMG
6jDflZTGxo7IqjSnzVy7kUeMnUXCt3h/XfRiQJXdWUXTTR+7m4ub+ULxlrBj0IyA7ugVUAPKlRSp
TUGY7vhet7L/8fmv1CZy5BbP0bjRFau0lDDg9hDAttGOq8ifk/QyAz/WfrTKIX0JaTfhhQncM0pD
s75TGQahlXemV1YuZlHoxLcwztkgaujQj8XhEmXGMS+vQZyWfQgntTLdhdg201fqNHnhSTy21yMV
f9JlzeP4QtzmNTvE/XGYR4+waquoK2CsmPqD7WoTWsm+OQA/s0/jrvY9RhGFyiqLSEakvG4FjBUE
dQjuYdp+p7cvefinooz3pmTKveMOmCTbYALRK9v7PYYd6VRvEBGoWcKDxpsEAiQg9e5NAzdskk3o
P7DyWzJNnLduoG4RFgMht4yxB82Dk3Nci9jaRDFPzTv+T7FJ1OOhMDs3ZfFG4cQUWRdtL96D1/6/
enHYlKlaBzjQhBLzYTWn5HrHzXU8GKtzxvoNncP4ZL01fuwp1/PzURT5McJDi9nJX0twNfiSnHDG
Cb4mvcLVrL60PEYi5UEQHE9WGzIMi8PleuLN22zmRd/Zf8mbRsvR80E+t+TIPt8n+T3+1KX0OkrA
MiG12eD7KoJXYFjgRxJ6tfPp3Yrsa4c1LofCmlhRh96f4/khdojb428JQWWvYuVEqZ4qCWnYVob3
kVtpndpB842wkZx3td+JtN6kOiS/zivFXS7iIY7hwq3ITmI0srm0P7iE09uBeJSGg953uWBYf0Zs
gWThJKEl7DeQ+L5YnlnDuDA6jUgGvQb6GpjnIdqAhfcEnWeLviy36oMA/CuS5kGHwRJOzD/EP5BL
uz+qSpPtfhCOuv3bmjhmf/6ymKsRZmk+LFoVwKa5cpTuxA1ZDzhp0WGe7Ph1L8elXXZcqBFsw1cq
4Sp2+N9pYT4YfgoS/YRo0tYo4aqz9MWSeDPTwqdvsDpPF3jKCeyosM+DSkkJmcYUzJRVIcxcnIjp
PyfrIXR4eB3fI/wg5qubLqJTiVO9JgKpxaMdVoQRqp2iUVWlkrCBNU6a7yYtcZZVLdms4jKPXvXg
I3trU1ACDbElb6rNYKQC9nP5LZC1gYBIVQlydtUjMGLVgUlreuif5pwx007M5XPcBsVvyv7eHrhv
vf7Ond/bgWIOe9SAPz7k2q6VEZJJxhlGjPWhRqUCcR9uq4KvAd2EpDUyKXRvcwsPZYCZL4YNnhI8
GaVyybkwIOU8EF142/l2UpY1ULgGX9sHssqvxcCdK5gq/WDMHJUXH0psig6Ciy9H1XHDFfKtFnEU
e5rQAKU1JuS3ilwCbQX00YiWFhPu82vzhJuFxAgf4PdrDETME8OJdMTaX0oa5eWze2XwgOouQ4//
4iJkT7Yl4xS4C9VFrvv3iAD33INbmHs0jM2iQWRBchwwzWa3DcEenPvpj2ljQRCPDtPlYWPU+HNT
hLp7f8ke+iPIR05IavRxXowgJsl/jhyTXfwr8FexYy6aGoNCRtAgenoijTjGLifrLrm5H9RT7ZiY
c1J0322TDgmwZS0KSnjbJ7e4t89Nw4DPVHFaG+Kjsxg8KSs5oFhU5ag5nD/VKmLVZwNvaqXky04m
+yU+9Y1P/pzc0t49WWN5XuE2XWBS4Y3AXCC0ygGDsFMZ06AlDZNa/WKJVtKAefF/CP/Rxxd5jYV0
tLmtE4EtVO5yUXowVpoqbTh3plsoNmZvqqk6s8WSjkcktj6z02wkPzjWFslvPjGPhoW972BNpSPM
yiFiHANDFWv0r+hkfgoBfNnkiIQgGdR1/M81GHUwRAp5d+wLwb610mXXNx6kRhTZF1YT4FFwDc3e
gC6QIGnJHudEy0up0rcc7bKubP3NYa2uw/agIteVtvG8Zzw1Rq3C+DFTSDbQwN2i9ZZBYfmP4YW7
OkscV5xjyCXMl7zaZ3kQbFAg+BBZB0fvcru9y01lLarOAFT6fw9KtoEXVZ/zy65BXeSkWmUSog8P
AYKqa3JiUkt2iPQufHhhe/enMSakjUHhUBw0pshO4/z+5rTaxhzHz9lOxO2ABrbVdKOc+c/nzpIP
F45nGaA4DVbdJd05ETWRTeKrEIcWmuaezc1r+u7T/ZjYTmTv7EOrcbq+hHfk5f7lSTFwkspscbH9
PQR7V2SzynJXX/ffqsgY8TtuTPIKnvYUe/3TDpr1h1HdQMxGix77U1xXG8vicBpIt2BNk2YbTJ5j
aAq6r8I666IDbKh7fn15O4tVEr7nGUO8V8ZCi40myHk4z9h6ltbqF47uRpYJf6/mdtdDA9FNf2cq
0r036cNHZMHD1f0SbLYWpWkP3hwRaTe5dvt0QPioLkMLwlTOYmiwqy5RPf7xNyqSwNqqMqVx1Nnv
jTqp6LpM5TnE9L9Zc7SNC92XceFYyFNggWmtIY4Je+k7CHcBNMyhmlzBp/tUV8cPvH3cC2V4GKrZ
v4GjSFd2F0dFxEfbnjG8f+Ee0oh0kX5kcOIW9n06PHYdYWmrpAYju1Er5c4kCD9AKcMwohmj8/lW
gEpyOmpIlvDRcYpRR2WbdnA5Ooz0hKs3pFMdKWk62uYq3fzxQKU9PW+om/Tu5RRXcCfTaejs3EUE
tNY1VWi2q2wJbbdr8DbjE44zIcHPm455jXaLJ7BQ5lUla9j0EuPg1J29EEkTcSFDYSVvTBqq03Dx
HnG51LjGKWxSw6bvuIOUYn5hGtkzS7k104r0yqRT0ozLRWMdv622hworzlhZpdbaVCJIwXno5zu1
Soepr1Oaa6SxOyNDCp8SnGa+zcpDtMvZR8oGmxb3SAH7qw3YdIUOaWy1NA4g1LfHxFwENEwDIob3
rya/Lm2/05ZBn/O4O/QUV8ZNcdZnEglSfKMXdTvG7iA44Z4gS6Tc18DI6JYu+vm5AisOwfr+jJrz
pS9Uo1N19fq2SDHD0fOLTW53V5lbuyibpzH/DbT6TxY9Fn98y4BaFaYn2YYma9k2jFAzGjJ2ewHn
bS+Q6gGljEHRj+DUzzCkZuUGnpjx+lM497nq9aiRWZ/R6/I8pSwn44r4bm6N6Ztixm1CYN4PvN/t
Sp1OmWU6y4Ib+wjxp0aeuDAtI8MoczkMFZTmByRXx6w8VBAFMmjeLcnH6ORjGUN5SAlA6Cz/+O1N
I+sNOPztKgKB2/Wz1XVGU35jjKdkDbiUXrgMTX+d8y64l8DKMeA3Ll6RARYfUbxDWBDfdp5cTKJ6
O0JvXxnIrSZCAND12mAoaBVyTmu7oZ9DOVJWhwJg21tqejdIh3+AcCCQhJLtnOcFsgdhwtsEXAbf
tQ+pUN9bPLmjMbGGbA0AK75jEoAMa5uXOivxv15Jdtyfgg6e4v7dzOub2EQLMxwcAAn5k0EV2rBP
tugH/IR2gmIvBhAXj9QmCNalqSdWD7ZS9VSjEWRaMiRu1S7Xear2pb9WziHu3qC+6c/x5w/HxYrk
QQeNuJmUO48ZR1rIATeQd4bxENPfFLVh23BKQHYdyBJd0d7Pi4Q/k0kamGAvl3jb+erFFreT5BPL
/Gf8EfD9iz7zhVF2/+6G/0JJUWQ3gK4OCsES/OEPUeYOgJzDo0jIg9tSkStTUf8mNFv1AcuWbmhl
z9Ov9RdoojuOwimOhdlzobM49eSHyhkLh6XORbwwR7SZpmTC8qe8O6WYkYkiv5fQL4ZITyTB22+I
ypveb20gk5HbtNFRoYNuaMMkcFMl+BrR4EUpMDUKhwKlFWQWjJxnYrV577oExSKLaJIcneoSYIWt
1GyTZKXOLU3kXycdsi2nGtAcHzUIA/cl8Rex9NEgIqkzI/8afPKd+LyowSf6iaAlbIzFSwtc1/Lb
Sr3TizXLCOoEWjA7tfo9i+OKH75WsvtsVYV69+H4Aci4NV1yIa00kpTB37UtP0b70XyqWHP1t/TG
L/zJTXJBPgMxBvnfUah/Rd4n+wnEoVaNeYS3q/4gjPo3cbnY20fqL6LhUurHjamxA8tvTMZ6Ekeo
oRL1cP1TUly2hPfAP+nv4bc/NrUNdYa4XYfgy353X2UyzlKxlako+PR7SPsZN6h1Jr63GMXxFy8e
JfTWxyJzFeh1jMwh8qsuihMNCQk0h0QuraS8Hat7CukWOGcNfDfrhf6i4YYrQcT2Ni71ieccMS4e
T8nhJU+07q0M1sj8JPXj15L/5nG2ZcwP8cwHEt5LTJya0vaMXd2CUSVu8z0/c2dldozIia8YAmaQ
i1YtodwbuUtGPX+SaZIAcrUoRjCBOwWz96HDt7kx7cMRzA+0nQbk7o2SRfznNQ+4KrPM9WqdrHZm
8PuD4qqIJC+4pNElKh8JxAr88SyKzx6F2UnFzcV/d0LuEhs7sphTV+v2Xl+00tKjE9Jw/qJAXv9D
U3Kg1HoNCc3EAY6MKb3X/J1XCOrOBnSOdRE6YMHBtqq8uoDDSNRlKIU02kTZmJTlTOUOfPi+RMrw
3bhQyMansVWsMnJT3UBvEws3xeQrJYqn//H+Dk2BuFbQ/d8nKvBzt/vRUeD7fKJyzXD6kPCES045
V217Uitd5BNeTn7iipOGHPKX+2rdsOE6xjhG9p1RI1q9ncPmj8SbTqfaEJVC5F9XlgBrmYk7Zf76
HQelDpTZIFrhk2ly5+lnpUrmNqgOB2ZVXPWjto5MO6DGJ7uOf+RMLrIgzSWUwHOIJqHsobQ8hQJV
xffjUUYKBsR+8S55+e3HqWDuSmCkMak6j3iN6SBVlkqgIfFHcUxlPzSCzRPNF+TjwMnG7Ax1XKL0
R7P4vkk5N3qH0Rd3UbktJeR1ED633h+7NCHr6ka6XOvKWGOqz9l8ma4n2tADFDx7KaJ406Rb/sDw
5jBgLyCVvlNQSnqUT0XtTd/TI4Nw5QZyX8S+g8KeeoBznkqVQbF9UrOvYWZmHbyosBpkXhM9IeQM
gY4NImfiz5C6NDg24kXlVZPuyFHNz1buPg+8LV6QLNffyZ6PhfyMea5hdXoRNIWlvtWyj77b6Prz
hoJMRueo/lm2qxiRkjDIMk3xhBVyIQe/pRAjCOjzQLImCM5HPD+a9IdUITgbHJsT/Aa2nflnCnBf
BBk5m5QVF2s8tYeJvRCsOwD/Rr6bvf1SYncNNXZvF1nY3ILnv4CbuA3+X50GYH2M0APSN5Dm3zXL
P92VCmZXTJE6gymodyt0twOLHMnpD6MScw59VnErAqmKnVQJ0jYuW97A/LCiY4OmarS2u6lypuhj
D44UQlUrc2PrWoE6u7owa0Rt+JlA3Yy7Cje4CCXwonW41hJO4AmPSARvfbOBnjPFVUI39FY4wzYN
kbXp+lPpnpHpKhq2cPpvUKVu7nxYsJ7nw9pciQaziHvkSbB3Y4qVZtub9JoOwGZ6KRc3WcxjoaY5
DH772K3ZeQeKa3b61viOo65uql8UR8Pft00vfJOjHm0vlSzmk9yAvXuT4cetr4KGwtSvQZhl1M5u
SPr3phLX5B9MyxMlRmtFL2rHiJJcCKAL8nvbsZgXw+vN9u9BzWXOoQLp17DLH3R7QHMu0aOEqd0p
EQhfTy9gAWhUb5Kcw96XG9xa8Cwsmsk1gx/YbxEuSBr5E9AaBlZt8stKN0aAUauuLnIXKL13D0sW
VK3WE8CMGZityN0yD7PB90pEMx3Se/eYXaNRg5Q1jPwY1Ojx6r49ASXdMSVIE+QDrOYNBhsCQOYt
1B0GeC0PjByRve0CWE0P0s4RcqJIeilnDhfmpgHqzvGsv5Ey/wxNQq85r8S3VSuOWksf4WCS95Tu
EMnqtQBX8WUNKgsMguE6110eRLT87lYelmalH1yzbaK8m3qRf3OxKLP1puACJy+iTxbd21FrzUeI
9ZsNO+ouhBLSRudGy6bF3P9q51Ywf6T4ZmhxwwmOzrzuKJaD+dPD2CDetXouLNrUoAP466WaGLWB
2W7qUO1X/ABczTXFhvX7HLncmGwplg7oJVCRRrmGnoX9c4viAOC04xhK1eYEahehUeyLeO+ONFP4
/HgZZAnY5x7m2AkUmSBG98z2ZUuW7ofQw6HwoWX0Noauj1nHUn+d4PFPu4Shgus871iUf2JglUpt
OGfr7Udwpo9R+GnkZQw5kHwAredGCAkSBfl+X9bfjLqMmv5jAI/BUxf+BGDC+vwHljZLIc7cu/rl
lHjx5pAVH03JBDQRersOTJaV9diT2u0aPoAiOKTT6LdBQwtPX7hu/TN9TYl0mI3fi08Z5XP+3Ml+
aozuwdwQjveEmCUZSRf0TqH44xOunQbAVfZTaRMGnfg7ERh+aFfLIxOLI9EeJoJYD9z1RRxLyb85
VK/6CQ9BIiwpqk/TT3rs/i6kjOUIz69fZ/6DEEOC5qUNb/5Ixq5P/kK4/sn8TiUKiK3sgqBA1HAz
GynBuKQMLsFSisyJxqgImZ6aqHcB7QAXir6M2bKhyCfwBrXokN29KG0lo6gEizIXIEkAt0At6dIJ
q1nybFYckuJRndCCk071Pml0/6WJDL7dSU9hYvz6YTbUzXwro69ASZYob7/CgVO7gHN8jqET/LH3
1wYKvbexaQROlB57dtEUoIr3Rue2QrVNZtaJUv+uqQMpdb1w9SLOxaAjjO+h1uRH2aPHPR66v4QA
Kl3zhqo9B6omiGS7JZyduOhuK08hiPaxH4p6HHCRwini0Ni/3DQQ0o6XKiu/L8+/TU+CH/OOwUSz
cyXoJPvTUlRef37JCAHOhEtnP83ik5C6TxcTBjMrvUJXlSySUgruLQw7MCfhbKdeS0ql4eLUdUX3
qEVw4MVTyS9KQNaX08LG4R6WGej1NiX/EiOuqqUjn/bHrWNYqW1KclTrqMlQukwhSR7ix0AFME6c
dPZkkHvUPb6EMDk/UiJ23z1J1BUiwrsRPnbB6wsNDjJvU+xtbM42D1ia/M2XF/6LCA3Nw/iHXxgy
Q6kr1okoCQaOG3qv79lDxIBCS2242weO96/RpDW0Gkd7i0YulNzcf6AWRsRLudrXYiIW5qqZ9uLf
hb8aaByvuJwFo7L5DD+KpvfyiKW1yPVzBy00uTkOc+tbfxdKh2pkc1FTqb8pe20mDmcjL7RTgn3h
FeTGBC/u61lhdjEhIMnkiU5IVcNON51LgUATzUJ5xc/jLDlJUK1WqVEx2pIEkIUlqmZCLIQNDkYU
6e1eh0JD4v6uyriVoDU24we01wSSRl1vbBwSyroAXMXM7baplMGQcprqPWOIWCohuod8V5XAATQu
KFRBdkmmIs61MbG2sj8wsvcCcGBdQuVg1VdcBh2KcZyke+r6U8+Vg5VL3Rkl3fqFgWiadhXjZR1U
GNPaTru4dryveh4X4mvlE9GSrN9U8ibwmNxG4CCDFSsdcAvUmakxZwB5gKFj0DON8S0siQoW/B6z
h6Bn8kIyYTs6ugUaD6LYD1CoxTrJNzbPCAOvTrQTMf1oWs5z/J5mPcxTKBu39+Fm5FaRA53n/Iog
tH4S7kxp1/bJrSO3E38GKLBnBar7Kvn4cQydv2Xaz2aorGht6M/4cg+4+N2eyEIxcWxwQQxetboO
Z0E+pBSAmxU5YmU9tsVla9jd/ODsyhVq5BFrDSoQtZ7BxxUOuGudPAMtPVrSpTpiC4kN7gORrAda
qjF1d5oJPdKFA+Non/9g7ps7sXSiPENTZsbRQi84Tg59D1xJixYn+Cl0mihFzdlVwfuN7UAy7kvm
EHZALrvgAQeTA15sRpKfA11OfG7cBaYTaJURzpmQ6ag3ga58LBXHbgUQ09xO66mgtCXT7cIkkRzb
FtW8nlujFU4wAA1WCM5mGkqsE97eSfynGESu72W9hFmtKmRXoM2BIVRCSpa0bW4iq5f8Y/xon8VZ
B1LzSS2X2HbAsD3DkqCiofUbQADryRyLImSpdTCwW6qrd7c+isI4poeEb9OWBwlyhHmXRTLIhtg6
Np7Ica9PyxNRA6hBuLpasmg2miMVUwLcEu+Bo+jvaQrCnvrmzubaOcFaPN6ddQraaljGAK6RHVBC
j6z4R+9LFEQ00ljPh5GnhUkzlzgGu7a6mOV7SzuQLJ25JAeZaZbQjZI5h03rT1V52tYjmljyI/pf
lvu1FrbuVwgX8osusTsrTYJcoxZPKq8Hv+IyCZy94FIpvuqXnZrUMMgFOpQGwbnhE1ci9eOtESGM
uU/I3+bIHvh+Jvxi1ZWLafW1HSJkywS8t9pG69RDEOJONJHX0RAYmhuNHxPdaCW/nS9jKujQ4jUf
KXt+Ri85Ih3AJqEoPuCE7J48sas17w6z36VEfi954UZkyKe2bMG/FfEp7PVcBd54JDElaB+dLd6Z
XtAvHL8o47VutWDM6ZB9NavfTbtt8z42jvdudDNcRwS4hjo69zdTbqAjk4rp8/PR8CFa0Lfh62t1
KFGfWdhsCiRVm40cTJR36y84crGn+QPbricxkaKA9WfMDxamG+umRJQkzLWd0tj7gWRDXZKut5cY
mHipfa2YlDWJCy5m4G6rdKW7PT2hP4bPT9gxN2hL9X+tvItGB9I/ktCNqGG6VlRZ4UW0san6e60l
aHP/jM+YjndlMi0EvFdi3dizcjTEcHeL+wa6G5MNpXP5JjDWOMel/b94pk39UnW7uXjklr2UlKDc
yLs3n+aaSb0DFSZsbMEEwzj+Ix7AX7HvNmF1BbWn2PiVJsHYrOiBsRMTd+5eB6RXL9e8x4X+o00Z
lswOVY5bIF5uO473iNZl4mz7pUQPLuDjOjR6JWjm9T+fGTlgBAyGXKZ9d1PVqRDUcQKQ8dfP6ZPY
02YXv0Q/w7miMhd6fAAYnxM2L3tMlb6I9ZlYHR6OYas5cYTYb28qKhn0E3n1rbpm2UUr43G0DqNN
ky7ev4PG4sQPmpiSXubYK9jFdk6wZ6blvUy6I+uU9GVIcYaYUBjWG4mceWRTyevN+BKeXFOjRtId
fT098uNwIU6TVIvnma9l7DIh1M6JwYyk3229eSN55cXUic7/RWVKGZ5BRqya0xEmF8nS73qkiFCC
QVTS4jca0uDmQoWJIVu1cA36ItBWHx3os7aISg0ZyvbdqOWCz88y09i0qWsp9rHTF+93T/H0RBW6
KLwd+JBckFW5Pew6oULMkMup0V/xD3K8YRwyt5tij4Y3aP+WyIfvtPp8JF5QAfXo7WXyQqm7AXV6
oy6W9SPAESwn9DLep1mjl50CO3F/3/1q+r4hlh2Xr35cBAP7hqowBYq09xfx+VznbdY2BipfFY7K
zSU8yu6zwFZdJbZw1QW7fMXDnt79rLU27aLLv1suGrXHyvMzvBmIhkn/qBI+idj+RW0YNtF13oS+
P9pjkAcPzIJtIv4e2NGzGP0TuG9Bt0xdKP/qsMMH8hAqdsTf8TlIMvBg8HyfdpLugqvIVGSacfG6
6xjfxHmlT9AeWWTGw9EaQ192pzmVGMTcGkZgMPVymk3XGK5TGS3euOCpFZ5ni7zw5nKlFwMz7tx0
R4Z+IcgXi7Y7S6tUK5/X0F6FTWCCbcc7bk75ja399y6SYIIs3ll1o9PGEu5Fwk9ntHZW6V4Fny4z
U2u+PMm2UFXbhmcEo9fYxReHiTpw4JfZS+1UFppYiulnd34oOJbwccFZMqO5bKREN42ilv8I3wZr
zPEjWibxlOO4rma91bwm+MOXin0wxYu8qtH//4fTqPzvqyYptqvITZK8cyKnovx4hFYxD1djItnW
4BDNf+JYrnPuRIUb2jqftiZPqKplb+GReyPyWgmz7xZtPnjft1XGKK/sTGJJfA5OQUBWme478RYF
kNrrvtATdzqc79WHeQUC+C9tMUtGMK+oQl2pUOuHfc4fK6gt5r+9QhSLgU4Z0dX5YvRyiSYb3elS
7SSYojUwS4lX02aFw69UBAMnyHj2iICwr15bR0QshNJ1T2pTz3zJdX6pvHvUr6Vy+R3pqAdJjG3s
UqIOdK9F8r6dgREJ9YWLSmCIAhbIZqp7OtegqU9cgRW8AopLu2p05jZIvJcwaeG4sC1JACfQ2/Ir
OJ0JuOFf/deMox8iqatWbutiCYFuR0cWnOTx/tW3AZYOZPLSVAPt24fKwMmkRvPmL8TBEVPs1EOl
MI2tralPHn/GjvdI8Ky/JFWFdr2Jf7aHFQeh8JoRJEVNVrydwj82wGW8Y8ZIxuKsPfhUBZvBi9b1
Pi7445iKQC+Sk+5Bw3ycR6M01Z82Iy0j1KpxN934gAcsySGqvDSmC+SF3QFuDUDVXPh9fAKSp7BQ
syTouA01GQds19d3TVi+C38ulgekbzMFiU/HqDAN4tCnzKHsqCEF3uTPJtmWJVRguGBw3/5tD4Yw
Q7KARb5GtCE+nxXM1LZlsRJ/7X/NiYsIu/4SnLLz/FgFdkL6BTwDK1um9PNW4HQoyEsW8j86H4X1
/htAmTTa5d1T39dgpRwThtDxFlTjxay5ujSLVfFgqz2+DIdQzoVC3k1tSFT+/Py+z6T/O4vuBhPJ
mzB/JI6SUo9k7ba7km29vx+0QPylcNQr7ZmURQNQlIGMX5Xjcefo8OCq2H+DE4ZnMNGzcAm8sict
NaLNNpjwmf4WemycaioUCnGoSBhj9xayhzJC6Q56WYxBNbnRqM1VbFGBTSv1uACjDoj651dizLGH
6pGO8OUsFoEiTWupzQdIOF4Ogs+vQqMMClU/xTP6MV9rqUhhM5HFlS0afRVyHBFx5pXSaF+60hrn
ng7UnwP0KrArjZGLrvCF+mvK406/EPJodV7536a7Ku5Qw56mXANyK3Wc4zZTOg+GbyRtb8loLrvP
SPT9DRTjWcqSaNESR9ZTFQ7u4A26c38D/B5OisypgCRUKF8MxKCpxZzoFpLUaajSk8wD4gO6mjUe
/vSQPsKw+04bOHGElpeR9QwBoZETChsNOAfqR6Lr2+ALSs4qVXTtxzc2NeQE6XIVPcYZrgKxHpkl
xUkEIwLbC0pCQjvIw2XgMBOG1/qWbO7ew0yhjExlZN4UL2d/gE0MtasA7I+SOtlf0JU6GWu8p4on
s5q312QroLOt6nbI8XOYhZs/nAmaPe5cI6zOyg53b1Rnv/f9DF0Q4iVgEuHAY7+lDnBUfdmNelAJ
MtRsn3hy5NQpH+EQrjjthl456TA2zGv+8N8Hj+GBCzxZxin6lPrj6WtxjxRNGQ0AvUqu3D4d1WOQ
94LbTSbGrAnTH0D3R2uveSsoUzlT4OIBui6nHNs8s186kdOdEQlTSN/l9jxK+tWEa60k3k+V2x2w
yox8VioY0M69VIOq4OZPZ5463TGlwYZ+dn2KUGaZn1/M7oj7YlHLScLvb2JlCOZPMGCYXGtGsg2N
YZzj/VF3GSVOg+FGqRCINvbZ5snWMAX1NUN/6GmZUW64Dn5iOmcmz61iIW1srnpBPdd2f20Xt6l0
b7/i1gTQotMUrctdo3W9CZ/L4VGb7RfEaxFGzHWq+4O3a3uCZgFPy7WJRdiAf25e0fADV9djI6wv
O7Jx8e3DjKvKScaCsJdiBp4RCKujjLaiV5z1Au60Tgit5ZkR5DbpWJzOkRpekUwDbb8MGF3BFTie
s0uUTKYJlyvw9UyqxqZVrWdflZtFRYH9F1Knnfjk3PJCE9uw2YvO+ibvmR6DAIX9Kro49x871Lme
hj6WIOrgkUE6UpngwcMgViRwIsfUzZ+25me0+XuW9775dbFF5kpy8GQZL6MQKHlSnZ1mD51OXg/O
JURBGojyYf8TrQCWdR/Tjfudr+CJ7o7aLrs/OuzAMsuP29Uxoxr9y1rPekfRl2eq5mtwQK+Bt5B7
ogQDf1feZ5y5jAERmtxKgZGVCmNit3lOMKdvFrd3+UqXj0aVtGUKyexwifXH5uORyIQDbKZpng3l
J8AnZFkum7+jvcXMt3Beg5bb7wlRZHrDRvfRR5isveJlyxy1S5c5P9xoLYO2CJYOnERhb84LoJjH
d3R+ZwwrclhOY6VPGD1njaSC3W8oURNDaVPRzys0XLzhB0RrJES+vfspAx59hLZdtZJ0TzUXrd+t
AKMxwJzHYZxFMPnBSBTQ5hBL9ANsVS8tCvSaeK3iGb3UARDSsgud9nADBD7w4Gn0vjasouZSz4EE
KWXsxtbsJ+lJgLv/EH3DBgYIUeavIfhfXMAXcDVLZnSOMkMjx2hkWd9GKsUXaV0XCM6zyYHg/pLa
T4cwDsGIyTrZ9XwZYgeqdzYneVFHHlh0pbJrlP1EhMxyWwLP8xHEiVuSYS3AYlnhqVxUMO0HkXvb
VtpObd5vrkyba2mmRq3Yv2Nzy7anzp/v5InAPteXi8nZYV0SDvrTE+YYwYPw9A+ZkMrjlziPp1j2
kI80xEz8EUleRfgkfwI7Wpd/OM8j65+hQ0JlE7j9YJE2zMgsjx55kojNp8p0fYiLn3l08Ioap/w4
E4VT484Bv0/1jDvP1cLTMR7rquw/8Fs1iC+hw9FC9uPxprIhzcupyucpqzgQqofsP00Cncz1O1In
YqP/V+MsZZI7C0iGYXQo4UUPutBaLv6A1lnTRSIv/02tp6MJKbysJEblUm1d5L1mhuWGELTj7H1Y
/YYIdnXdF3X11BCEbOBY4WrAtxfkQvVoLJfJrPKS6V7lgxfHsQsX14CybyadlmpPL5arad90jCtO
po2+G0uh69dlLn1fXvXIDhhvZpjuz9NgPIvM0K26EsNSboPc3hRG8XHX4QY62Ci8Gfoz8w1vsxl0
P4l79LEjAVhKJS0SQ97P0XrPK/o5mbM8tEt5KxQKLHqmfjFhN53AL/s8hGccYcYc97K2D4V68dcs
+0jTc98YKfcLW+Y4h/aCj521lDIKvPXyBg+GZbYDmVFhhKfBJrs+1ugPuc493XnLHSYy0OhcafCV
Ucb02N+Wjwi3ScKlO+gLyeDisqYeeedUkdmlqXOf7BupWBO3zPFtFgsfQvGJ4ajbVAFYE+mePGGz
uX1hfaysGJfiIcro0QPmFFiJ2IA7o3p/JPYeEzyvjNmgC5dnyrJ/dikrbVmbyYxBohDDTdXIRMUf
iHQULh+5W1NpqSV/TODzjGXZSx+mdqkcIuJnMXGQk82l2df/I7dullSKRruLfp0Mw+DsaPH9AQuj
9KY+Bgo4uNGa2FqQJCF1znyph0xmA9wrPokJ7TWs76TAEnjhXKCAc6fkbxVKfkOT/EYmc47qP32B
87CYgsu222I3WvfM0HsQTCrs3Vrlhrud6kcvNDgXzOf2KDV/x0LfRKa2Tb/BH5FC1rEyC+9W/5oI
m5eTdLW8DkrWUdUaOqRHPWJRQxvUi5tnG4DsnciATu6ixUwvghdAXeGd7RGtgUPxDnz0ZtnKTAR/
CIC5Y8OoB9j2p8xbMbgYGBfvrhlevN56zw83sOznwtCTBfpCAk8Q3O/yBWK5wItBc06wetDh+z+R
GaBTKqi3nNcAddu8TQqJzU+rmxPu7AmbXPKMh7B7WMUTH9ywPMosWSC/8HDUmDkoBwcvWXVLUlzx
OqWFsNkjczR3aRAB+Zb/1GQQjcnf1/dyLSL3cKkKJ7F+WlsUaVaTvF0RYVALtwycAb+7vzJf2cXW
H3j57+hJAQ/PpfyrkAXEbO5e1Yhos111R0jpZVkkqE8fjDrq2NWjxEGXdx/7tcByspUP30yWfcs9
KY12lRGStrx1LiBQ5wJ3R0/0Fg8EwgMNirBo66mjLq3hsPC/OeA/pVV3EIQxq+o3fRJjgPbjn5mg
BGkGRmshoCMeYNBDAbc4DEgCMbhpsJrtPcl7kqekC1NmUU9ivkXmc+aOMqYO2fH2HBua6BHKjSV2
4EEd7o7vm4AGzWnNMYuz9iqUSEO0xOUFQdG/L8VgUiGm80KKxs9HFbBV6Fl0GtLxwXBm51D0Y4yb
1h3HzGeqcKJeRKkDZknPDGif6EhKNv9bppYx61lUSszLb5zquIG7nE48o6+hIV596+JdWZ7VZYYz
20Ty9+NU83ft3jM+WF+ufp/sFiVN5gWgEj4smy4KuXboozSIBpGLSPLElz0iwcOgVwC9Nvk6r34L
jqa4vgB+ce8mXLKZpoJpE190EdDx7uaVh9AqqZOuB/zLHUAQTbXfOjeqfQp+/Sf3YGDUIEHyVTVj
ab7WkWpcG+ocwxB5+qOBF+ZqwY9lJKxSuvWbao2PZJ/v2sLGbJ4euIXYuAv+GhUzU4dCVQ7rxBCd
5L6gl/8Icn7yHad1k+VKvoOzbWHv/NyzqA1B2KIqvLVX7lZ4NThaPbaCLJd6PRShqcjeXa8YkqFt
7jvs+4v4nLnypiZfuA82M9+TJmNPlACWkK5pfzHSQ8YXHewSdgPFEOhNJS5ay7/lO4xSRZNTiEfJ
/uznu9W60dAJrkVRHqJnFTHM7X5O2mzHoGdQ3vncC+URR+AYNIqBrXjgZ+LcdxXZTP01N07szwvc
6pIkTC90wXLVEOkVmNmkTelHjgQjOXpNSEOt1G3KWpejicW0iZi2nl7rxrkIhjHowUk8frwA6zy8
D+4DAw24f0oh/xbGwHfVh5ApzIP29xyaPgV9v7WMpsbv/gQ4+laOWe0MXlqhIf6XPYjWLxae2vyi
qk002Sa8sKvf6XofTjAfAlTjJVsNGKnW54EvFZOus1S5k92LWW0OBnjZxXYMEEcXyERecT1rn6QL
HX3aeYqTutQE2XkkUWKX8YWBw5XRU1U7W/juMDGTbeqBe8jDKhD2WBnwneoavJlvR6Hub07x4EC/
NJj8ZUuHqk+lEni9MDkrkd/ftadNsXSN1Z3luc+q9cjW//IYf2ZVrjmG+sQFGE5mmNUxuPZYTmeW
lxbtQMMoJewCoJk7WGCTov/0xS1yucwI86iKnc8QMd9j52Bh6QIkDmZECfF6sAa2K+Slebo8P0IJ
WLGK43xz8JSbVaLTgZbHCXihF6hvD2BbahUbMhbskNHItGf+sKFVmaETFGoQ0vJV820SEoIuRrJ4
HNamX4Db7G4bGPM8n86CR+igv7vi4zQdbAiYasI6RlvTsYr+t4efQxa9ei76s54PsP8nF50F9uH+
3E4SLl/ppGlZDQXIYE034xUw4veNsiOo8JMTGn1qezwvHnC//xAwk7Nlqq+GRe0FyfIVLo+/sJwz
7qTDWhhwoa2ZE9+1Mb38e99Oi+xosXYHfAJjtDaBbpV0WM3PQT+ivV8aMT+W5bFPEmD+9GqiFmeM
bmKV4ktlaqREO2wE9rD6ip1h3oXAifEX87/LbPkxrSU+DaJr1h6sEa/fCFnWI9DcJETWku5SuLEc
fSyDLU505gKCSR0C9WGVmc5pmuDJlssrgRXg/UuGTjiSU3dZtXPvCas/FZVFAO0F1stlThNfh8RZ
9E+Op01IddLLZfKq9Ro9Ef3Zg7E9TvTZE7psnGYo1BWheGUOKt8kxttMHpjGsVqHgYV8BSsfaR5M
QJT5vyPTgAFK1i82NjKOIzqwoRWrGhSOsvWpJD/3a5//pFeyQpouIi+AlMFcDSN8EW0hjKrvsAZq
J7gREYWsZiY1D/ZZW5cbgUY2EOmdoDP5jB/L7MgK4vZbu0T1wfzUJvZvwDkdie2MWdABawnT12Wq
9fUOyecFALbbhEPsCzSNYixglOGXdeFsYdyjmdYC3iKIfr+ikBAfHCBvjJIRRBYqoNlEne28UXF7
BSwqEw9ltBrsiixKDluqdPW0sCguE2qbCW7g5Q4YTJ2l5b1Eq05UHSZCg06f/vCPNU9v+lGiM9ep
HMSOQp41B/4CWoz8YcH4Qut9ZowuCR3QNwTB3TBcCxoC27CRc/ykOCQrH9BPSpeAFsD4Uc7tfbFB
1/VNuvnrNfGoHgTaNWKUEJcI32s/HJJVQkX+n6+xqegwvO20xTQ6uxQAPI8SYZfBwVLdGEy6AXLg
IOf4MDuuafMont+aIv5d10auR1b+qYS0I2bufz+xS+uLmW7uZgAoGriLdmoTVB21v+G+1karjDdt
RwxCTwpy1duCW/m0JnmGlDPEkVonqOtBGDpKqWrSHfv60/zmNxIO0/C2x+aMGrkkKBOY7C+WFBCQ
ZNOCudd/Rm7p/FJISol+Mp8C8bzKCmgDRrByLzR4BKsWnGYrdXxwskaUByHGtwIPUaONiMDOJWA+
79N+ARtqTE8fF1zqLbrH43ihdm7pSKAzPR7Y625Ouqc0nKzg9T1shxwjB02GzDrk5Esw9BYKMEW8
bT9XaS2NEaEMDNQF+XeFtnIr+M0wVNIZssz/QDa93Fqszdd2cgpZob9iMR8yWiNY5W9vDvOchjlZ
CKKSlqlEZsbJtbafu4AZm5aU4e6OJXwD/Yqx+4QXejlFlVoHx+i4tYmjpEim2GO1b9rPVIu/cRD8
lczPuPOkTb+Ztcdn11G5gKfY/bNuqUlMitNcT4i/ab8dVoCEs5VDvnfQm2QArG9ZXkGywxHzYWSF
HpiOK/DYmnjOqcU11uC7g8NjqmkMmBHJI8FUyOvc8p0a5647iDf5GdjQrnQCwW9Q/TsNDvlMRWJu
6p17T/Q1rjgjtq3Ows0fb7t9eRwl0ZYPc/gIpIje0rmSeSTCvDqu5ZvcEJRihArmSh6TMH0RFrqB
fKr6ip+tQB7urmRA5BmRqXmtB0OQI/T98IyepWVyPg+z5m9jLsQfbTTe5M0mtR0dzaveT0A1dR0w
j17oZk/4wAmeNDeuK0FZ4aQTgAjcP9R6cjroGlSlMCyl+t69fVGQLjv6hascRxe3G4CQ0PsRZMCB
c+4Gu4nfiBy9eBut7vldPhwowzcfj/uRHZhtRue9cHv9yXxcBnkeuzRwpU51kCxBsuv40/c0bfdZ
ZtR3m/fcQN2y1y7HZYWt+jnQGAEqMytQRD3lnaobOlGQ9/7hKl5cWx4WFKBoGZHDREsNqM0BcYze
zzilPMo9FY4UI0UR+SBP8lI1ZI1OVNszfIVU2WKWHtscRn6eXKkJ0MZV8uZk99ekgiqlcWpZAxWb
R90xNX67XUCDJWcOW/y4McYTQ3bLOHr/TP1yzvosS7WMTGXOZrETIwIGYkscHJ/cf987IGmm5jf7
y/rdo+bxynzkF8maFQ5W8i1mnvHYU4VCEb45M2ZrGP7dqHbhPl6HlVtle+Y7bmGsn92j+Mq7j3ek
dDj+v7wffJ7co2hJLe42dn5vyaEy0EszWgV3qPZqJ+9Tb53+dOeGyzcCjeTgwnTDuIbe5wv5bPWY
+C3cyl3G88jJDeI+VIYrXwl9dd5qIoYWTEaH9RI48Ch2WG47xdW5lkv9TIQt3eZ8+ERVM99+JPjm
UMeXokznx8d/ckbvUz74jfFlELRSoRxNsU01L59k9PXlRuanCCmoewV84pS1gj0NtgJ7sJJPQUE3
ECWEi4DuyJgiJ0+W8tsgwlYzeed5056MmMzqR7Jhmnthn6cmN/MbGL7nNbv0/30NQGxqlljHdjmi
MFYrcLn6aPyPparfvSKLjSnU5gGX+pFsdcLeKnTZ3Dtfl/7CIa6gY9p6NY753qXgd4edNU+jYOzo
Mf0suvKgWVKGiRcIMrV9AjrTws4rHEbRweBIhyqWCaUlkkyPOXLqZTJJVZTiFhMnRpixBrEjgCNR
0L/IFijAWmkZN6bTCKbUO8GxH767MEt3xR+y9U4346zNW4iz1/O4zleMtK+Gxk4o3SYchtOSswCU
60wqvm72ai8PB4uQnOG1ABn83JU+B1cjwwYt0X7R2hj7KqWyNrxBPQGKk4aQzyMBZL/vY0zOvB4Q
S8scN7pa4AtKPky4JxFCFJuaOH1XPclKAo0htmvtvhlGCY8V9bpLvwjZ9bUaVKIxmQZY5HlO7EDW
moixNAMSV28mEUwmlrBNId03ETEk//Pk81iu0aIDwLmnNxHLpzKjU/qUzAO+ZLfmzzT+JPKeEVIk
SqM6l9OVCn0LQHyUF/kOxuAJRyMLeUwMlhotfJaKh0v3jFMuQZa3o6OePFUbYotdf7oFp3otxnuR
VKrcPGVN+PyjAHwSEZt4c2xvtEZfLxkXDZrDKGo1F0mTudYwL3ugAjwnKjWNgxVidJkz2JpJhZtG
Ct0vh16v1o3hoAMDwNbaPtoV+dojQqMiT+pXSNEmgetzwyYrd/pKNvCItvQ8iFq1U9ao0M5uaas1
WBOKBzzWqcgekRpdhq2iY18+bdnNoH0nprSeRMufdc/IQNavgf4hKnHSt5GY9rxjl9/QDNdmVAG3
Z+rt2HESJdD9SOJuX5BkS1k9KppoY0lo5SyfYjhYYvD+xzVr/YgaqGlw4D9KoQZ0lFkqPPAZLaRc
jLX/bztlEsGx99CX3uZKXzSqbjemKhtlEdH8MtW8fTb1iWrCZMCdrqh8cloEwYuDicD5esBH3hdI
+r1x/UhsqDOgp43xtkbW8MecTU9OLXAtKHAwKJYPZFBw5//qZElfCjRK/QnUd8L1F8rBh0CQFloC
CEXt6eZ6zJmIC8HpLFeNFywktSa5sD/Bbz9VgJl/P6GbSVtqajTmulAHsE0/HfjEBzgINj+wbiHc
3iJURi+UDIIQxAXg53Pyo4CgWrjPDq+5l3BwIACmW6JJaaHS7PAl0xGVp/HpIAMDP1DifV8mG++s
1kK7++cZ1m6otbN9TYNwVVdUp8dnVPNYfAKX8d+BflcWhzNNooPwtqv4kQE94cKtPY07JsBpuCAo
an1gMsLCITp/zyumbDEajwNI96IlOe90uuoXEdeIoO7BmhHhJaf8MksO6p158aRyAiTIs1Ag6zb9
C0Xn/GEqv6NedG5GENhzSPUUh1HBgRiltjOFMx6O4qanx5eBCrOGNZZoJDchwtoud22Rv1FZe+Bo
RPoRicolTDK8TqFL8COGRuGr7/bUs0DmYHLISFRKEccJCuJ50Zck2Z4NwajNre9ZmeMY9wo7K4Vn
c9+svad6iOxyJDKXu/0ZwBf2XB6CJxj4JPtsWO0k9olJyh5+taRr/vsoSTUx+LqmTb9O65MXqo++
MnXEgvm11apxbdFlcCKznJnqMcYT0ljL0Dz99E35V3HCU9Mt9KCd4E3HELKH+PRLgeSKwQEia72V
3hINY+WdnomyssVdqJIaHl4+HcQQynwyIz7paNobp0+cT7SnLe72tPeIYUbyd2tQvHsXCMKIeARJ
8yyO2pM24Ewe4cGV48Jg+84rSWxgRzYhdETH7lrDv7JmyIDrFbGiLxfHMiUgSjjcmuXE0d9qOl5j
1712tOqgRgvu3SQ8btgLS1DcYIdigQgw1zHFnMVgmzjrbLIMSaydmED2uzxYSxcsnIJQ7FhdkMuy
AxLDabZd88vGVmd+LxHTV1qJklT8T7Rze0SIybf950ER4/EcmH6emJ9RTME/tYS0bx+dVJBGnFyG
npedCxmX2RJYiCIhTGCZcOzvKlpAV89RXTFnEeaC74RZY1rAF2TiiERTmgPgvYG3X5JOkwWwFP5o
riolIFNIhCr8LcYhnbRhiN66jBvFKEL2zD+q/wyFyeqJrle+O2uj1MsIBZ40v4jM4Cw+McqZT6Sj
juDjvfoQTT6M4HyaZ9/sTHB+WQ5DpC6UCbUh4bBcGGzoTJ2mj/knbRuGfxbQ0IMjDq9fVl9D7Fm4
TOUNLFlOu2151yF6rF+2emAgqiSKcH2zzjLmoeTPeChE+kL5F7O/B07m/rklVms7SGyOBCrWlZ38
G3hP4/SBs/ib5XMRf0ssTRdFvU8PaGOJPMPCQcmISvjOo0N2YHdn4DRDFqVwA/cS0/fbHf+wFgXM
odbX3R8uaUnnMSZDK5akM1lAbbQCZuVlk6RJFiGL6hGUTcSn19cx+a8ArfV8oUR41bJPngdGesI8
gGfBZlOEwwccNyLztKYBVQc8GKqfvw/U6eduB6hfKVu3DwpCP/MiU0W08QiCscF+1jhCAI2ysLFX
k/fybCdG7p3CW74l8KjMq9V/DxuNw6zeTUZig98c9Pe69X9OOHdHU1/Kg/6seEpML0CTJKZsF5IM
xoA1eog8QqRXNs2rsOOm8DWZjpexKxB9md4WfH0M978dRpyPc1DGkdpzFH/XLgRAlM2lh5hBFULE
ZUwLIlb34CgyZzQKjDwM6ER3dB9+YggCPZ0YCdsG2+AfcunbyIYgwb+3JLlMQKpNrhTgrvfXUUpM
ckSWfCO4G05hL3+s7+X/VTM84tSPZpPA/CLDl2Zh7Vt1vVbYChejnxdNphKf/gJxRUIKDWUmXxja
Sthzfa/CU7Wc6fj2w+4J9pn/LhdaTV0Eb7Go+Ungksin5B9jGEHahfE0lUF7OrPfPfhWVX/tl/wM
MHuydW7/V0L6v8R5/W0x+mnKDEvncVfI2eR0GRXc/7ysvi8Sag8GPckbC4gboMu10wEvhWf2l9P+
o0HPj52sXFXuAxSZFwhtoNgz5dUh0vPIHlyw9+D1AKAMnTZ5cMb+3jZiVunDhgJh0sv12n+aIQya
wKu2iAYP4SzOJhZH4NSIV9cuYxQbkLyoiI9PjZFDG0ufCZEMCrVHPPxS9yBGr8zBoglm0fwhi/iZ
5plMBf58Yb5g06G1kgkXMOL01Gyck9tHvbX26kVKs6K8BZSN92iUYpELASnGJv3vCzoQSbaS7oZG
gQKb0l8ph37RTqHayPnDEm7feAP7wXo2ZYmlXv+3kgIXJl51SeWC6t6mpaASsIL1t0AbFUtpo5i5
MfPeGezdPa++h/VdmVjav3roLFqSmags2mLGS6n74Dy0t76M+yQ2w53RSOcaokrfn+iNZkadE+rw
gVWkVEfjOjR6RJIXN03hhFHWLBR7BAROqw0DL9R2mG+s7KEX2m8yI8g0kSgN2gy9np9/1o7VrBXj
/spi+PipA7NZalgrakShDfRtj8n9gFGnPLx3/GsakHq2hOp4jDJMlh/BqS/vEL0+HEXjDntn/LzX
7RXrSRw/V1w32ne2pB9DHA2/pxuUfcZBFiW+x2UZsy5DB2Tgr1sUXQ77SR5BWXLqk7ahiH82Pqc+
IsRPTb31mF6mCc5vWt58PkXGqOJ6tVzbaVePZGh19vwvsjzt7koYMudZk9DbyWAv7I1bQyWtyzig
JH/A5rR1wQdMQ9vmAyN2kw5UtYbGYmnfmsLqrmRhIsMA0ZuiAe2+IK2E33qTzyMvcn5FIsDLbQuy
YQuCAeKB1TpdqikTOuGXeU98sHJb7u2mz5+bl+XNnheKhEGMYrp79OLS+YhfnaFTpO4ynXwtwFC7
iPnuNqvGqqoAaVEcG/F3h9N2Oxxe5oI+D/+XCTVMBFuT8FZs0cDqHeCmAln/i/kJ4lmlOV+aiMQH
yonyH+/le+LOvXC/xYu/c6k713gz9bm2DTptwABUbmNWhmxPA5GkKvJQ+pXEi/xuDEUg/CjH7Fb4
hNC48vyHzOWTVv8ZN/9acOJBEUeU/rJ7aKtlFnzg+ssun1+PjUAGXfuQvZVFG1lN1aHONEfXoNKa
pBDhThr8l51cFr352YTSXz0vDNfhBxLCs2175IIypvOJjEeEkVKcVtfthEbWO3XajveiFGPbgYzo
vv3TXqtRzo+MAafZcJQVmxk1Tv+mODXfGEj1ZMA4+S4LjMYxprZEQUaJF33Q3LmbFnTSKq5ccZoc
kLMu+/UcYcEoMkzRn1LXA+vQX1wxUXk2jsD3vZeqXqG7eZ3PisEgqLcZCTrMuIDhf+njViNxds7u
eIHsUQrTvpZe0SGKSzGYgIdOMaYJ9zP0urGTmQzfWhLp3giTBXjlXKFCs7PqN7xiXqL+mibBXjXs
FPqjkLonBUeejA/CRhI8ORf640sq82ol29uFBZ9jZ4U+p334i0USaNjz702In9uNVI92G5taY7KD
nAev5+PShvJNFtwDalsSJA39h3V5NLVmeWH7wAN2yBqpALem8yuIJPpQ0OfNlGCQDkjpZhs34ssf
BXbXuYKx7bT4UBuJxKJ+qCNBrrMCZyx1Qz8kilBrst/LkavQH86KCMXypLgXrV3Lt2Kz/2zAtMqf
aH5ipDWVC8uDtsaH2CUB+KCaLEtAkuNtplW8pkIiU91cWb/IdRlO+Yn+LKL7o0BXam4HrBNEn7hM
JbFuwXUYv9+GKHlm/JYNgJJMW6NTq8CWvJis6DVWyDaw1FQkIMxKMHD6zuVt8MJTgHYGXOj5ilMh
aOf6u8rtVAXXTUOdF1+AE6+E1Wi/zGUXBPviPltpFGi88KS/HYnOUR+E/zHtZjScxrfJjpYxk6Et
YRGCQX1KAnhoHvRlGgw7ykt+/BxRYWc8tyv5MudIbvNIVXj3rNzBXttgE4XWsCko4aLtdI516+Nr
yORQSE8bX4eoZ+hzQCGgxJO4pd/MEWPWK5vpcOdWIF15fURFRfaILpOeMUqEPZmEXzAh0QpCaQcQ
Q17sQqWxmt7mz2p4g9enOuxiJD5ZoSh/xW1FeiuI+iGGi3KQmQqh4n/b9uRlnKgUbTiBr5B1ShD0
S9eM1GbKNe2Az4519mEL4QNdgkHZUZpAxnp9l90O2zZirEGtqk6SkU6//wb9ys54fiQVGvey/81p
TT5iwO35w3jA+o9TZCHcU5EX/0C/BdSAzWFO5QtcMXqE/lz9jpPMumqj5JblAiVW0X0ZA78jiWV+
ih5dp1RgacFb8aV9Tk/dME2EFQ1vf7/NJbE/IvQwe5jIYdz4vu6ji6iPRW1gvwjQZUrMWoBMQfvG
6y8wzu4TcIlXdkrm61XlSQeopKDnHzQz9WKpUU0FXJad0k2JEQTlUOHMwH7PaLMfZQY8NE0yGuqL
4uN++bGaJBalEaai2ucT+C+WKBPl1NwFXJ/SgL8MzLUz/aRZgIKFoqwhVEyCAKBADL62SOpMkwtv
/GxiDZj+4qBdYYB2sLow0Y1Hs9r8oG3XwO3d40dT3sK1EaXym46zoyzx4bPEn7nNmc0dB/ThnmBM
bIF06z8C3KEc4u/YXjYDcEiHZAWwqPBKTJCcnyf+ui66RL43xI1alKZBWKFfk04UizhM1hKbp9k0
RfyLvDCbkVQzlj0sQ5VsPP6eOaxCdCPUBaSlHXwvdtK70zrkigNRNQ/AsINM2+f+ychzcSe7liRh
Tb68GELsL3tsAOg0upx0fCH514WOLJd1pSqamAyf5J2jnt9WWJQtiXOF0uyiOfyMjfbdWIJOZbw5
QgZRrl6nKNpQECVh9dGCHmFXtw1eelDvMcOmAB+zYBKps9mkIlWqwtgfmetrx6tUhL6+x0JWQrVr
hPKYaMmZHRwAHmyxAhSZkF7acmtfI/O+c7/tI5qzXhsv7/amSv+Ui5AQ5mC0XIT75zmayWJKrEep
MAGFfGSdXA6jd5WHEnqGnxcZ9Zhl0LLWOyTan5Ak34gLcjmHfrgefqXvivvIzDMzgb8QLUutG2RA
qb2QozKxBw4T+aMeH6ts5ebr/nOWNwJM8RPEbiWQh2ZMHr3tO5G5XMP2uRhyYfeTgFKEgob9YnBm
MESeLGLw/qDqVU1e07+1YCaZl2Mk8fQkkjV3ccWK3BgXjss9CeAJ/O4Ze6tVFJ5c42CKGTEfxhtU
FAerDkQtBgtYwn1rMouoA2BO4lcXhtDi+H0ZmT05dkHSAkVEc5gUhZ2poY4/el2evW3DRYLgaqNq
XUgMqH0znm/tGOHzIUcdvXsOdvE/Q43tWkie1c3nvNRglO7LaRo5S9pHzoaFrz4R/66xfBTQ6KGt
lIHxCRWtdnm1AkREQf0h4gcaa1wcMPe5VtLDbg4eibVwRRwwn5YHhfD2LXQWQdJR+RH83fTGsWo/
BUeNQT/1Im0wEZmgAegnAd3QesTu+AxKewoCoG0+aukkg8+7Oz6sHJTmjVl0PXTcvHuJ+TESZz/7
/XArV1VRNkvbNiJn/EgOm8I8KUOQf+FJWLmjEXfi0uYRvfOieccyIBKoN9reaejBVI5shpKAq3+f
zrskNJ/mUJHlHgo8EOamEaCK/z6D4/CoXWHUZYfBsCQu2pKluZZ9DQew945ebD2qEFynf9YTvhwV
VBgyMXl5XG98BLEY6/J0TX0xNmGdL6+3tsQqnaP+5VG/YZ2PqhUX3z8a2YMQVYrI2sWrIWscvT5e
zIYyoCKDBWErnhYYui6psdS7YMXnLMKoEoZG9PGvGEN4/Bml8JhbbU18jtakgy4kOKhaMX+s3WF4
DoX2oNeQ+nzfMQGQo7t6RmSLHteL1KVHgcfoRtJLEEuMuNdimPga9aOcCj2Y/VkDTWJJw4EvsZSl
Jdiw75kZNMceDNKy2LIPI+Zy9PMz/7bjxO9x9H0gm2LhQNlf9XbxZJQTiE5q6KeeTxEtwymQ9M/C
Th+b9X2G4CZKSBeO9NxefxSEz/MYvruYyHrRnyeJv7cKN3gImLebABMokiNq7To6bDe4Juosg2yC
9g3jUo5r4uc3/qTkMfr/zNdakbKW3Z2ZyCCVZXDvxsnpCnKTBS9BvP+hJAGWxqvB0PjiNVYFtlVb
8cSNLEuu8+trVR+03jff68DlHqBNnZwoIRtzPpYaD2dkpTJdlW7GdQVTcvL+/MpGGuWlt2G+tvKo
ARPoFfGJg1uk41M18WGlcQO0Gp1aD5cRvBZMb2gDeT2mgYL0LsnOE+mU/XITeznRnZyl5SntXXiP
lVh0FgA6Bu/lh9crwkaevzzYs98Hx0jj/N9qq/Q6s810ZKJZoh8DHN+614mgEdWGdevEIJlcMAOe
U/kivPgSmxs5/vP+yN56v/ObifUiIicB8lBOKEp+xep8BNRnOrtTJUzPVpIwmgmCkffKjfCu1d1p
+uiuRlUywlpOHVI45Dd+ShTUbFOhl5q9RslsITBErIdnP3WluE49PXms2Dv3puQ/h7nnjjUeQy17
1aKBDDlwRaAO/e4wsdiBqtUYrjQniVlSH4/jWf46yuPMqHVsGEddseLY2q/QRIPYXCxQIHmIehxe
QlQLsX0nTnvyWuTcLm1ekB8VnORPumkXlflPLKDGmzrrtE70oKk47ztRFVksOWKrqGBKObKMKJlk
ExGaJl1ET+Jj8U0fdi5aEDAPFYGTIHv/nlM5GPJe0pMQ3T9gz2hJ60bbga5nofeWQtPMpvQ4fWrF
DseWFqqHimfFiBI03D+Fieb4s6qUiNHqruLlBxEQyUP06pF+CyOObtI0Nik2C4A4mNE7Z5jGUi4T
ZWIQFBE5WqclWaswAa9nRq4vGkC/lfY2gmTxPqwPF//1vKBbrIOnzoit4KBpm4B9FXOQDwmTq3hG
yTZD5UTYhUzq7jiwFm1vv36LlnXxtGD7nOkupdoNG6etaoT/dkLOY7g7HQOnBglT3lkLaEL87XT+
VGVJKoAP9bVKa1NRVELDI7r+hryPMpBwjOCeuo/e/p8ZaWhGdPOMAUFpeRerZDv2BMSRm8HCUPif
xhu9xsEa90Szz5SlnlMbxGO2CWWsh8Mv5Kp9v8myhxbmICjmp+yfzUwGDsvDVKkx/V4dZVNQvKLF
TRbJEGHcr/oLKpDTJaEqqC5COvFZD2jwq9HWA2M2Yleq6TYa/hhFngYMfd48d01Df1ZElCitZ3Df
1TUQNePhACOiOvdK/FXXeRrkFluqUVYU0hW2+sNlfxVqTLur4+OtaUwZjBoIu6uQCNMwzR6EZFEn
93UgGrnZZKa7Ox/X/yHcn6oc/Y2BisVpfS+DUeVLQxtuw5GUxUqVdE8sUxdmUnDHZFeEHBvTOA4J
yit4mNhF3Nra4VMJCFy3mjvXFsGQszVClgF6upfbLCT3k7P74U3tTCybX3rPFMwo+qV6Bga9nFc9
j4k9LASg1UP8rTKAfPc4aiy8DoGj8S+n1bFDvqZzGbRQksNugKnlnAnzO1qyXEMtEQeizQQOh4HY
zN8Rb1FpiCXDdJGbBnBtgREAPnQf8nGMX0wRUnFNRMQXiyURFOcxxpRx21Sz+Gc4Fsh2DCL8Ux9a
qRtqT75xg8EpK875U1mlzkevQAP5NnA9xhUheL8voKtBXr5oNu8btkfnE8QzY+JzTxxT7NkM6Y6P
9Oz4/i0jMB7+waCf4T6OS4gaRox9m8CSdcW0xgF2siomJUPnJSRooKHAHKWx0v62DMhR3qvMgVEw
I43vJFwzhGCxAPmB4SWnSehJLI6RgnhUuYlt3PwDOKSF8Fs66mQl0kqgRRBy7ssNX4Iw/5yPJZhR
Gmfi+HbrvwoDMmL0ktDTm4CJZo0a2MhM84joZsSZRBZdvbTZ25+Rsu148amOdsReix77LWN/5Rem
/1GShhgYWJgEhHHqTR+FoZzHbA/x982CfpktfWRx8NSA3YUypCV4JEupNXxCfFat8ODIDVdhrR9t
28hi5dp4KoJTr+K1n0uuexnlJ/itCO/l0fXxvPXoxnV02Ihx7AHWPV5pF0BRcOEI7xFAzQ5fJq8t
T0lJYpAFJ8PkSYOgHAxVqWB1g05OzQRp7176Wx+hCl46Pajw9Mk+0nVd3pMQeKmYswJ3CJi3hvMQ
N56z1+ud4CBLvm/fzIUAfe6AJNDCTgVhd3UdscmHP/nBjff8WTM/f5AGC1LNcsCE7/kOhozOEkHM
ZebJP1Ih+iIvImmQiS9XSkwKc/H5v/VQAOT7q5/fA2Ibv+Ho+1S3K7UnHWfChFcILc7Ld248g1/O
qsvlHX1kN5Ce9CaC4DuslfZ7jx/TcKMIQommILF2G/CWx1GvcvUowUyJ0oXbb+phBbIp1CdKz8AA
ZPFyFGowBIRUo8MipmDJO+Rp8FQcA9wimjRaPOBQTstU/2xRg1dXzXdCNqk2VL6Cr+4W+S1Bula0
fbSmx9JvFxeSFFF/zm8vzME0+jouiDHE4etq/ttKYUFef8o03GGcznpg/CurByakmngzL4X2s7F/
Tn+xWzNF6gbMSQyGpr6nvKKgSGEDyd4varfStioEeVlIhTA+iy+ATDBuS6CTunI3khvgzI24r7W6
n9pmIp5FY/sqZocTgQRNGzmhadj0EOf8CNniVyU/Y7NbbtXLD/UMe63f3vgHOm+n4lpm0Fg5uYQu
Nxzjlur8c8KmQ+kpRX4DBC3k8TgOEKJ9kGHZKVJWPm2+U3PJZ2hRfzLvw07Zt+HbU0Z4Ywto3ywi
QUeh+nEUiAvKJAxgybg9Mhc9SVRROrXGAQAniWh8zBhf9EqhtVdnmGkeGKIo21CiA76vAuRzqnkm
GmO/csc7aiKYvKnR7HptW38gCIsB31bogcycP3T14CZB+bBdUElClUkpVgqhAn1kxENplE6H0cLY
Ld2ElK/4CW3UVM9M8D4caPIajnZwDmpsuotyKS8bnPhLZ45L84m08l4yJ+21EHhmFf+E6Dwd+Dl3
GZBFIhCsvVeqapiyMSDxGzNuWNEPyXF3ZX0PhOkwskrlvykb1BEP8Og4T9H3AUfka7qTmvHbtS/I
OvZFtq06uF3VmLKZ6FdWZa0r1sYCOTumpOYUR4zpQPONPe9XbV1yHgoJSWx9Dhto4SeBgCz9vgyK
jOjLqE2uC6+GLD2+oGUBdy8aC34/NIG3sw7SToeIILFWcL/yiGofJP1D+NFZ7Wd5WwkOElKqyb2B
OduI6uYZTUq6WBIaW2E7sBU9fKqnNpr9VsAurgEz+1lIHrD2pPoDpe725ncGTiCY+ISBNzL+31jn
uHFM8/TJCu05Bf9c9PJroMxdlEjNG+TTXnk1j/RU78o9z+9S0JKBiM4H23xbn0v9XGHWkC+lSDbg
xgDzbts7XucbE8XKLg2PmyH+C0FUtvjQ4gaFzU8X3/7v3k3flUC6TweagrZfOVyRqyU/liqAhLez
664Sp+jznGPXppiI83Izpx/Iqoqfk32BBPAFMd0ix5nLuisn9LrVt0+uKeiyJvG5RyvOV6qeXv8G
wxNjl2JjldE8QBBrAQ6gQBMtAmO3f0pErTi8Kgck1OrSfXw1y54yNl8QdfYApW4CO+dhI4sQnZfM
Bkf6DZqZPUVNuKbxGz8K1eZH2D3iSbPfgIeVH9NTY7h0H1FeRa/zeh/4/Jv6z0eUYp4naiMtweN+
MPZ6R+iqgUOAgtS4G3Mqi01cRNDVKD20U6RXObkP8wj2xc7492ZzU3IotLtekaFIEW10tcTf3wuE
MTYxFOUN2vIrGwoDIWc0oku8JzixAChY33zVRlwGpiakVyOA/DdrLZNTVgcGXYpDuQAEAB2xTHIt
ZOxfKr+GFiydZtUFtABybGuPzqSKXbg7yZIolpgAMufDNa04Skoo3haxqmp03HHDhJkIggXpePGe
iBQxxUJ93Y7J7QKa9yDM69pAOEXhvLoHbvYaLSR3m7wZPOS+STqwE/H8rot1+ovoQ+VIM8fKZ0lw
4dtLXb6jLcv3mAWnTLSN+erZJp8UuYp+1hTmNbZv6gnAVw7J9ytLPWMIV9MpidtqYob30QVRGrxH
H9OIcCeICtFOMH72LwsEBGlC1iJZlM4zaY5n9YLwqs/MJz5+YwccvcUR+NdjtLFVevPM2Fm2W5oT
VE/nFOrSfNs20LyYhHGvogGKJDgLhx1aEwe8yajsrNnR2bxrgE02xMD+SV5uwzgsUcPcP61+j3LJ
QVDAYOQO8feiFNggqTu5yxSAV0/U4hYj/0kh9ls2EQy5vMc4MfggoOXwqXYioQQaczlvVhiBbjo/
MU4iPypc1K9AnAVSnnoe/Br2ZOM2KT51fLBVm/7Y1LjpiBecaf+vNOdJ6geCLMXJjKz2oYMpQpmO
V0t8cxYiDdWTGaXXNhWcI5owJxgS5Pj3gBrYICr6aabrCCgcnvaYRfRjQKAP3bPic9VKE2TUcsvJ
/nRjvwAVZ+sL886U4Ab06rIjBxsbpM7YsbuLmT5jeVkoJQ5ljRs+mqQv9bLIufhIUou8NqYSwVwi
Pcl2pSxKv00OeWCrXnVfUuMQIraka7jmjvF6Pl6e+hS9MYdKcxz/U0cEiigHbVsf/5DJBo4FbbUx
vV8nhp0AthcDup4AxcoWJLyTSGt5Xscm3Loj3+WYccHLaPH4/3/0Kg93nUL/WDN107tgciZe2WKn
RCyi81lC6ti2lARb+3ToaqzeL2+ntjB9EIukXK3d6KtCffgSVnkq15gUr31LIh4aBwei0FX6bftc
MBPNdYbm9/eFCVSlHngNS/GDqpViQ6HLIB1E6BBD9TMy0vXAPrmuX5XBEObTuG4N5we39J0QYYJJ
p1suADyGmluTlXowMbhAdB5Lkze5YjdZBofEIRP/UYHTvRjrGdS6dooNYcJDrkvsJ+zRSyqXiFxk
bzlr3W8bOAWxSuSK1HChy+9KSGf82fl5H8yvLmiQUs4fBrSrsuedOXwsfM+pkMpAdaRCtdWREfO/
msQKPscqYmSYEvVyLVgeA5bSRtO/56YWBQHeF2YI2dY8ctV39NKX1VrqcbGcypREJLjA3mYI1fhV
CJmbrgcV99iZz61nPJ1OJ3Qh9hAWXU4icEymnf8jSO4Nijm5rytfFE+aXpRFXnGH8sPhaZuSX+NT
VswjUs0eYrTKMFKLxsxQ1uFZZ//ZzKYpnBA9OHdD5w6LjxbbASuNm3ZpS9kuAagdkA9dfzt+DlxZ
hNIc0RFqrCG77XlFXqm7/jsWJ9dVMgCgqdgJR2MNAQh/SlReEbzxSbjNfdQTwsf1aaby/hRsHC8K
qRvVUfJ5OfGR9n98W0rC3E4csV4aurvLtDVeNPLkVjU5JqJOF4KWt/s2BskhhXUep06Hb7cAYilw
Br/zWR1NEfpCQp0AUjBiRkdJGMNmdZztkTKbPdSe6CP+CdTJDF7Kru+cMC03jAzNuaio+vb7Q2b6
WqGj2N4VnSmuxZwRznJH5XQdfpTUG2N2PJJyUmfFWB6L7M+R6TTq0Uv2//F66b2au6eAgXBZgYVY
q0nWGL3tzyOuNOQ75NAgi53kymOoD2EjQ82MsLtCEjxQCqaY9CNbscyDXcoqMEh9IU2MjUwtGfEV
xo3G5YdnxjfoNn6tHYqiakvPaiwUmBBv2OrcLCJrcjxzrjqWqP7s0S0KPUwp9+Abtmn83NY5wWdm
WJqutRzo+7pWGQbY5fEvcgE6I0sBxh2LMj4LOQqp3nV0oJVkBMcOc9zzq2hWWeH86LyCVfKEFcQH
1QgoIADcmu2HwiR1SHhKlwk+h06wQ9KeKr2Z43tLPyP7pN4rAIv7vTfw/2Cu1I3q72vgggm3OZOf
MQuxZimHng88DRh5MmxkGwcFf9phIf561+iStCxjp4A8SZBo8zSQmixP5ueLvSC/vnbHxKPB3de7
/TzYVZBVrynTX70TQCqSIuZxomNOx0EDYAddjh7vSLVKDbfNyGSWsp8nWM/Dj9MnsFhQTqxQjxX4
80s7b/Hhfu/fstietLZNGR8zARi25TlUB/R8R7zQuugzryMg1WkpfO08Bv3nWKzyAjKnBwHDBdQy
FskZfaNLIhXbwGQbTvL5VDHn+7pnFoa7A0F3rzDCELaLC5xqZOHO760g97ENHMqRkBweJjAlWciR
5NDOluaHX+rnc4CyZQEVdc68DBUMWiiklyaPoHKgda/ZUOCSmwLKoTvdabIAM7aJ4yPh2i/Vw5D9
zSNIDNbx/GhofftkCde2Q9zSEvtopixG6tpLp2dMOnyWcYkqxEaOrRIkz2cVXkEAp14s31CR7hgA
yPc2uHPjk4+dGg8Z83eRvV/CzkSZZPu7AA+9A4ulN24kOMDNvvyZLiqIkkU40IRmy5PPR5UpXzQm
F/Ocwbzlxma40G4KE1vnXVMwyYgWScGEkpJHaIUWTYN4Zs6sm8Ko0ABjXiAVyFU88zOlrMBzCZf1
LSvZk39Ep8KhOaGFEh3DpeRm52W11lJspesi9m+nv5Zq463ZR2/pRkJfPix6aUFOz8qkjKgNNYRC
debxE3196fyGeon10h19xhLE+gQ1jvb8pgXhYFUoGXp3QCiCCSNO2nuk6oOn6tR+88mPzt7OCnFR
+78hTAxUvuSCSZMPr6Y6G5+j589DmoPK730GmGg+hdal0KjnEJPuDRy3AI8QsDIAfOjqGP6bRT8+
Qoyq6GUbd1DEXhF8kE0A6Jr63awaZbOSwFQVqhUoxHvxguw3nhpBghkQgzZBmch/NbTvrYgWSmCP
IU06MaJmn+eZo0/xyK0qv/Ci8DJGs1KHyQfjYGoy0Dv/hVe7soN+/Qdez086KASiF1wKiGiFB8+j
jtx+ABEZo8EcSDP5Q0O5vcPGl2l84WQN7ZUZ81RgrWrFIcszy5eine1DIRHp2r4ZXEyj6G3dwAHI
g++xIAc31CjBwZCozuLm9pVCCjbZcQzvdl/Nsgl8ulWyHQO0PZhekg3N4gUykQKNo8PBcWAFznXl
SePnSLHJCOyfirdIozgutrxAx9e9XZVSWqwoDOLRahSOZlxAxZCSsHnhgfYmBsSMW81fqxPeeEoK
+9cK/iT78S+fJ/HvBJqtZqL8YSBYj2E6/4RPmQ7cfotTS9zH9EchcE/YLVDZtt4QIvHIW0Uh14BK
zirRhXfw5/JGQ/hTNeEI1dozYUfBV3BQTIPiquXvqIez6tfhQpCWePn5d0KP0HMsKAl7hEpviUo3
wHmv9W4zWEDpG64TbDJiZNtGf0+ZzN4vQrNpdSKydEPXeUgDZ2mRZ7ksvgXvZZqVKxpVeLnCmpmD
XkFAGcXWTwkKe3yBYKuNvIyRm9Tauaxo5GC9ptiM1I8qnBmH1rdkaSGT2GvtpD/sI2k77OT0l8aP
zzrKLegRnhgGEfEYIrQA6cFfwZfnSsVSgQLNHQZxQeaZ0UJ6N2YVaMLb0GwGw2Q4LgMLC4Qll5oo
8CgvKO/vzuTUoxGXfVbQQnOhzINoTTO+pwlY6frLwvDduIDMbqHH+6TOJ5I6etDr+fpV0blREptY
a516j72dToKV/nSU+eldDIhs5M2Duktn6OyoXTY2u1JBU1/3RpRhQVplV1IGJnTLoyjQOtMfu+jm
IaThLNo/ruQCBqGPPpiHPrQkVOpn/ffLqM0sdxs6fvpqXRNNIYNqb/dOaQx6vRjO33L0eW/gIj9e
qxtWVDLucu4FTPFQkc6wBp0TY1iN/mFTuWpv70leU2sphVs+diwTRmPdduKyHkipgKuZP6mVSijU
6IxOqOopu43/i63XWKlJX1YxoEHOLs+zILJjcAvDXO2cWgVaDc0Q32myRE0M34DW7h3/b/VE60P9
f7xNDSFf7hEa0AuvkBL8iaLhms5g5/ugtbtFjWRuSeR/GWdhNGcTuEPbdp+2qY3J8F9FSSMK8F30
8gbNMvTUyULXGTRL/1XUy9+ZkKQFkbz14niXJQhIFCV0wuY0+pLoyo4R1Oko3h7le7+LmKFvetsf
ywlp3PPhKwcE5zjKaxTfwdTibiF6tiYkXvhva6+/kVFTKKWCpWduIRRMpm5nuYMhm6e65HuibS7z
/c2KudCObFHuo/0paBaHYvle62+TABrhxCHRxv0F8kLIJMesJzqqBT8bwijKNuGjJxBNVKmVRGmA
GGegnNIltUXwWVnLulqvDvy8V5yzTFegUT8QVJAjf4p917jgfvNbaX6ZDHCSWGZOF/ivpXbUG4xX
4lDK1SQdueg1/GodJJNO3b8EuYtlRnwyJm5lAlr1KQLoLSwrumTfECNWhlqAdWEVg3KdywhONd+6
7kVC5cGiQ1eZOnAdar/NF+O4y5Vh4jhU432G9hGJ8Hw9nu7i9h9pbhv6QqAkYquw9uXYT52OFxRu
cLkRLxPNOzTsA6NtZ6OvdjK6HXuzxSI7WnKnT7lR+Z5KJg3uRII+8QxbCbAEKouXHdMkjc8iNz4p
6gdJn89fz/uMwY3cIX3Wpw7ogCErsBwoceG38bDhLDnca1QarK7iZGZDgPCVKtSQQIBf20cehiTa
d6hkaegFHIfCW1gxA0jH3vYXVzRet/XcCW/pW2sxooKohZ045abgU1eNR4h3Hm/XXITp6RxRMsVN
7AYFo5apld2Rh2zI165lu1kwj6tE02kdGII7iWU/2S1jc3dIYfUHTljuyOIHOn6vVnYZKQYZ5Cxt
vJ2O6Q9ygnnU1KyBLkwYDUlIzbTCl7JjycplsfKeZWcMys/cQiPzHTTgzVis0ZhHV5YkIXsesyTo
N1fU06njW1ElPJJ+NqTCkjOZvczqYo3QQeW1dBCZGEiDYWXwIQPIA7P52+qjFHCcGT7it+Dq4U6U
5SCu3FtWsZ4Ylz70LTxaviu3Sl+sfncOFsKbfgN1eA+6qKsVcvLxhMPNBR7WdPBy2SncOL54WGB8
HiRvH87rmoMPeDjyGvdoTetjSD9D+RQbm7YpS2E6AecvzjNuvXmC6LZteNn4c6Jg06O2OhIdx7uL
7GPIfDALx4Q1R8qciQ0Mlge1mltURJUFkEcH8yzIJkX0mMCA50dtgTin+GQqZ3QuK+hJilJAXe/n
Xm34Qp2CaGE2AasibOyv7IImT7lg9ECfmsDe1kwfuZTQVaEYPO2sKS9Xrf1/SXbb9NUKC00YuAeF
6Zkt5V2bSo+UG+fzO5EXTiOraqin5gG6+X6fBuowQL3orlaelwOrjp33kpHQ+ZaqctiNDJuBk+u7
ftLxkdT6bqmIi8wnC7Y1F+EVQ3Wy0iF8hjLTk1RyJ4Mgx3SxXSTMn0/P9eXiwwMg0EIuz3RGmOtD
UF1XPQ2sRc1MZ87JGIbQI4nizyaQi9AQ2cZFtyKLjU8W5zilESrymKlHCO2qX/kw8UcAIe+zRaYv
QZoT+si3q3oGaHGRNFUzVPP8h1hhY2J5n3WTTUMdSAIFa+XIG+GTKnSb28nozQMKKmKhNADxxpdc
lntxFkg1zOP7iHhULReC+AYe5ak56RBURLlDuXPWWoCWBbzuCOm1pGue/0sjQB7u5stH0/zOk/r0
7YYa14xauOki+v2+C10M2SfxdB7LMYZl+npFI6iSRFV01Vjp9fZsva/00mFslDMHp5dtNCdS7dVw
c9ds6vMsCZ6r4Ow4InGmVUIeGQSph4mTIX4ZgcuRTLnrku0cEMD55WfNlKOeJ5ykAEXQZqKD+6KK
DkEtk84/TWYDmLJSLS5U7W7WShabjGK1shTkQXYWejwCS6AtBk4pN4sPbEJwGe6JwOpe7JiCFpLJ
WaCHGnR4FO9uzSZSio8rE3DLoZSQ+N4BqNeKDc52Dx89n1XchANhznziGmKTjm4+HmTtayRRJMtM
Bh2U22NwmASk5zZXjjwm8s0+VmJg2IlqoXhwtCFCCAaScYBFYeKq8AqGxDbOQaL3mComyXwRr4CI
pJ+QF0M6lVIid5gABbKLTMMNVHMLIJ5j8sTgncMFz/SBZvVGhF+vyA+EAiG7dtDbFOsg4lypkGb4
M/TjzSYjZMbxXFtWEDyIiIJ4ysrNoAVT1V4n+Ulz8KzmIvSc7HfqaIyVa4LZ0W90R3XxMaBJqktH
yzds9eV/j2B6UJisEEY+OUVtIqKZHPXNPjX4I19XME+rtn3wGWNAwVgqAJKFcE5ULPb92y1CGPGb
B+IUBvQ8VPImJnPXr1aw2RuL2u+5unGa3oCAmTykK+Lg/Io9aYNUU2C5pRQGCCX6Hab3eTUi6p7K
hemN8gtNdMhGulXytp7QHoOvjzY32TsFzJhrxx820F0iME67puzmnU0sJYw269A56nmfgJ8hwSEg
87yF64UPL+1tw5J61FRRwov/dcrSrOKbtT7Tmx4SFr06RNuhcdZYV0ZnmooCv31zZOZi02713ep5
qTivOGXAejGLBEGzLUk3cb+HHLLo7nghHFuc4D+PEEvf+qgGXDPDAvjtkEbTc3vewOAbHgSJFn9W
/7mwh/f2auLHhUlpNIR5xSVNe6Ts0esXfiYsUy0Y7soZ5djTsTZoER8Cs5lTS4G7A03BfUtu5Rjh
ixnEkJ/qM1SDf2tUcGg4ki6wBrXYxdUivBWCK6ozAlHcWyVlPA+P6kRre1fj8LLiFncDrRdJhzXp
INIe638MCZ0XOwqVAprZpqdBbMITBTFYNdSDI4iDtq2N8eFh36ts7VRxz2zSgpvuaMZDdM1z8/bn
Ey3nAT+XMDsaLvFLhIbBrgeSiCRsn5Z/vIb7yz2G1yk4T3BQ4jxbRHeUQTKMws8txkUtkRb86wEY
8P/WOEIWR3tMoaeRi+8GhoPljIovcaMa6tzdjlijBYHjQdd4Iy4AxwV+q9FaMqk00ntUSUxmkt0l
PuUiidnHPv4KEqlYrw5vhPeWxdV420yjVV1PyUyQGl2FUgAjF7HDgAWxKctWLHfSMFHIfmjN/v7h
pSsqjR6W3HsaXpCBqKKr9LOG+349ZQFTPnTnXa0vA1ZhWCMUHEcaP4bykfS1dIi0D+5BtjJf2iR6
UmJjAkwk5ubK7hiCnndPn6sE7B0DEloKv1DlN8F7QocKcyyac2hDylEcA4ynuVHAsY1NcMyvA8Rb
IBaOJAuet8gDoB2PnyFD7dfWCBRmwdKhos0PjvEyd399HKz+CrQT2kuz3jfnYF9JOvfsgCt0rXyg
wntwyh/HyyM0/sM+4lV9HCHBNHbfBxsVZo/ck5umsApDPNdYsHEbyf5AMlCWVwp4cDKzlyH1AaI1
kVSQg+lMT0Ade0c9hSw6VRPMYC/+pPajglIFWjvtN/ANYClyNI3PWMTLTiPnSz/iyLt7JG7bCCMM
tScahPiRUYJHRIjA6elFoMVHlpSgyTD6sAKZqyzdaDW/WTY5/0eDohr63u3Hb5sa//DdBytv8ACJ
s3t+j6x0sm4nMiwiuEzbwq46IJj6N/ChnM0AYkip1C4mDwLCS0uQMkktR092P1T7M6UGv9rP6Oo5
PYqR4CaWytiC2n5YYdWrZk0ZyS09Ed4wvwoxInENJr9VasNzIKmmiSytxtslAqRy+6euCiOS3gW+
hiauAXVOn9VV1zFGgNyqjPM7cFCjUGUm5151vMV7Kxum3aAUikqcM8IsAdkr6xWoLkoHWB0bVTKT
xWJB+KjE7jl60WiOU5ePsZBBiIXIG964+gWh5IGNYyQCdrYyeRiHZpGuEW5fOHuM9Cy1zzBbl3Lu
fq8kiluiqsgAe6XSuFxpM/9YTNUQhsR2at7l+VD7eLKo0/GQ0Juk7JBe0DU8JY50BFtdebR/1du6
ywG39CLXRgskSb3Zu8y4KvLRFwQwpLAYzhqd2Ec38Pg5wx1eD241gyu0hfQCWrvBTO2zf8P1G7B1
+OrEstnfJcrfQ52pBsnKNtDY3bTr0SbzPHoInQrWxDveL+jfd83/GeuSmg7KtoKxK7oUARel2/qW
y5nL9MURYgvOZcbsJUH/KzPGKq0WoVDtcU4pKCMh9ei1qyC/BAxCsxzY7P4Gaayuj9beXRKJhkZW
uhJo+LqjQIWPc4NSiCVkmIKpESLQ1t/pBKGhkE/k79VEUcMYMXrUv7ztyemZp79wEpFKpvaN5eXi
HHP0tXT+Ku5cXb5OF1eOz/wUiTOWeIMwzt133ot6W6al7v4CuJxO8VQWBYq6OvtEk8geC8Oh1rJv
YIYy9MNb5LmRhp000AnS4H5AZ/mjtfRnY4zDgCVovkyKAqk0x5n5jO4Stm+5db70iFZ8rROYxD9w
O4YtFQcmQRd6Ge+yM8nMrvJhYpf/83pWZUKvZCcjgj7QHwHRqujWGyv727dUTtmETLz52vMZn/zz
N+N05O/s9hgrig+fObhOaqkXzTgLJVcdGrl2xOJXmw+pE4tGfcMCN3BGpPojqfoMY0jMIbN4AYzU
sI75vPK7ZXKxp5UA12a1JMPERC6jKN9CwOnnKGGQAh1gdf2ZS7XcslVC2bUTPiQI2Le3H4pAcLZd
BDqOF3TOKKu5hPnkViSoV64l4FbSkF0kmbRTvOK4yDTRJwz1cbiDbLN2XWpjQJl/uWrF0+ddmx2m
OZ4o9CYxr6QAnvs7gn/QBv4nh2dqQCIyeK91fiBPvQtfBUmqLm0hatbTC3gJN35wLFtcpp9rcwYw
hdkdweSxqy/D82NwAiSf40uDoH+m7eRrfPiUJfenMildCI53haEacaA0aAPzqrigTo9AUXDyCCDw
fPGZE9nGXoi2ksHzrRRdfK+aVVNS3fn/VrgZe1/dWleN7jzRed0HGwkuN+pGLYcTLfBEhzyRsorw
U5//mo2FVbwJ50c7BsgAyLrEtS5Ni4Rusc2TzaR2fgtVamsg5HFn9U/vxvljKfsHto4eOlvZ3LnO
Kb6YAfzbl/8W8DYb6MLWrQHsPcSWhAH1nXWDezXIa08JOSejOh1uxLS2y/zIY+wyNZdDipW5mL2U
dWccmrmAXhkHBFk0g2EoyEnaS6MYOX6sjcsyFK3nFUqPEloVgJsehyLQp2Q7jGyYxMTF3jaNr5K3
KSAA/zYGsjp9NcLLgFMmqAivwFOfBJ0gucNJYyFPe/7z8jw3NMmOLDEKb9YZEOE+PeSuwTBBHH2R
zehAgPUiZWZ88uvNZFsVdy1GCC7iKr1VUn7O20+N0UTqecsvOhyc9haTR6nA2PShMTZOD8hSAldN
BcuhmfWpoqELNcpwJcGcd6f/6aM+eS15cwiWMwSgOs7AGRw38TQ/TiEUoqpUWEEgULw7n4fKvnT9
dVMuMRl2taGwLMwCGi1k0atDVJ7b8XTex7RuSxOfNIg2Gu7HKFztmIVhV+u6Y83rvt+gIVftJl+I
nFOO8qiLqqRKwzyEN0vApfGgcIeaueqpY8E1XE8MV6Fz5l+tWFaz/OLBOsfen2u/m2zpPmOShaFb
ADe3vBwoxM0Biiq9djbLFi1s2PjRGFBqQJDVXztj0emy+bBzlIJgDQ74BGF3uQ4e5eLOwaFEH6l4
UQ0sV7649SWR8/vYpMGiFNfP4f9bC36/9WGlA4hyoLvMgSzD3/t2ahiE/KIlX+N1yAaUFDh8ZI6z
MGDZLW4jxH2KDAi8+1qUYa4ayz+t69A2FgL1V5pSELVhRQMosAVsHpbBmaMidcEb2HAm2kxdr65A
nIONBn9FBTDm+XqrHZdF7KBUyD8yiF5rQbHwBN8AgDZLz3MQmRYS1fsydiiWXePEwQVd5zhgHyEZ
SdtOEL9uBMwng5kWbUh41FsPb+iFLg7r1bJGmqUIDOHkcsARMwJHgbdaFWXFZrnsOI2VE5mrhgpU
PJpTKYZRzn9NiTOZ48B4Zhwpu6RCKSgdlasTi1vFzu3hoMXwVpVdQGtSMRk6E7WIiykIFUmqCu8p
4bxsGo/8e33IrA+bhxUi7h4Vg2dPk9EcaFmZ2KGJWRcbNYELJrBLc4xVxOIfvl40GL/WdQOhO9ll
MMKSbyMXT7kSpvbbMftcthLHM8R19gZdJVf+PiHuiy/PHP0uuVsxqgaul2GOVZyPK4XY7f0KeCyo
wwvnAm7tjZ4To6K/6pzICCOBdkTaeb9cZKG3syEshVZ9kukWn1VTIgh/Sktd8pLBu5ES22CuWi1D
+/22E8cqIGPx/rbtTwQqpf0Mw8t7Q7fBRcIRgJ/2TFGMJ/Ri4oG6lJvMhXgAJhstVaOpBPmW3aJF
vNFEGqOLEfDJoNBpCJb53wjKkOZLUYIespjmzotR0Gi9d+IzBknP8uaMpWwep+rS8qsOuzPqQJlS
pHAKvUmykmSgt3ZlXjtDrE9UoFBRVNaarPuZs/beMX38Ay4IEw8Ba8K6Yk5MV8+UYro9MnsD7kxs
KVcdju9Ljd8vpHLKmdxXVS2YUO+GLjGBn5D76tqA25tO8XCS5W/rgPsPU+T0b6OO32tavTaEbKn4
e3TS+0lexQAUbMMbExTs2Mbiokt6R6PQTKTrfaetZPIFxYAsJzqrDwfY1RQZiiL1HMpNNTKQchMy
RfRtCOHkfKMfFOSOrx6SfvxFHjJcF3Nb6O1eiX1xModNyBpQLGfQXe9unDyHU1bVJT3qn9V/qMuW
6N2yUTdCQpztwXDQkMdASvHgPDx9F47fvUpynJVd/HPwoYy3PrGqu0N/eN6sgZpFqnRyZAOK5gUw
as8aOYBYwFuea9vrjUHsmcUQLaXJdeLgxhQXD/0/DO/ilPo4bR3EluyfD8cz2WF5nIDBGqV7ygra
BTl+vUr+ByR0ijlhcmMEw56JYfKtdChiVZ6dNQvqau5OPaGqDLgjNXtLFyQnlyKvzE3Gu4XP4+KS
nJS0g99K+Z/Iqz4jptkldQgc4n21EVaEGYG2oUAGg+kHGb7lWAupZW1SF0etj9Brn0KcHWtpfjkO
SPjfDFKg33CAHxei5fcZvFwXp1+FcBy2hdPj4fnCZ/M87Y3oIkzhKaN7bmwSRTFY7XcBzBdB8Bd/
qbvJxQoaImEwQ/7C65pWSIDorbFJQlEEaPctSDdGsHRxWIKwIeAsAiljhEO82S1yeY4EqM0Kilzm
xA2oUUJXwG8wWtlxav36HepgHufpEJ+RAUt89RxVzMbJ4Ma+3HVX+4Fc/c2/WOV35W9UpoTz0EjU
/x0w1RzkKB8XXEi2TYknZSjALs381pyhF1TqC+XiFtpsEjBHbGo7bvv07rw4uEYLBEtG6SRGOHQL
4i18hQMqXo/4+Hu/9RZZK8EvcyCLjVnf+qSyZQMJInazbFU+IP+pyoae9L5GDyR6BIbOJXpOwp9E
TjH9mpmULOsqrWdlS7X83pRitsSawciuxhPe4qIWxvR3epjdKDi9gBrCffuHJUvfU2WrCS9ZUtgR
2Mzi960OmXzImbFKGY7Ocm2NDATERldyquTSTwGMh90yoLzSvzKFpUO+iwv/+6BQYO7Bizqao9N9
UKwEDXL6nJyQhM2N8lehbH8hVRPl6D2hZ6+MCq6ueb7NRUBd98DHI6BlkYE2gsjbMgI3x9BDvX63
Hk8rFuy1nvPoMEaqAtR2KzC55qQ2Qpk60o5kXBMafuv0hs++ucU2TSSomzpIu935YJW02jrje/rm
zolNRLtGTxeObNlMUPuyu9gDzSjn6QGDKuWaafHvHoyaMylVoAU6RJWZKjwsMzMVY0MDmsAXKXlx
rp8o50QXLdvaOPwlDsJBnlPPpfnNa/k0lHZ/CXyy0P5Aob0vaWEtdr810xyZ4Xc+GZ+1vJGcyMcE
fc2rOIs4yywqOqjsKKVrsldJt0KZBgc9odHRrw4wSzJGRkCfW/ed6tg70MfwKMdJxZU9QkvUwYgH
bSDHB+QsjzXmTSJqY9gOMx1tBoGLPTaBv3ydSezVsdMYwdeDeNzWunB5SO65QHNod2idwaOie9uk
J1dss501ddwcMmnS8hqhQ9YrpzkFYpk84+WOUh52FjZTR19BJKcLGP5KSd2McrB92mimghsJ2sHq
2cbjqDiC7fKSvaPg0qU0sJtBIleWOqn9AQe6nr1GUMJOwVKDiIy0aCikqaytu+tPsXfqyhdcIhKh
DzWoqQODZdhoRDrERApifdSUWnviMriix2Lf2sM3PshK1YNgsALXAX2vXJdq503OsIDhoY85ESbm
W+fMwGfATR+MRjfc0D45SMa36VesOAVkljct+mdPAwuC0qGCcg4OA+77n0AxM01TNIcscY6mocD2
9Yiyg/qPFPZIdly0fx0u7ZjzQlkq/Gg2ofq2y5pZhZnKeIU0njp0aGY9K0a4ob+9kf7s7MqzreB9
d+h8rWwtw4obzpY7Axr6gs5yMTgGn+kKZmFkQXRsNa1ToWQyxtvK90oUVLL1B3os5cOlrt37vQ2u
giNk//v26oDZW45X2/d6AC0JlN0Yhhdm3Eh8r1IG4J2BaVOYs0mDxCKHVxdSS1xoqYu8c6+KS8Ei
yycS+kMge/IxF84DdQAmEIOdNa5QXKOg3GeVeRWG7P5iJoqTYUdNeX0+2me8X0WerdLaf7t9rYyK
7MoE2252PXqPMwveeWVSCZ80UVYyr/haQDqfyx9g0u8wd/jBQ2Jqo+f3/lZmelMFpRZ+gMsjFn2Z
sUqNoC0gBApvmUumYn+fYCzS7Jpwu9qYd4mNV0qwPMeOtLosnmn8FuqQTwMzqpD0j5dEylna1SXx
Aqs+QVgiTN+ydCTEtAS0u1OO1mTKu5em2vSMMVO+ARYBjCRpyoq1VOiju26HVM0PwXntLveKl3iG
qLdjr5qO+Y+7Gx8D6w6zQggDTqdwwkyx4d5vypeKjKFJbphyMOhbflpCLvG1eriYOHRF6GWTrxYg
FDT3TTAaVZqUMo81kZPwyQsHj0ufXzV+f4RbjdzlCSYItiOGPDiLed5zyDBpYdI/mVaY6AffbWzF
/cC49rZdSuzVZoQE9yDBa9yeTWFR63F+dlvjF40IzOlo1ryjr4qbcs/UIKfzT5/y2qgJwFLJZc8E
Y74V9Bszm7h6FsnrQsaJFjzYmwCbHi31+Z2nvw8nzV8gAJbdUrQG1hpMj2AH/21EX9xg903I3PjD
1ERJC/wCfBT72Dw5yTZtdsVL8Tesqw4oDRCIW10vLLuBvoPNfHSCGta4cAYP1T5i6Y1L0DShWaub
DzLfnSymHSIPlTAwCHVgOpLeTCxbzguHPVO62Wgpaan/qX9QDl52OF7ydOFtogHKUH9vAMihLcsi
Qprm+lizzGbSN4/4v6d4dFJp0RyGFEWN2PEW6SscSQyMuAWtShjf+TdBZFunQYVOCh9yVH8KbIoF
SAUBMKKAeBR5onJ5JYEBqJoXWTek9EPv9reDtWCm/q84PFmhWOSZVQJZubeK4D0zVDHOSQPNwzJI
b5eUEsOa9A1Yo1Ll7gQcWOkhgBxJ9V4+YEpUNZI1P75U0cfpw3U105KAZKxoxcopntPPZiRhEv79
LyDhaEswXpRdGupKRNN5A2qB0DUzJyi6O+QhH/W+tRm78N7QUZCX8OvPBuKyILYV2rR2Hp1egCOt
DE3P95z+g8nTM5sUoj+n4mQiG1zW8QRiHmjEl5yh+x9tdr+D8/0OoObi/7+oLt0oJbB/2c13OD+k
VlzfxavnhSaSNA8QlYy/3XjyYmB0E8V7C3HejEX0EtB6NggVKXDg45FyY1UxOFklFDCI90kgANIq
K35nBhZe5hE63/RQgJAoaKhiyECirSzyM7yEWzAmO30YSBLOiChRXtBd/05dCnAAgjYqBsN2EJaR
+KXQCP0fVgbyPY+z3r0YENXZAxuca18aUdQ5AXxm0x2sjG6DyW9lQolCDzuPPUMQlWehgMVrgIVX
5ToOV4C5PQcEcxNbay4MCb5Gv8OBbUcL8CUiZJ8IzPRmm2mD2vdSvz/WLbcKLvZlLHtrSINGJu5o
TgTsVTZfj9WU6M8f7KBywk+5pNnotQnorXwla3uOjd+C07zehlOKsCpVUb+clGeGXWAuWX4Fd0SI
8a4H5i/G0zuLGoASaRoWxIgFuCWKKqTJ7/GrTl6hwaeh8KiT+ijQMGsMvnQqmTWuxIAsFs9jW5dv
GSOWBZTUEOgA5hWUkKpDMS6QdVw1GuCZnGP6Q8JPGkVT/IhrJQ81T/H+tTeBChb1S0muPOjGp28x
wzp4SnUcgkSIvdtXYnNAnVdDFvPHMp2bMclZSC/PkrwQIOzwVhTjDoJ6wcSYy7RUNTZr5gfcglwV
G8ySDkpXT+/ntfhnKVhRaZir3y0pi0V490P/mcMIrPp3gy1zlFKdznq9cj4J8GpJhkY/l7G003BR
d6gjCrixo/0cbKFUV0q+qpu+v++5FljmyS4bng2QZE55kuNXooYS9xL2cFJKtDzMAeM37OqehjPk
bz3+pUg9PaMHdxPjouak6mZRKLwfDXOeNKdkyR0+8yfr8BtlpQtj3W9FNk81e+tm6PUpVkN/nw0h
HD8k2ZdY1zN0mpyVM8eQ13cyM5r3ngliLpbh7zcKi5pG4WxbEK8sic/UqbuUjHAjw/CXmTUIcVMe
sFECe8fv/Q7qlUnw+RMgp/N8Q4TJeb6Hs9TJgT0JfF694o8MX4VU1ursoLxB5G+6sHTLl/KRUVax
zr3GV3krlMWIOzIAPAIG4z4D48zHaUEtVCsHEU2BH9V7xlb/iSDAQx+yMHvm1AAsWg1jmbvcvtPu
1sMt7K+y+KydMGAOMjXtz3wtST7EspSYr1yixIt9lwImWoNV65wQRv1hOw5abmCTZIPMcqvANTUE
/cMDi+R86bhyabRgdIAjBT0UA6G5sGrFXg6CtYXnPZEHJ1hRVRXzVacx7CfoHkXQvyh2TkXmEUIU
ZWfiFzYD9VlAY2Jg2WAFeKL26zELSBAZrOYyKMU6oa1OlGoGCX3ZOyYIHrpFPTWd4rF7HoVQNlO/
qsIByq9Mymhp+Oa6yH2aOkra32cNDCVFpwfGnCT7N85kCopYhqX+iSNYbt4uOOD3fzzd0Iu7Kwjy
cFmX7aChFwt1RDtQKAS5oAP2NCH52bCHWyGOufjowkaNRQwK/wPldzdyTjoCU6oC0uU7drV1Osjd
qipe8do2r/Ce34/njcvtXj8Fu86Hjn1ibzoIRyknnspOeWOpuVJFEYiYQDn9AorwqvII4ksZ+N6O
pEbIrsum/5c6rRDosrwTeh8lI7uWJr+X6AN4Ag3/OivICwpvRqR8vogR6dltEv+LJ36TVqoikhqE
xFf0OYZS1mOBfnyvnTF5sbTtvL4mh9SrFIigPzClgNa/VRThJHZrS1JcFi8bkPFSBXrfoBfgy5X+
cT7NRAgjtizWywYVRzKTQ+Q47/pvih1Ac0se3wdzA24ILeADkZzfhBwB5h5bzY4ntZBaIkYtZGXn
jlMBHkngrA7fIYIVUorWjZI4ONNLehjX4my8NVWKkbM9uWUYv0nvgUDK26R2Su+OZTQ9+EBu0VyI
A1B6gpqgPzWN5j+oBVeIbOXYiOolx2tDWTMEABHkEw+sZim2LJlqj2S9Fu2Ndybn2ysOjJyVqNIy
X/v3jf6vH9CZGfOcQWSbSHCrpJ+a6+6/OUbZlYk0bhXbhtlDQXRJd2hKi06CTtcBR2E6n0UYDYHM
LTOwYf6mI0M7EWpl6pbuj4cNW2m8uQbl//vBTXQ5dynAETbln7lCfb0qXsas/pqZaL56IR0rhiOk
UIuR1JBSS2UyW1KhtcK6JvD7f4e5yT57mPrNOu4xCiVBDbRJz/Zhu5V+iX6Z533Muu4R5MDhT4NV
Knr8Lv01lqSYo/6I3GM+V3DmE+4SVR3XbTKfKeQY906FriyRmmfgvoVE2aZcNk6bMWaTzF9YMvQU
2bEpH/lg7Mpwjm1QrShCYyYSCF3lSEB+xYPeWerB+AaruKSAybVoBH4bzILZiuOySNshlMRvI4eV
gHaqW+EvWtNA3dNcGEg3UIjfTbYN7tGZVp0PEN5D0NrramENkxzcpClhflV9b9noY6z+BDEcx2mX
XADrXNX0uK+urvisUyn5mzE7koFSCsBuSrN2P2M3wLvaJ3U7On2NbiffaeQvP4ooiJoIjXtK3C1N
ap7yJIP7Xr+GcFZ88Ds6fiS7euoBKMsi+MDdE8BSKKSFSRJ3AgMtOJz+XfIEOUlA7bNOzz2+4MWF
m6OU89Ud+SaVPeO6O6Q46CzyPr49VFey+xzK/Q82HWO73bQuLanQIMbL9UG2ylIS7OM49QYIA0XZ
gn++mScA26MkmXuBmZ65ZND3dSxhlVnshL5Ve08bSJ+Vhvl6OHRorcUWHr3e2JGx4TCYczP7fXCF
qSvirmVTA2gpIWaO4sVrgUaaPUqB33G+VYMsUu+9Y/zMfxWwC7lL+3oIndsgkFhDmj0BRtFgZnMP
4egQ1CNEZ3rxQQwj85+Ze8VoAorMVw1moTO8ciURQ81bz/4HQuujF/GYxPtGSRGwHtnsotDXu3UT
i/AVI4l37eHW4Csfa0t0CmXVKDw6wc9pfTy2tXwedoErcCf3t7g1Tuy5v7zwNFIdRbLhvY1I1C+L
IaF6XT4ds4Ju836S/W/hZF5H6zbdCiLHFGqqbpJ/nuBxT9wlPaq7e/NuPjaW1JuGLwB36ZfbTgqs
D+GIJnSA11Mseea3Xx5KgkJ0gN10aZ5GxBw5c005uh1NcWCsPjACXic8ZdOX2hY4CQIFq5HTMS80
+uQzz6jKOXLnXvIqipuez2U6yIKIp6v6IW0/HZVnetMQyyOsoGx1fgXZOX/Ce6z5jK3GsauBG8sT
hT6/bA8ifZ81x1S5hIAFkvwYEH/auyO3lwfpFxxFaFlUdw84FGSpdakWBrSV6lCbizDigdHNDlVw
2w6Bayh+3tSwr78D2WRo/TyDRZfqHFdQzpjokrDE984ONVJQXZ8n1MYDlcqvdCa3banyNINvjmc9
8DPOaIw2DDH53GdXNdFAiuJ3e/RFMknXJV4bXOrv0VXgUivlqsWxCeTkeAboGYf28KkP/NtUWKy5
6uBBJ49eTfPqMV+6NyZPXRVMHT8LsJkdbav7B0EkuPqU641FVd8OciNtUIPx0QZuDHT6cY8ryc6u
Be9walTDlB4NAhWHy+CAFrTpAxkfcSwJwS+FDxTFRYH8C0tYNpEww0BwVbbnNUrIl48l8QG5lu/X
2x2I63meIJQVCrSrt2izC7KJjRJfNP+D9EbTsQw9l0Yv0mMirOSOCsNE+P8BuApmr7n1TOUhTmYu
K9LNehW4FoFmZWiripTs9Jtx1pLAHVV9JrQzE8y67XchVOF3l69xDth6ile4vslFfXU/XkF3ysJK
tdji+Hv+qdEYmt90f2S/6GLV2UvMml62+LDdQy3taaUjsMgTfNd4txONE1ZeDApNxTbwUjiVVwrN
2zYZth+4RL1A1F6xkQJCSz4rHS8UIzVOU83t/5i/ETGyyj1+SLDTaImNVy7Qm+ryD5U/leydpbI1
svCYhZGJNFKfxX2WLrWBIJmk3c+XlD9/SWR06ohuek+JXPV6Pp2U4W+nwmoVjJEdbN/7pt9JZjDw
H0dKsO0ZB3lfYGx9x0PFO4ZEt3k6aT0Q0DW9MsZmOZ69OjNvG4+L6gMqKyQ/QEZow9wNK2WUfteN
ou0FGnM4eS8ttBRDVAaZTN6kgPR85VmLZvavagWR+BwkunvI2YMdv94iGKvyvYDHk3TLTQ3Z3F7r
9elZ7yM3WX4iC1OxPQ80z7vFyFiphOlcdLYVahKZw7/wnZhAu0CEyHPPOxGOImFmHJYDsD0aGsg4
K3qlinhMjEb/gMj0b64/dbvGz6wnYZxCy5xtqSF6+tYnbJzlMhelEbEK+L3WXIYgyxghka1zZs5S
PaLgKFW2P4/yLyVOaw2V4I5dBR8ownrU1ixgjyarhpQ14y6Q7b1KHB+QfYyRUZfhC8UT7fkdjz/s
oy870AA/P3HID1HCXFot2DVcpMmLyUFGVbUTxNguszdi/HeVvsxs0qYiRo5H9Rl+tUhe4mRxqLaj
bqs0kwsms71m0rTOybbJCZhfCEVGwRDkI8B0muk0zeQquCLtPyqSIdUoTefxUkg3Mw7mtUJbVXDw
QQ6iXbdtgr5e0wv5d5I8FjaFydkZJzkXbZb318qH/1sUa0YVsx2jC+8HSqRbRH6GZiIWQ9Ak/+vr
dCnQeSxGk4wVceDMrultMR0KeMbqGDLy8LU546IlViS+lN11Eq1cBvCkdA5K0YyaAhPEY1Hfa6dH
YP0SY+JyF21+okAIzQRlrJGNN75raMazdnymGNNB0mjLdCAyyyynEvQ4iFz8UqeRqaMlFnGmYRFV
wqCV1fA2SO4I3mBrkt9DC9OJcm8Ow85v3UdQh3xGntPmaX4QBrx4rdF/szht/9YvFSGL7SkiBAWP
kfS4jDtwW390pF6xtR2ECk4XL0pJgVEQRIKA1UxSV2A4tSSSKSVzcvUnJlcvGiBSGmF/m1CKA9q+
qklC71Q17226CPgYBHuMFasAt1OSPKIwPv4DbaRMMKYSOQeLJktCleRj08OMh5BfPkb+wFhV3s8O
noBBnZFa1eOqSktjGAvTDaUtvS8tr3ufCfhG7f3IWQhI4mBhoBzbNT0U0RgOqtcHWITJ6i/X0del
RBTUvXhpBhShDP33we6OnOEu2E04ihzSddswvz1CxSVhVtGWil39ooyTGZPgq1H4Xqghri3DOuk6
wji2/gy2RktP+KNYJrXxa2/p46BBiI8s4cDCKzMDzBluRctQcrz58K9CQCA1JuTsvsRJVY7gWQlQ
ZxPlyjkthFn/4hQSstSE1F03RKD1yH8YsR7YslgWuNsYG6cKXhhdN2+CoVqt85VM/2CAm2XUiQ6U
acZ8vI2lro684Qhe3waLaN+S8OE1GNgmc50C2J75tQHFQLKKFMerKYH6AmbZfpfJbiSkMwyGTtBG
Rmj6esQ3Cxe+9vC5Yq8bfmJiZAz0M2a5DAzPWWb1eEor+NxM4/MVEn9caegxyw5dm6v3qGLdZkLw
4bsXx+YMUvkeUd92JQR/NhVpHBorSh1hVXm2b482vLXIa6PBKnGNTqNAAn9RV7QLz1sbTykWs0ho
Oq1na3/r8wn7WivyxNra9q9g3mFL4dcuiJZ34RpniD2cgL3VxNRne12NOSfF2SwW16Ewqehm5yqZ
OGdsuwgiAEfScI+Lk1uP0fUs3INjsydZrYwOOHuLNPNbNZU5eamPCBOnk4EP9WEZBLVSDuvisGwR
1agsR1A1mvaKQjHShZT04CTmjvfg6fzc0HVQ3gIAgTBQsMAZ8nieiCSwBSIRIGTr3Vs+3410lH3o
OHjVxhttLXKDravg76YEvRBG9WPIoEmU47Pcz8AQ5Tje6jufq0NxKCqoJjn/YQthN9dwhfsVE9ue
Xc79ey+L2ByV0K5jvW9MZYXZg0k8pFEVQTnUVvMpyhYTAFu+kk64DZ1dBUi3haCM+Ma5zEyk36hp
57wdanLBHCOxqSMS6HN61RH+nN8pesST09vsg8CFZjtkJk+ozaq2iX3aa6mMau5zISP0JyFOHcnH
Tq0J6c454MswTFteDk4WJeOEUC/6jUVMEDucF6aKH5Gql05uYGToeCxK74NU7SW8hFSqjPa91AGY
g+dThB0ypbHkITXKeMCvlP30O7lT5OD+DACx4IjF5zNyvBLRwek3+czDX6NyzEzHLSEVxdNWGK/T
TryFkUh3gpCvUQ8p+9er3pO7+AtbNWgx4EC+mE4cIPYEEd2T9/pmTF2NtAwQNktbEFyI0g+jh+Dg
2Dg4vMc3q2Hx9Z4I9mEYhxX11gs+4mexas1m1+iB/Q98hDlMXp3Twn6Do3tiPflpdo0TT+uCVHz6
YUiGntSHvA3N6YtF0eMRN3BVV/a3b1kaRT43Cnez5yiummyZus/lYuzgfWE4im+XDkCW624yCDG1
PWccN6E9GYZRAxkASj9v7N+v5J5tfEw20oVGdYdHC37i6Bortpfung6+BNp8bZyLCMw27SFU+eLC
XYiel4LKFzwY7RjBiTZ16yXRM+0VCkBTzGLOESTw1d/uoi8M2XWidPRuU80eOCznbI3e1UjCHc7P
QsLNlZGPfiqIjnquT2TJDFFJnTpx8FWhMkGqSWldvh70I7w3dIB6SUgBqIyN7bR1HGHNNhrVVCMc
kghGk+hrDs5zz6V1HkdfiXQxpoWNf4kqRT/e3UXw4UUL37UNfCCcct5XMaltT1HvGIfEXXjFRUVb
O2IRCcCSR9dEc6AK997Q22Y9+SBRBSBYEnyFYuHCHddDpbYQWeEDIV3fUiKU/bIfXpTfGIGeGccY
XF34On3sDw6W3kl8l1FyUQBaruYRP3JGvEjcUZ5OnpiVFxxYXvsL6aYb21eJCqVQKJaZRoCwyVsN
n8o5if8iUDHRCui1c5hzTCcHjIwBxSdU3azSJfAkyeRkvhTg8VBw284P+Rd8eHAKGE7GVrcibeWr
0EtD3jphbjiEYbqSSnU/7bHtGJDQkGADVw2UdGsbVucrIaULLuEZNu083FO9P/gY3zc1u4e0E910
Ygf4twIJKXPZSNLe46BaK1vTCZW6og2jsS+4lsMmNCtMfL2va28Uz0aA40ELT2CxYfwxSQd3Dc1B
cV3XLcn1Ok5EQWLahtryTtM3g+Gl1hu5dxeRj6BqTDfs7+XeW7RIJFexgw6b0L6o4e5ezYURW3Vv
UvcY6sygaXUc7TT/lnzo2m2ZHnzjQ8QL3wBLZ86g54FUqqGRB4dGYGroWlTWb7qc/whKvlZr8+HG
4ITmvq6O/qt3aJ7Vwvq8KGYZpWKm+fOsUmNg0Pu/+MOu53rPSykHLA5EnY/7o4rmHZcEzY4YPlZf
2kTPaAe30oFuhO8iq0I3XI3oE6r/YtGrjkC7AvGsywVdrHSqC55PzgSXDpN/C+oZQldjGMpkesp7
8DOAK/RsaogOAmNRKIerG91cvPEUarEs/Wcq6gMT28ScLZ2CifCzLf/KkCsTjEvk67p/wqO/m6Fd
OD6PxQmFHF3LPgvT6lDMHMIS7g9BIhe2L4nHIa/txzKZV4aa4YlqKzbwc33DQZtiUA8YgWbiawcY
ciI68jpq7jCMtf/YNPIOQL7YcHKTAUCaAavicsokxxy1edexeZFaMWsfPZEld7PfLKGocsiwfQpF
YGztUcB6KGMumxr8pU9L/N/t1zSb+swvfnZiPtX1D4TxF70FBw/NpFkPKvPcu0kKaGoNjynjMFFH
8ebzJnV83Q0vxmKPQGbIj4gYbVvJathtYS5TrerAN4oVJzPlPZG5pADGVja2l15TY+c6CO2Xh3Qx
aq25DVVRNd+/9NQLwtz8ApTRB0rgmtL8P2NVZFNoIQz8rjJFY8OkaJRprmpLP69EtNZd5Anx4Q5f
1OU/N1o7Oi62zNnQBJE5zJ6wBg+mKexfahYFpPJ9E1lKJOzHNnujf4CUjAX3xGMDWpEW/1NGqrIg
JaL6NjJ365uMbA1ueEqciSpe+CS5ROAyuzMt+/Ec7Egy8smpAubuZ5wL80yi6AhClmQlNSpHbOcg
Wka3+L+pWvbW6nTccaKScHfuZndAGopyNKCqaxDdEuQkhw9k2JVcBKYQX/LjWhA44x61zCmNE1j7
cz5RPdR8ayeLNHcFiDIaXAH07eNgkVosqprad2dtCKp4E9b9TiPzeU7Kp3FRkjyoUr7sq0zZez30
iop0DunyEGjVA981TfVQ3LCoTtpJXLiOSKDFxA793t8A/V1Oa0piARb4ccaCS1k3eVyL+i7iwIb+
VlN8Uj1nvT2t9+iRLR1cWRTLvX1K21brr5+ifpwVX+BuuSjzAjJgNR/9ngxa6BFTXwfh4sl0IrB3
pPq6XEzTUaKe7PlSm/Pw7rgocIvE3RGyRi2P8U7vorD1bnsSUAsjxFN/ELeiskqHHG+o5EXqYev/
zu3XHwWJWOC0TnxOVdVIjrFj+RKheeSqg47e31SCG2RgC6thquFioI1F5ILxz1hTF6Mv8xUnImf0
NpXm7DBGFwixt/BGI0fH8OTCg1CObL11axIY7CRY3bOALIbjZ1C3/Uht/guEHcPmeKZXmgryPuQt
yfjkFiTdtT92QVvLI6VaL88C9TJ+cYzuSe6B5VXsbTirL+b+sdVlpWznBpey5XD/tceVUSEz+Bcm
nJuLaEVGvA16BGSfc/3aLoSmdMkTD2RZmvaUVu4omNX93xNY/mp0j1v0qJw9prYWc4ZwN0QWDiQU
ryNz00HDmnpp4B995gDpvu8Ja8U/gkuNRu7bCyWCCy6FZcNRB512q9bjv3APNkRHXbG79yuZloGk
RJWhdv/Nb5JiM1tsWzHcGqYHJ/FqQzQ/w9ci/j5iwtovRYreeajY74WTwlxb4eXfWxLkMKQ3na96
/kp2mrQWpjlr1lPmQOKWjSCRUgerA2aohh953q2zw34+QY3WSbxBDQf718Rgp9wbVzG9r7E5nEYQ
WRyS1qrwRx1ftuUgWsyxMB7TKWlKrV0q9m4nEtAaH5i7lUuqwEaIPJ2YTaVLkqu9jWTy9dDHfLwh
CVfULWY8auOodZBiIT2CAz7a4NRD651GJoG1G6gbBQ4r0XqCv/tREWybCDIYGJ4XUnUU+xDe8cQb
9AvoSQRPHyyGsTXW4zC8w09GABlSwcWwZjmD+u2s0n0Pcwyt4NrOHxOrcScBTPDsLbyMdNOZGUcb
nEcsYsXHP+9oB3KBk6M+dxGzbiwcDFsjCgtOUMTy2MrERovUD4begNUWzIsdafdAnETyDJC9hWbW
bgHc58RuoqSVzxns+zhwTTs8GMObOGD3mZ53LuM0J+ltr3Sr0SCzjv0PJz2ss6CNwyot8/LlkMeJ
HXgWa5EINK+lohxG4UTv46a8XFzwUmEBWcsHkQLrEEEyEmjv91X9CeZacEkgHwx0HrmbcMm/i9xK
uZSGZZLOhUK/CnoY+kH/e9Wi0szXvdkh+iiKWntZd2VtJOUO2cysuRO8mh0326RENfJ+HR555vbQ
3oqcUkZyp7q931xJzh+7oz0QhR/DkAb2Z3whgOMexG8SuxAPbswolPKF0ejHN8KUYhy5a3N85PJp
6wlojGBTmq/j+51HFZ6xQYSAQqwKsSMDYi6ZoyhwBdbmIcSKDifdAOSyMP3/N3ZAALA1YmCcu3G3
99IpNpWXGlwfgsIj13JJeC3SUMpOscQ5SqHeAFGeNX3Cj4gHjvrEX8xptSgHI8XobXHIyucjP+KG
zg2sP8ryptGwD1odfFP7pBIv7fq6iKHQh0jI65KTS3/dklwckOTB7jx9DZ7rKhjQwNwgVRhH8DEP
yDDZxwsYz6dqnoDIrP0RgvToPcDGnC6K1CLKpWSUYglqOhXnm54bVLh5tuLyOitUmSIMjTpDLJom
8QKZCI39EiOVPJtoiTk4wbD94ZXEJ7xmNgLi2gluwjRwvJYuWq72mnI5d5wgvMVyPD732qHccJQn
Y5/BpQh/jZz2tprgeHdIb9Lr21GctlzgzBm5i6WOt+lmHnIFps8aPCOVRlXdqVUnm6sMrPA/rL4Y
SmXAmEOLwISXxMjUOPOqvUJg4mNg5Bv9k6paQRYedTwnl5GDcazDnGKaqGih4d6EhgrTh4fi9u8b
7KymXzdlJxHKrYhnCXYwHzaZLGHvN10WoLCi6fdc9788eCcyvIFVcsWPRS2wNvtQr3u4FJyeg6Cs
fA1txpDFprGc/ZmLZgFCq4PrKODsIyANRBUO5IuDdqIrR6T3FKjh1jdhOxHyeQdgzyyNb307daKK
CLxQLD6dyp4548uK1wZMlaJ/x6MMp6aNK4N3/jW9060MOs+Sb6yqn1NGDCKj0aVl3h/n4H224vBI
5cWTTpT67XMJMpeTgZ7V4ghXFQAnrKLeRgl6YrySc66sGWKejLxEEp98c+4WH/tfn+6QYbRgovaE
9rQ2y47FwrxrX5zxC4EWgv6UDi35fXM9zLyCbow20BG9rlH5MvM1tU54cSXJa93u0MpHkrrQDx1Y
soIXYnla3tVhD++ehGSk+Em2y4+pD9znGV0aNmyjHpw0SWvApoW9s4DF/I2DqdF9+1XkFjl9yP82
0CuUEkoAu8tmyiSAOOzmdW0CCNhfCat1nm0UF9WHTJyxqY8DhFK62cgJE7gCO8In/SKXOe+uY5Wf
ORf/BCFHUzjJVU5pWU5A7AybimOnDVRqT/DjPPJtefHknptrlskWmO8GDwd+8U6NvFAeVJHAPQl3
f3VuHnp0nZA8xQpbmmf4qoOr1wUd/UuCEVpBd6SCS7wCjmPZ7i5iqu+hME5pswETEfCcb2BRCaWR
VN4Bp3jhLSPoeAaLw9xHq+NMvedzrJELSGjFREqqpKfGdr1h8oxJ8ilYxJD4G50femdJZWvkhs60
hyKGTiiYoD6HIxJDqr9uxtUKMvsdrIqCIl9CWY0PA6AA5obqyhGCfSUuUOmVzaE6XVEA1sI5+9RQ
+X1TfJ5jG/SATaIzE9VfOlxZYW6gQsc2qr27jEMerIiAR6633oV0ZfuufrKU4dSagCJrsGIK/OiO
841YPdJzLlYjE7+D5vKw+OkHCJFhuN1GXXUltpRWWCRFTg/FZzOciR6E5eefoL5KwepJVT46TPVp
GrCIHw/W4mpdJT8tc+XGM/4yGyPkOgUVtuaRMaVCKmrHJLPBa286BVhA3tlVAwVMSGtwG2ZucgFM
Ak2JbkmC2DuBGdhdBN71x4yP7rUt88HuSmOkMKVTs3tF1MrXYdkOtMBEvwXirX2SLlMfjWyMSQHZ
hK/NgGL4pO48PJUnfCkbD4fKm9HgHdI66NDjq+bMimXzpW1N1wqUBs8tUM24ny5qd7BvxXGIyyls
nY9Nk7OuxAs0VrmV3tGi8fbujATR50E3JOEN/SXa0/eT0B5yyGoze32zgtalclsJDC0yxMf6UTyP
TZgIKDpqONYTyn/XJPIlP0sOym6WUne59pil9twTvn9VB0Jrdeh6hBHirOE5JUTla4aZcBHpwS+V
2GvOaN74k4Ng3x7bChjPD09M7AFxsXTpTaiJHwRzlK1kSA3B1Id0CwhregCaxKyHJFOMmgSmwBF/
o8Rkl9KZMOoNL263iz0iGtzS728TRR0R+d6xgf0TbY72MOFuvL4Stna/RcMo3EcUUdEGAOySS59K
6Eio5mjw11jBMgqkiWAKzmgrIkv4SQirkixusZ/HsFacmaUuZDImJqMGndTcpco/4g4FRVFhqNWY
IBlNzAHDTbI22p6az1QD+fIHYvI0UcdTUtDHlvgjavCc+1TLAT9UewWxLw0/kHy5JlqbuCdukvKg
9/beLuTX7oJOhqHCqnre0crx2LF3lqolPtTpHBlEaBm0iPXsw2EmoCs5pxCd9O8bkZGLQLmLWMgo
st/buHvPVl8QsLRlSqGPRfN6D40axPmxmkuskZLploA/hNi7t7oo0B5L1nNsA7HJqIMZarl00Igd
L0Qv+HOmNLyqq0fvUSmpw1oNWy9iGtT+UbVNAgOHKK8GdXY1p2eMcaE6flztzO5ehZ2kbDAYwiCY
jrhFomSUEdC7djQ5jmrRQAKRahljPqGNqlj6UBosr8dFkh1NoGuc1HzWsmblJhdHCDZybERvj1bk
UGWd0NT6tjj894hy3VYhKM8Zd0QBIf6ikQ+mux7sTUaPMMI5YBWH1wHyeIprtUSPDUXqKng11z3O
lEExG7m0zvTDcd0Oj1LxlqwplurI+CB6MmAypc2i8z3ob7hbIFI2nEdtGpvoDfAfj6aahYdb1POq
pLm8OP0/lI6bKH/HlYmJBY0sbuLu/vKi/PtIQw7mW/Fptm+JbwJqDctetlQEMA7tWeY8oBXeDz7u
UoFnT2wmHRdd+hObwAuuxKwcHsZfDh6hUqdQH2hex+MtIhHgsAx7Fg/xnjHtLWyxUzrgJ69wkemj
F7idFbvXBD+b/V/dzPwyB9N6dguo06lQtG+qu2VtPxEGwtzVBCfM8W63hft8SASOoK+kBo8Bhnnx
/SpmAGUdtOBao3/CtNX/OBuhAkGf1Ilz6HMI1ZVXsgS2Mw2l22wy+lI4qXOMZqLEvhFQI3uFelCV
V68V4ZtGmpP4Bmc9Jin8bcU7eFfVQWk+wHJTvBEm4NqcdLaY0gynC9Iq+N6tGfrK4ajydNuAfcUX
cyNK6TT01Zu2RHiRqMg1J9PlSqmW2Gn6sOaMs9wU2JTJXfBXEjC1OIHxi0IxiGgd6xQPzudN/cUO
MTwPgD6Q/uUqGDd4owkOyTiAO7fFHKTozGXrkENSbzTjtPN5Z4DzB8xXUKaQi35m419QPo28+rQ7
4KVEhvnJNJCq+f0g4p148rqesrIEK3tcPM9ZE7YkcDHZ1WcrxaeZ8k530HmIt1uKZDVumotrR9vX
YSPgvEWVWOXb9Nnwcq+UqpD/9Sno3ssx1epgxUYhtHvapLh6h/ilBBounEVpscLBFXozLF35SQIR
PVRDWnboG4yONR79d9IjtH7JlaFJ8yxCJvN9HcjMpAtLqZtXhNioRtoYbaHeHfzKqUczQCdU6ZsW
KnB9jq0MmHu+LXT9jNpaM8gGXF0i5RcW8DR0+JqzVded9shUYxu7y+Tt40QwxvO+DfysXop4rtq0
oLiUvNetPanbzTKR5XDp+28Hn33/1+4JjGjlqpR8s9VjEyd9FL6YDmlnd1fs+5bAQVxe2hx3MuKf
PhRZHZIaKZRx27CapSIi+lHbkQmaSpxpJsKfhEI/wQGFAE5AWUEzsRuAO9CtZNDgGrkUIddi2oIq
uRFba8xZ+BFVt1plXdYUZJ12SEtqMaZWGFp+xLIp5JFPYyBuoPGQWR2tu+IKsqDebSu9d/LaM7mr
uSnXl8JUHiEja6Twi8tnodCwNTmuq4nPrH7s+a1xjQqji0ItR1yW/tl/jkHhMXCMrEqZfqWk/7PH
zrq98zB95r/NHaXmuXBNhtLDTE0ewOxc7nXixH0i+6l5R9vgjVtG/3u/DJE+0Ls4Va2W3V1SJCYX
XWB9nLf3v+eteeIreUzoVR5fz/98DLJLGzvzVhvqqMeM5qcRSX8tLrS81RgFz0gy1SEGCGd1UKHD
ybhLXkp7vRVWGTFArOHxdbuq2K9Ve6dywkdr+Ru1p7U2VBg41wGeB2BazdzHOQz5Ow8jw49cv34f
jvmirBt7KAbyOuODgHmYIYrf0Ap6BphZcTLb7r3lCd84vfNJukp1sEH9aMlXFheY0wGyVYzQ+//t
iwllvXBU+NvDMqfKp7fILulkQMlv0JyYPoRoMS6QGT1yrPobRRVl8qgT1m3rPPl1bXzcIGtZyAGP
6RWHa5ay4LWJ5Er0lztCRjFeRyok4TOvQ2sJKk0wqw5nbf1auTxXFLYJ7sXl3IvXg+g8Ft7/bzWd
B/86LebMkSjsLv56oeV7iqv+M3LsEn1eLUTyUF4/l2jA1pIuiWjTg8TVdHvfCxUoEuYmfmAA8qMv
cKC1/FT7MRGDn7LZZh/DdBX7+/r4TkUz96T6a4KQuumfRZQuaejd/B1qUOoRyrezK1ka0ke0D/K1
Fbah9a3+h9iaKLlKZ3zi0VOO+dd6yJX1egn4tMmPXVkpQRJ+5cY1rAVjgjW+czcnC0XqVwzkuwvN
uKq0SfZr21kNBYg9HBPEZ7x+hEFccUzZmB3OWI6CPyfDsCOVYZfLSF2IV5Ns8j69AvFok1Fpuc78
dDOkX0hiJyxQfMLHTAKvofPbApl4QjXFAX41NLU5sxmDj1LuR+cur9uFTyrPKj8fZTuHQzCLHl+t
hJZZkFtxTk9hwmiEtHU9+QHnlCaljAWXreXyOnxKzEp6emkPJi3TZcZA0F0W1u5IbTmNwbuxJDP2
/KF59oMT7+vqCjSRWJwKXc1KzUejevtLvhvLZZAJSP54L8/pu5ZWFJTwWzCSU1G17nJ6NylZSAtR
Gchpe6KJIfUeyKJIEvrcfDYjVQsJ4M3/PD4sFBv0IFB9deMqnWlG7Sggwpe34027uE92Iiwwvhqa
Xk0gkgGcuSl35kcRDpFBzV7HIbA3DMU83FGNkrqTmZgdtOLLvdAifgVI+YXiIY3MypPuc4RD3g2o
24LgXLwSCwytohhgG4jl3rFTG3iShMjXtLTGa3eCPpVcMkYM7sqBqK5iq1WMmYb77kV0V0YObLQX
vWcsbplwFoDVG8JaV2w6ZLSWK6hbXIs0vghU1k3QEzKfnpAJN2gKKmD1OWqaN3EkHB6xy56a2MF4
GQwbf5qAAru30l79g1dnRCBmABjbUE1PS71zWOCK5RzQXhjmLtG5PqRC3ykH+K6X0Ud6xeI9/tUo
1XRGnK9YYnrC0eWqjfp7/DzashDVNIyE+zB8cMbSRtOH3PhxO82TxQ9AKwNx9U1XzAEC2Cr7hKLH
qeVQ94tbQWoA1N4wH7JGxrK9JdKwvNRgmnB1aDWOjRulmbdL7+dN2Ms5wmgKgt5lq4tY+9MUOhjG
at1PrmQ0NHYQYxkfLQ6BvLHKknoOICAgk3YdYQ+ACTOdOaKV/kRM98tUP9nGrpswbdQdaTHwJHga
fWMPEbANJzPLv2yreVIczu4biu8ATJqt0CpnvDpMRj8fzhGFVcc7dcgNJ610shyC6WbGhIoHd9VD
DxvDn8SwIzx8k2fXMXLlhLmzbbBYX0ADZxMj4yXbPYClkR/ruVles6CzykloKYI7sSR8r+ZCXl5s
+2TPFQ1I6FK5kVsAS77STW3WOzr35Na8ANf58ubRQ7C1m1ysZJbwxAJFWbD+FyodV5G3n5vcNmBI
PcC/zTHWzXBVrCbJtatro4UAYTha8fmXrEX3fi4RJ5ooth5O6vPUP0pnBrsWqeFkY4hyd9v5kZSQ
puQVrfRiueQVON0u7CgYExZsaFePvDYmlOwehSrgPjocZcOZ2vGbZM5jnHswNGQYzdXAizZ07D4I
vd3/lN8pNHeDtv7FtpTYIR4sLvIbmv+MpNy8CdnCxleJfFzxQQ6AHmHCN+oZ94tdTcrwDjawmAI5
A9tQJpBX3fZzZAM69/LDJTr7DCKmvtS7384GD0Q1lGkOdUqqRKfUuJ6e17CwThzwNb1k6Dd8Wtoz
a80XM0sCpevSOEtuQeRFziJzMqmvTMAsjQDUVBPErVppJejArh6PxAZYUKASO8b/EnDNnvtL8bHc
bsU9NQtQT5jFUK2P5CIb2Uy03oDH0mexv77hy6s56ulCTAxem83J9iEsKSgUbTp0jqZzYNR1wu9z
l4SOgOGRbfPVNV98eSwgcTvH5qrwLjmW5MgVikYrV8ZVSaWws2u97DldZMnbK4TnYti2vJ04ssJO
Xp1/JlzpDue9t6Y19jvLlAbShxaxkc0O2e2+pY8R1YgE2+v5+EgjQSWreQ9JV/BgUcOhsqPaiH+Y
cUn3pwUOEOQJ083p0zqhy1bzfe4gbkxfeKE4ywOhl4lVtyHIqatm36OEGapdsWHJ7IY+5IAoZEST
w429sFTKgRkgkDgYJSeNsxEhJ87ZVlDloekBrs/roxuAtBGtwLmIZ1D6aXcASo45pJJ+Su2EIZFQ
B1O+Qc4PJq3lX2+Z8N4vP80bjnJOEL01VlyaBp6B8jd6IOw/3HJl0Dy7+GNDLycnN+tJRlmIaPUy
kI8+8yvM+YMbN7EqF2iYUUcu1FkJXr17b4DKWHXsG/sfErR6WvG/S6CBCenxUQZKAfDc1waUedlp
F5rO2VOHjvmGhOLuI6EuV370e5yzMvaYQ1Or+vztixMqqq5pQ/65kkVrsY3H7ZENKuk9tg4fdu/z
T2v6z933awUNwQ/okqVoOKTrgMEVvPqqVaYmTIKFIfpccBOlhjpy3vDzfhvP+HR2guSBt4gysqGJ
pFlGSTHf0CGudvi9/gqEmkGXjH9X7ydTCeWEABqb5LKrPG+37UM0+Ek79lZrbVcEHdvd4gurEXfF
dHBGzIsv8kIBquy/DjwVBsEYj6Qj4UYnsBE/nn1PuxBrC+RUqfxhefKD1ODryET+thW+OG3srH0U
wHKmwzktt2uE54MvabVdaYc6YN2Gj+DgOu1ZbBGCBIGvhChNVP7RHRr3+Qo/XIKodxXdyakwcYe7
t0ubt8NPX0OzE5NcAJe5Rh00xZ3ZffsgYIDzX2+PYMw/Rf81SLYjionTKazfMKKh3GKW9PHM+NCt
pNfb8PXbWHhHnWABfyExBebdja4UgyaxyFS1dRGAqg09XruoPSFgXgPwn5a7fXykgmZzelP/c2dx
HLD8lHB/DweTj+KrRz1lzVoiSQqD2SmTfkHcoxua16BuKORdwip7UyTpk0e7dKL7LwThG0rB5/Pv
ofR/FsgMlyMp0QTCYIzAM50nLwJ/tvSAmCj47QaCgKS5y67UIkFIc/5Xm3/yPURdS++4r+9JFtuH
I26fSTm2YILnxw1RRDkqprf/w9cXMvpt0MGCo5O1BUEg/e7KL9LQ/aYYWr3o0vTN8fvrna4S9s1W
F3B52FW2YAqCjHLQIziCj7qBTj5bSepOdKFYl7WhVAuSaL0ZsbQ8/K1pVQVISHVm09M5lhrqeN5g
ezmbYuS5ge8bn6PlUbURbSzKAioEQA10WKsDSgl/CWsldY1yTskx7AOIzCGCiu7eV/u+jYUG2jlu
qo8MMjKaP9EbWlUzpmXhSMnmSasKjMukK0hqmDtAElXSrSdk3r9Q8BAY/emJjnsBAtRP/eX6vtkR
nXZQ/UE+LVqLZwaI7i6wYTF0a9CMQS+sgmsbPwVfGWZeSMS+Wa2CF/n0WCLK33f6L+x4Se80s/Ra
MJrgwxMthEwLiE2zxtvYkIF9VtqeXPtfLI07Si8L89lvFKziQ/Ui+aF2f/mA7H1DUAuPBDR15vLL
dNmztrrFC6H4wbkoLtAYZhvJm8Rr25dEyRjiqzwLC8GWiXR1DpilHatd71C9+odVHDsS86Q+3j6p
uEB4SZr5JrLNgq6wJHZFeWnLy+ER+UDh+rJYIGZcQB1W8Sv1C5nloakkkvhyWgeE8samw9hS+rQv
9U8aVwFFqTtQ43HNHcTt7cPNLCuONRBxxqzHeVxHGKw4AfuweLQJzp8BcdxFCMYVRO+kjMPUM1Bf
qnxIGZadT9uiNGlpkcKeJ6IHAytysrYgprcuGYGxorSjerMfwwvgh/aGEKNF7y+HAlOUfBg58XQ5
mUZwD7RwbExdfouvTfdrp2P8eE4mlTjplMB50kbHLnk1lN0bzm4uNuanmQNIsYeOcNdBg94joXto
bLzk+wyV5ue1CyUgGhDkfzW8iuiZvPFP3EL2fc8ikPW3JJ2+OUyEEkHMzK6KL+BVWsehByCmmOZK
saKdGELyGHmINxxPPIRr2Ht69/aOqobs7WMhA635Ipa36WsyMkVSz7nogSLDgEmJlO4VnGSCKAsk
94qMvG32kgNY+apcqMJ3l1mqNItjmjkUHDXQ+gS4mdZtrdE4BlYvfWgAwUyU3OZ6VsYtJ9YJd+yB
AUuMKAzMa0d+MBj++/fq2Qsbf2eARyzxpcxcgvt5kgLgk3mf4cHywtXP25g3X+BEUAlOCKxjP0sN
zP1d5KFKe0Q0LP1xFoddehvGR8E0PB66P2Jen4Ys0fidIkKkXnElLizbsBIKUmf5oGVC9L2Gcder
NOggdxb7wpVGrz6MouongD5038GzBMUxpW15ivMalEyDEJFyW3W629cPOzaT9UU874SzTpb3/Rwo
Lf373n3Nd1JpFT96nq5ps3loRWFrl92gAmP9a6l0fk71lcstUEMLG2qcH9zkFal7LyJpZN11ExTl
3UwFzsD3LfbjqdBS2znOOyqRiQD8vujnpPvPCdeMGX+XZmn/4EQNmK9w5fMKUAlDmeonS2cGpKmd
ozT0J6M2H9EQ/j7IfJlPO1yhmb24yMdw0XPylrkZksMUvGrMProN7NnVS8sicKDyUnXgTBpDlVDd
yVU5FAjqOsPDHO6tZF02Cu2k/FmalBUHs1Lr/vOHIahxqH7ML5DO/bIeCWx8TKAbWuQjGXyeYz2o
mHNzusvVshpb2HAXpvqxIq7X2pgdL6NvYjOAoVl341cuEBIzBchhVWQx9rneldMxa2yQXBMKWH9m
6PacAPO6yFM2Aklkq+fltHkqEqqTey1xkSk5D07VyYQXkbImMd9TYx4KusnZv9J9HDjNCW8jRsVX
Iv6yKpoAaMFzdAHpDMfOoS6Uy7VWwpmEdTJuBel4G8/tK4TZZ8TeUWKylFXEhISO8iQnX4t6W1/5
cqvkwkdhW66St7i5lhsQKtmvLNeAVaAk6i6Z8FrFuFzOuAyOP74Sn1yALJCcUfhGff7qKicShm3Y
0tyVwBcKXrU1n5UOTIMG+rWM41GDhg+F13NYfZTFjr5eiAvIcJ9eX8eWO5aA4FM5F1qHQZh5mGP1
qYqV4y7aoRwaHSMIK2EWVkwPJD847sqxnLihmnq4nEqi05Ol1X9I9r8WKSolCiPhq5VXTUuTi/gU
WwaO1ojAbPUIJChixNBGgOXoE878RiGkczYEV/17TfGBZVboEaUAyevQTQRir0GrqoSEkkAfC98t
QlzFOChV8yM1GA+p/8Tiu7T65ciP9YE6j9GwQDeeLAOSi4EJYe9/rdOZPtfgymUYnrRV+KCqMLtG
B+CgoW2DCCT6r0io9P6uP/aK1VVarobVa32CrXNGVFi3X0JulzjKB/qDn5zwXbDx0CzjfEzntA/J
mzi2uCHVXnSvdiS3Bd/czuVN51rzw272FuXHV1wOHlFf8elXwD0fe/XGxSGBe2d+zYDhJM3C2ylb
/1YOLLxc2KIF8kHPCtCfcU4e2H7UJuMpflvA4JKL7UG9Y4hZFuUQiVcY8cp4dsM8kVt16j5wbtzE
wHtWmMHk4951iYmXmgmLnZCXCFe94ZYqpZzn7MzXfto6LqvYYKXvAnbp0QLGdJeg5uNuaDvPhsR0
R19PGiTfyZv1OwVMA5MwWCYmNiLq/4Jflb09ng9chjnj1P6D0VEPvT2Fww4uXUDCaEK9XshEWSEI
Gt5fH7DlZRNQOAnwQZqkCNZOCDlyaGLN0SRakUKvL4t+QRm5lB0fOD5Pd4Oj8LBQnFr9Yz6ZeoQG
YaO9EPKcB08fHdCcNYslEqoGLuFh6zSKi8hRGCkk8a8qdlNU4Qy8KZOkv4GFAeanR4zRoqAfZUlg
mU+YhM2Y86Z1Yi9q0ztJTZnEIBNGl4ckD/GiAB6CxqUFcJd2gngVyV/VVAeo4mQPZduxeile3p8T
vHi9V1o/33BDrvCU3swx/xpJap1NG0hfdUXW8xt14U4IsPi0IQh00BjQ3Fqq5p2AbL4YhX3MZ4nI
zcQ/D2N1xGftgap19rT5lG9JsbDYUwzImA7VQ27ZslLizc59ZTAxPNSz4EK7JClYbvOGDA3p6zZN
gsow1qGoBhqlgVOR5ZSTa4W0UMrDFjxMJL4lmTAJ/Rod+PvBoectUrKK4ocyPxqhCRQfFUNfMNWf
DZnGv6ZwTB2LmAsr/akAgCNvT1YD/4J9IhyBiJcPb9vvJhQMQTrGup4HMV+G5KUqS3j+5PrczgsA
uk3J+tnSj2PPSMRWg35c+R6DLGOSdn9tlbYM9AoymUwKbY+Jn6IycJPS0As7WZ9ioJnJwuKv+ZtS
hQFKiCh3PTdWrNo2nq9jN0CIjBHKM2Ee7Kxne1+322Z9KNUwHKyHuap+a3WuvUA7pakKJNTfYCT9
dKT9wXELj4UDFlYvu20++k5V/1KpoGo1GYPQn8sWmxoL+ULWwoR3t8DjC95p+Rs6I8kQfnsl1MIX
VRqpRuHwHsLBszQBZ9UbucNOPaA158FXeonpwNCSBElXG5P4Qc5nYapniQMaKFyOewm0M2jDVj4e
a0qnxGHxYKJIPAarud9EQeAnPLeqsyGdBhmfIKUbUpuxPDBgcRIK3SN2vt51FyEREyP/qySiPZle
QPTe0dy/sT3R6DOBX2bi71dkprKznYkH+9hlnSut3rzAqhqLrus0GVkunwc5csX5QESrVOxPb0Oa
aTPS6E91mQRA2CRvWT45wXSm2d7Z9ezMFXpGiQzA/Jgt4y1tUnuvs493HZwppYHRi7zdjW823YyD
XzKAncfi60vtqRxtaEJGZQA15cJaayNAlMSpLGxpq6COD7AcMzPN4yGZMJi7Eu+QjPFzjsoTUDXA
nGTK9RKXncZKhx70SoetA/7RKWyDPJsr+T3Bbo+ZGPg5jpN0dVeIC8H2sLADMuRtaQFimAEXv+gj
Uq3JfqBymMulYVupF5ClApoCKMU20C6N/6lRtEZL1qH/HVYaiNcVjzbgPLC0p2TC+txlEc5nm8qy
b1gcPF/DRAWrDTplI9S6NYvQyLywXYcBEB/WhlAUrqVTfiZsekCMAYxT5Y4YOjj7YiQlS4kvfLiJ
1xQvjbPownSXJ+E4XX6LonZqYvOhXsvgKbF2TLHa3vlhbaWInPBEiw8JvBJxIu/DMDg10znPDbzO
8G5121WteiBndPoXX3l6wFmk/HyojbChRfc2NjyGaCsdUhms/Fb+ym2c917I480vasybDipZmj93
0yRWjVPV7GfDD/fqUn+5fFbiMJGhXlFN8/qXIBCI0XhGK0wqiHXWcNDbmHuknaAfv4KXDb+f3hyQ
KN5HqPM83NU3tlQRPjO5lZACK0J2JQ5sw/8zSwTBuTmq7CMBKkQMv+bHaCaBzj5GA3kkmkgf1R/B
D1zRzueHVXAQa+XMwwJySsguhvf2U8lBYlvsEAynnDHDe7HB8ALQ+gDQFLGRG5pty7XcwToSViz3
ZTvcrgf/iXouHXymQTbM0oepuOfewwub02vGTGIR7NvGWdPorjv5fxJE0+GfMH9HBY0xWe2pbrgw
xA6sd0RKcDo0KxNAf1Yi3pgmbFMR67cbNmi0VNKWOYpCy6Wwgp16aGYKFoV83AQ3dlOQuZmc7H5z
eUm7nX0Tpey0O+c2dLFtFp7cb3WBM71HwxwTIJcjB53sI5ABbldYKWkToPJOoDZTi/i/XyFLkYFn
qaaKbAqL+5IWfLmvCgdkR9C5t3Tvbj8OCShQ2Dsmazl185Xg0mVlQsbKbsSsmcP2l48MwiK/IinA
rHxQfIgOXSHGGEfm1qaLgGuLhGSanDQx852C+fbbVcQO+A44gboLxbDg7HU5R3vZGe3niUR0no47
i0W7tUGS7SmsgTYcWLoZG6mCRzhIVLvKI6PKf0NHvxeDSfnkGUhjAI41H4Q3zUe4+7f/CxYOsh9S
zFSCn/Mn8BT8NdfCiNWwbkiNc2Rma0VUNWmZKTvT7wYpqnvVPPmAVt8oIQ5yDS94Yg9HrZt3k645
YLH44XMB8sSgxSuMG2spfJeurDQq3WwHq9u0USzIQU/XicAkQn1AdOWsmv5vdhvtoFJsV1tFHH32
nbJUqRElt5TQXeAXl3y+sSosC7kDMKxJBw+1HDluG5ZzO/rCxhoTyGMzdLKq4/AnyTOueDDUaZ84
6OUJJtUrLxOtSvnXnLYgGZ6XSY1U09vEjKr3rgz+8IvCC0N7oaNNFb7iUf7qYKZaZY6EQdBHBwiu
GPEaLzRJch0nRtiQDDI1YZ6Yx/vWvFKlqdO/l0BmnWlMV1XqOXCH1hxjQheJUNFGHlpySca/uTGZ
KuA+S8zM2wu2MugFDHXCZK+//TidYS/s50Omt/yp+bugX55s7K7wqys7AMfsfb2p9tsPKjSkQEeD
ngYZ+TkJuirud8JjFb5/UHpXn3nvTXJlLQnv7NogDMNQInIDgUpGMXGDnCILqtEL6TFTOMqAnjAO
NTf+5etEJWSmxxucxalcCQAFinsdeQKSwWrJjf/kFBh5eiW90aexuVgG9LeC/duS/YzUC2bN9bgf
OSm9mf5FpwsX1HzR1HkBkSr1tcbiB1711r5Lr7Hf+nj8CEW2GNyu/1kVpuTX6VRHlJelDkSL5SPm
f9jHLy2PaCZOCeVF01PUsmQuc76aok1q/5VjAgGl4/28vUffOwtVdz0N47bO6NE2YEzwRxI6wB7P
n5uS7s6lf5ulQy4YxJBYQCSwKemUabe4F+bLn9YgmYxcAb5QHRh/cwEyGIHDxtY+RfPJ91C0bEkL
lcjHelHyse5t2z2E4eEyuhNUhGZ3H4N1HFaHxk2eBEfoYBPrLSBqp8qI4aU35UfpsNhXuLpZ9EQ5
okesP/JkFW+D7F7siK//UNBVBFKOLeLjd+nQvk3Vwz7xh2taxcunNB6sRbMJ0iwXe/x/qp9OcdhP
pDeL7rgvr3Rs7IP9pY8mJVsYzgnofo/kzYM5e2I2uMOx5DDVT39LVKycjQFDzsoWzMoIucFbIBtZ
d/s+4T73xmkW/cEXX7LBbg0TOCWlurYW4BqXQNkgZWxCDfc15Mww/pe1qqrm1jJ1KUEpMxLp61Gz
OJUkTTOvfvYu+zVcDVHCbrBJ3l/H4mM9reP3Goxxgm0PkXGbERgRWKwgFQW38KV2wFWloXEbQBMV
wrfR7oyRtRdfCe1txSUSAVMw4ApCqHNjE0saj7l9qwP5q9ypjGBoofbrAk5SmtDBa33Np2XvlnmT
L7F1+dvkq3TNAiirmbZ9OIkje8uJhjhBCp712MgfjxCZxc2Q7cZRLxJE+NXJRNO5+qtDsmC1PCif
B0T9poGazxrXOzs9a4HzGmKFyknmsXXxOytbtOOjRHZQxj/wcni69cQIQ4E0fd0nV96JfthT1/A9
TZZKlkj9fIPA6gFadCz7h5rHpqs9ONcascktC4Uv+s5DdSZpnN+gRRkYyk68x7AJ29nTTiD98Uos
j8uB5hZE4H5JzWVOMJ2pohl7R5jr+HVAHsM4fofnoplOnA0Oo5mxaDzJ2PWpoAOAh6mfGnx3NNmB
pl3OAfSQakKoRGHb6aI7JTj297HbbscDQX98y7Ltz1zj5YAD8K+X94IS5QPQWjMVRJT+3RvjS4ny
yO+df8ey86DWIpk5ABP3TvbWUkTSbKXHnQbCo2PztyMgW9mie1VbVImEIhmKqt2EF8JH5HIHLAhA
4JmvUXBkgAOg9A99aXBcVLlbbsjy0g/tvYKhkuFjULPhX2LqGZh3qfb6lMQUh9HviWhY7ofeuKq9
y35ogABcocIl1WTfr4ORpsn3aYkrj9bjpdeJlwlcaPbvKN5reBt+j0+izFjDeZxb+D4QQHfXdlUj
5GinYWnZXdSD24hl/TrbAE/9Kv6A5j7sp4FdJCWsKSFJjbPFQj4HCJybNneIa5yigXrNqqjz+6zk
Nh96VvOYepaysPqI3BR9GJnRqMlhmBFExhS6cJhew1FdBDPA4RxTKzli8gjqZOZEn3mc5NooUvtP
4p+coqsEHxHGiEguXctcgTqFd8Eg/obB8rtM1zuMzKcxwwGKA18JaqS6ZgWRd9gNb/Vk9D0sqv27
ED0lYNKQKRQHQQaE8w+gYu7xnyzPen7LL44hG44CIdONk4stkw+3QbxYsj4fn9imUv7hYPpBMVsJ
Uba5oM5QVxV/usF2EByQABTGX0xZmXiyGI0JSW8hYaUPc0FLfX5Uf4Ru+q1rh9GGQmins6Sv7Wh3
U4SK2JmOJ9F3xF8+xajF2+kLXAt0set8da0jncYk4Vb29p+2sQDX+Y7VAmPpUjqIiCvqdJHbArp3
fQ8JcmC1eHHH7DsZ1BJjHavMJjq1PS9gotnAS65QAsNgM/gl6iBu4ftfqj1KKX0SEOKnYo2UaKHi
Vn+pK0JlWORU5EMOyUbWpAG2SBMN4bXKFVTDDxplIBWK0KXNW6sVIaAFd00h6YVlU7bWYu+ykIrP
f+VjvFregceBVqATXXNKmCqH/+5KYLUdvXcepLGcJ89g+LDctFq1uf7oRBmRiS6dFW5E4JqSYj0H
NbE8+oxFesJftiyYVWH2nQyZraRh/1223Hz3Wk2kW/VUETLkvjWBGdfWQ94WZMerGVS617jQVVIF
VhQwFvj0K+NL269CFSWsR3wOSIjKP1ctRfkXXesqPV2Eue4qlEwrEPhA+AQNLSD3qBR/TycbT8pE
tOhaK/smKpEUWkj/IzlJ8IvoiK6yRD4ogfNnWBddt2mYSL7/mx5Iqur4IUiUCzSvizSSJptYn78d
UFh7WGKAMvrag+Fx2vxoc6AC+s+Yhb1Y8AfTDyE+1UX0nF8avbcw53AQEXdq9QYW2RA6+8q0k6qi
i0yw3RYUwTOdWnYtFkuWtp0hQyQKWY4FXHB+fEOmW3J6EmCOXTIdFbuyNndlGaHsNYOaNNM8XsV0
vx+0jyysoGAFGZrl8YcalnESi7cpvWJy5TU2qwZ6090kZYEVD98OHaqajfPSklvMCPYMNqjuxosM
vL4zlBJ+5CN49LtY1D8kLRTN2RUSDAB4E1RUHyuOC4U7J5edqjSy+wKnwcirg8Sq8ANW1SRxWsP+
DqCeqwEoQtt+3jtoQMkpCEzOPGddp+p+grhSJV2eqNNgwdWBOzs8Wt/C6EsLgUHtNH9X8CQJbspj
I8O1pg7iHBXX5nrVg6+wtlRyLPJt2UN8TV0q2nYrT74JdlKf+p3m0icqJVUyqXMYrXZpI2DkQBcC
0HdHGviGiDb1vdRD6L5Hy4w2iu/tMbIFc7utkakf5/Wq7MRo5ZMU7w0jImAUVX2q282L69l5oFz7
PIS9pyR1hEGZ9AhmNF1oKuyVG/uamMGaGnpyWwjj9iCYJlS2K0iyybAT7emvLMsAHUc37Jr/mS8Q
CxdBo0dyTCpbthS7at9wDbaMXd2s0kqVrd9+mUtagrpAD0VFEJcVkSou9o+nlE93S8MNp/vlrcvl
KoAkl0UGU7FozluD91jCk6uqukgjfCmUmBxam4lzVyQ8G+JfcoPmmn7t5Eqr88DP2Dh6X8eadmER
PFz6vV/uwDrUfFuA4I/F7PmkeVFLLZKeR+hUvHNGKjznXOuQrz31voxthTpL9zm1Qjsj7NMyxAM8
opr69HrW/UGadVP4we6Bw9eSyl7Uc73PEUIFfKyF0eJLX23qED5Ynzj2M05ghKF8QkX1gD3wAw/O
tIDkADhJYZmwMd8VniuzGoNco9MCSfVzgfqw1IYqA2ceRe/cORQXfiNLlnQjLjd599jMp0de8u/X
oxornvGuLWQ74RgEUIOoISoW8SII1vAH7Sa2VimKw/USZzg1apUNn7gaRXO544o2qkAZaKF+4yDT
UadIpVVu9CrDvwIDmezB/igYSbojNjm+sMRYfr+2imUSqORKzxLve3L1aDfpvvDrkyBr80zcm/jC
uzpL3mc6erFdMgphFMYQVxlmDIiCxtM2C9WlPeT6mR/KcNZo9vvu7vZU5vKxm4pz5LAU31oe5O2+
Oim6N7GTxRSwJ6KqcGu5TFOar+6FI5gAfe687zhbNLSXlRO0W9lKNFnNitzrBnvt7fE0D3QRCX4q
+brLWvOFZedmTHAkWCuS1f05s5hjoZawhT6zkhegkY1Icgybs9Cn8wjfT1tozh9ReOXwzU3BuTYn
f7euWpbQIVD84yLkKFB9U4fPahS0vBbePHdkjlitCBavBQI6HjRm6M7Pq4ZXoj9oks7PQJg0ZHvs
37PdxNNty1V4fDffDsPr4Yf7pxscPa6Dmx6vlOJ2nZ3AIUICLuDF/78NwSf7nyjoraordmw9079A
ptTXWgM3BhjZnjVhUzawvSZ5V9GPbuOv6fFLz2T74QPWXqiCiIB/26zj2jzaNpK1wuZqvvUGxo61
iReAtwXFxF4Nfy4vHR1TISV8z3wOSSPAkxQMTteAa2Aj66JefDC72Obvc3aM99GL6a5L0PFO9Y27
v+n+rq90a3S95TXJG2S2Xk+nhoYLn4WxXYV/TpsCNRwQF+rm/9lQdSfYG6RHGYL7dKbFuHhdUHs+
jKyNRZaP5jAgLD55IkpqnNdaIE32yl/qRUkPg0iEiGq+z2ma61cqJL1GhV6sqkuxqMgpIHlb+biI
MlZeLCV5/SEDZQGx3EzXCe7fvAoNDeAg3yha0X5Flus7LuOQUCGvzbhP7Q6b3Bg4HGFmgqcRgY9t
LsNkuKeiQeA633oWjPcoOb63zKRtZpYH2hXJkzaUBuxkZwTify0hkVQAFIFnkdk1BI73nnlK/bSn
O2qC8ZXmREN+PqQNF1Npds0pq4TRgQ3iyj44j/4hfwGBe+hmso5N6tiIV/GPsHBQzfrCVBiw36YT
Wnpz7HkXE2D4NzuhncKq07hKGYlrYYXEdJHXv5QrmwRmt/P4A+nCmORDEd1XjejJ4HYbO0j/L0Ix
39cHun9hygJkGu0BzI2nzwRMBGTF1bz4XASO/2viOpsFTT+ENsX2cQpP0NPFh0n17/8ZHbRXRPcN
X8tiRnRPfTvIRLwA69ttj2HDSsYQsB/fjA+wAYET3j7Fn4Pq8auuENM8Bbrh+1COaIK5wblRNkEa
YEqpLdC8Bsy35zbOSKoOKcdpWZEJPkhi7GDkRPAGEx2V1UtF2fOHvqWrE0Udllf6XhLB9NnbdZHg
vCHB0ljxPzjXwr4RF2ErlTRjKxgV5qgwV+UmFHu7+IMHkQ3xJJks1LAvU6NoFaF2onYSH1mqqO0V
WGMdxb4+tvM9LqKB2kLsCPf49yBnL/xdTLl2i70gLlnapOTVBtB6fuLAFODTLBXB5TD7OFJf52px
B1WG2sssj2siXwoJWpkCQpxPnVhbu2KO8aOf5AsTpUxpas4qvDZDkDvgbAbdqyyyRUEkAzO0ZOJh
tDPQMkOCVroBEnvTyfrXhmK7W8A8+XYqB5ezO0eJDUqYtYS1qSAY66w9bS+51a+2X2JfSakIP58H
PWvI5zyDq75O0lo08tsGQQV2rA9CAKXJSdQEWXYNR5lRAwo1Jw1Q4JTbb8qG78YFfqojmguxPj/T
f/MXLH0IBwTcizAHsBRYNYQlpmsmefH2lUgBMJEYPwiLF3tDCSPZw4Cg2n5vB5FFfy9bcqa0MQPp
cacEgh89Pow15a6r88DXFwuPgGXHTxQ0qj2eNwR7gQowwbxlIBFTwW6TNoqiaGmy7sUAhs0RFBng
2u4815XVIaR2J0vrXSLgGizHo2ImTVjYck1QDI0DTsSmlbF1frqbfc5FEgV/Sm5AhXlURaBUiQ+4
7sWKPeJ+usR5+wiBQ2ATLITl4A87Apl1ye2ziWUcZzSy0jLLyOyV8Z4ReU/H4P9hVJizM/yE/Ft2
EnSG7rf2iaFUuSPSiHNh2KOkTts4s72ckMYG2FitnxUicnQ1IijhWF9M+UHCurXCLDAPaguDPq06
eg2zT5HQveZePck4CJOuzV5xIc+PNcaCY+aDsJTHPOJ1lnDJ1wojS5cAqs1M0G4OHlmOH2nAw360
euWpjgLi3ObMKncCs7JZDBrRh0fBiHVIUG0O6fHdTy2TjCoiAoVv0Rs/t09L+jQ/kgp/sUhAqNgf
4Xc95kznoOstuBXpV0yQrKnlBDu+MZ+SJ3crcx5yy48OhxnPx6MG126wjRt+7UgMHLCsRb2Rh6+B
Tf6kvEh+jB3kgYBUqXe96NRlr/sS1W0pIfamX0UhFZQolLuBlafVgknSSP3nooxziZkX9crWetA4
Rdb9nEOkTdX3FjQAuT+PgiBiG6SlK+o8fnhUEqUSsavL7aJko2eF7CvJGVctOwrI7a7LifFN0caS
BMa2uZT/za6rWg8RhT8LQVJPs4Su6TnyAsH6XDXWKDHVLrIqapKU9TL7Z2S3trsKnDasM6wIuA6l
b2hFtzKyCKDY6B7y3csCrARgJRXfCfnv7iuPloIyzOmUn6MyunNYzxzEzGzisYWVtbg8k1NtNmp0
fTJGNsTfVXeIw7NJkL733XQWG6v+bZYe3i594o3U+guiCGLcJpYZWR6u4oO/jE2NtQMzL+m6Sqb3
fw7fv67o9A7QYI2/GDJAueqO/IClbsAfbI+aEHl2m2+nKpb/ynqzLSRUbfx8UxVzYblffInYCcUc
2Xd95KwZtRWvlgVGqqfz1vPhjpIhZcbycKY/wKOU3Ou79p9OMvtSt5e6UXMK1VppgYKuGK+x8wwh
6gtMDkLXw85DSGS2g4R3qkf+jwhny5gymeG5Uv8PJWsqU/hDEuInka9Dcog7kZ+rFgikLQ8n1ORP
yWSEoJVSRWd4Jw8+8mVP9HkVt9e8o3kn7ELkIwVorFM5DVPwJLzY1zAk9sPrS1YYoG6ZnptOLxtp
lrADLjhIjXmSWEeCHHkw2FbhPlRilvhiSleOnoIbmEoMRS4ifSVvlfmXLV2SOYUPV/shrzdl/jTw
psG/u6sIa9EwDKT7O9UCUDXFG4c85H1SiKegmVmrk9DlQBIhdGtOdOnpSnUT/q271iaMw4d/ky3V
eKIJd59JiCKHaih3L+rdon9/vNEX808vvm6Nq5RJLFaSC9hCXHenRB1MZs/OV6NvUhwIALRC6ETa
KotQpWAwTCa1zPEtheFLbLKh+/jNukNQGucLnZnH79qGE6BmgBqKsyW0srCUH6i7O6FHpF3Zo68N
rhZ108Rb0//vWErcNxpFf+pg7j+LTf1lt0+GyMs+frrizdQWDdwyhpUXLtDF7snw6bzKBIX/WwpG
FiCgcYDgcfxfH/Px52aD7M1b4wFrRCDnMbxQID6qZZ5gPWS6uSrYEX4Uy5s/i5X//Sj8zNRUvtob
byeVN7+3MjYmukLRtHjSkyieC7GUUihODBKB6xYZ2y3YNWp9ZbwGwRvKkA1UGjk0XpTWoMOerFzQ
2VwAmWcvGBnOn0hOQIZeRHfAUzc7u0JlCXRFzfeEBiwO8klLh6FdImWuWsIIvlXv+5gBL1EO9867
YoYLZx4U8/QUHF/nTGarHzY2saw3RH2hlGERf7WjhW4PBwNxUuE5wmBALXbXSzTPwIuYhGJeIbUV
zzRdmNBQngPqaDXCk1eAjkTLaK8o132VLKIXNeT9waY33RwqjPTyZKQU7zEGK10Pj/NYQ8OC4waE
AYKHVfFeHGGk4oRIxpj+p5hmCEmzJJf9Z/2LfbaLYPZwa595we4+FF3fhDhv1rEfGaWzW46uhLLV
nqie5KW0w44eBdaGAYmxRmeH0YRqAYCBcvqQMKpUX9YLalMaMOU4HTKkLRDUU6i/WbII8ucOVqY/
Y8ULh92mKQ92WcHHNeFSJ1D9t4sRouvtTEEYa9vwjz2ZEOQgpzKqF8zBaM9aw6vgnspnC2WGLQud
pc/rnF6uXNQ2rtWsmzPxJCg7dXOB2rCHWgrr5IPe3nF8Y1EhuVfeq9U3FY4u8kKp+VEibxC2mmEy
EZaWIVj6wAm2AJKczcUhMkr7GDRE+LJkKvadqIZYrP42nTGUw4NUYEK8mnR8nr9Zfyf0k2ZrXTQV
Nynjyjzsm6RxaRc9XSmPOcH2yBGiry0mEks/myoi0PIVGhYVxi73JtyzGYT7MRlIZq09VkyU07cV
2XbzFnRWPS9eEKGU402otmyG3Jaad6b5r1gd+2nC3CBVekXcnFvWZbrqX/Crx2drp30fJc9fszo+
junVhJj2t7HD67DhJsPBSmC2SgNaWdlrAyZ01hvLUJnMfFdlPKhSWno5ytzU9Owpav1HIY85+rkw
L2tke9AKJT/trYLzSGOSCWtBVSwnl2yWGLHQAR5WuSMjInn5nbZYT9mPIq2gDuJv+kni4E2m5JsO
OjbyWXXSOHh7vYE2E665EWjPXXG9Tws+C1YrhTbq+bJ3fIRBLZW6DFb8jG0i8ctbipEPuVtbLO8K
OY63ePlO3vZKeJs3f7kD9EBgAfRWw/dX4Byg7zWe5v033tLDslr81qzIVG61axuW+stFAX2P01rm
pEavJyjvlFONm2KAlw8ni00qeVM0car5/5+e7lEFfoUo2XaFeZ3lQSD6brjbu97mD9R0ij+/PPQo
KyFx0I2HFPOpnSYtp9QT8uoUBDYfFqdNI4f2y6K9d/aOQaVAyrg+pn9vqkyI/eV2l1imscIPoGjS
9uxDqi81g6TvfKtXCePOxrHbQSI6XoqaEMwCdp4vUIzKGV6SrcAnhJFxFHRZFa8RmkPEfQrKtpNJ
GT2t0IzTvUSyQO5AgHF3DKM9rdOuZ/oxao1C1LVyx1MnC0v7SQxN2NsfGl1NWAgLLU4lAs2M23pS
SjkWer8oEbRkGmgDUfOPqCFlAVXSm7rON9fzyZRziQ57of9bhenpxcZl8HQTT4h5Wg3zhVSOox1p
xm/c27Bp3BKrZQ7/xCY98GnVtn60IFd5p/+/vLVQyznYHr0u8StOr8o1Xq/hOjkjM3qMm8xJPadm
zi5sBlo7Nbz7ju/bbL4b9zOqVbXQToJa8oSczSfORIlWyvyX+UsZPATA8bNeDsw8+oCX02h17omG
5RSR9hy+crNHJyjHNXZS3iBGD2DJBQJTfyOWqnynKIIkm5qJapuX1MxHx+jrWP1YhurGkPOo0UyJ
CjNziwMAyZ/6k3r7HUuZTnpoVJMgXsNLLc4P8zwlGbJZN6opbx/RndT3mGlvwKncsbJeuigyRv0Y
f2iK5ki+E7WgHjd20wUP0OcpD/4V7jUZ2iIrPblIt1i3ryHt2rPnNp/ChCq/YiOSKzDkRaOJ/vkD
bn0le9f0EtSlZX3K8vAeTLGEzfMV5ODvub83TeqhQ3bR8o9Ayp+OwSOurC7aQ/efZCA9NMNdwfYF
KKj09Kn7Fcybc7dOG6OEv05q6savHc4rnfR/nTiCll5h4JyfTGx/YvMxfcWul3nCYBVipcQFVz8c
jh531T90JQM7H7zf0V30Ro6KCCJuOlgQLfUnGnDTKS1LwWuB2d25Ls1ICWEAyuuKThXwfEuNPhCF
4z8d6GFP4UhjWJJnI4q04N+Vk7sn1HV2wSQ3nSsUvSQTw42Bz9+9uaSXuxp6esGYdF80aBU6JTty
VzI6uUC5szFqvcWBZiYFdHqP4HKsgIrOpHSLtdMm+ogSdhiCzGzTRDF4TBU5/6mza1kPzqzhl7rh
AHwTJcxXcHz7hEY/w2FL7hAvQW5TCmMk3mu2fYggSkWWfPewGRClGCOsCMyklwGNPFeO4/PyPRfX
ShpLhGUC6VAYTyBLGYJq0O0VlXAumBQs+7Jh2sl14KQ3HQLCH7PwoktLOwIfVwKSXM13W3knOBVX
8TvPvery0/98Ui9TCewJVTlQoq7EzjVHDFW2/tRGtCjyJ2ecVkjmGLFHIOPiAWSC09QZBxurXxi5
QGkAwWuyfbBZReRQvb+iN7oTJBXphOua2yGpayY8zTqVWFkGIbcOpRPYV2NWbRdPQ6Nj7vLOTN+x
mEbiCjX2Ph46FEUkk3bX/dd/2dsEN7m2Vkn597Di1oE7N2UzPmAqD9X7sE/rrdosp3bzkc+1bGX0
hE3saB9zq96OO0wxczgKkIIUpHP3FictTni6Ku6nYFcZIyq6BXs8laJFcNph6aNcpfEhscaHUvQJ
fW/QKYhwdvEJ9v1gjJQ1xC6EkvuWBt2D4P82C/aaHHKFR6i1H5BJU+LunvE/pGQ3gzTghuS5lNs/
4e6BUrRs8Pep452+4KaauX5BoehGEgPZIEADLmsDGuhiwwE+ld0wxJL7dDs1bxtDs2XNhpIpSoQd
0bGuZacssmuBzWwY+MiM3yz0MTaOSTyccspRssskvJpxHgmz15RbdyjdMWipbggwehP+/iDWKy6M
lYwVnJi2M1kxN2a6/VrT6aWevXKvuM6Ch5ytErA++cZUOBC1Gh/vgsU0Usfyp7htF6qAvnGbyHXM
OsHOceIOUyGwwmlIqohwCrIA9FDK5mdmQy1kaaRNbCUX89Wo3D17passER1OPxLJ73mG40Lxl/wI
HoE+EwUDhnqCZpZwcSMEEN0PhUhvUr58CLZ+SIqpQd6yy8nh/8mcpcs4xHEtGEkA+fWleC6f0eVb
pVP6VdNB9N2MFscM5GjcXQHoZkd1Mw8bEkz226XFHzxqRUB08PtyQnOvAiWg9kGJVCczii+jcfKg
xtEK3otsg7QBbkPTEhQsgJ7TNqow0vWqKYQ85ZwX+eHckn3PkMqYUPHtSAnzOTzwLk/Q0JQEQsZU
UKXKgyriKCESPaM+J1lu1X5ijPB4/eB3cjFu8nBV6Y/0SDrikgyqNwaJMmWBWI8VKttZ8Exu46oD
0/wwSK7z8iVMAQ8IPfSuSwcyTmKWuyax+VRdvC8rTaRdG+OY6appg5NFWWTxN4JSjRA8NEdbKTCm
0C4CAHfXzNilOr3edfHf36wH0fudqgpAvAuCZKJITDWScHCojPEWLJ3/lFadefsXvfVTR8vfFSI5
To61TiNbKwTL/0w0Qu/FWpDNhuk3QJCCO85/c7C1/5QcYI6MXm+4KVYU7dCJaGtnKaEcb5U+B5y9
R3TcqNTl+yTpbyyw9tyzrXlJ8xbJSNxnXkSJjdjt0lnZY96BNFzCEIywwOSbcvJiYSUq3T3OUrnA
GiRWGdTpBdeW8H2BMqKv8p/SfQQDK6EdF6PxZQp59AUfiFXJwWjMTQxIgGzUMmKYGRmM0yTqEPaJ
i42rlp5Kk+un0RmvrUDdF7VR33pvzV/oFl59V7a1Bmj8qrTgwpfmg70WlP9uZylG1X58k+fZWxEO
2qW+HrqFmgELi/EhmLivr2kCv9nhQiugpP7PZvC8tLsGh0X89XftzeTPy+e0+XjZ917Vff9GA3Ad
ZGKqoa5PGwBrStlLCOHg4VkRxfw+utVbz3BhQ5qTSFI4gHi6sxEJSXs3dkUn5F7YDWeU/mIA+a1k
aPOjTfpyEfHl3LK1C5s0sntW7KBS8McWcQ0jpHPMp1MUZtPxxj6BnwV0BTeEw/M5IUK+z2iWDF7P
l0TIAxEFztQVjmHkt9HboUAt+U+dLtB/bBIvhC/iAjYz04XVzr331ABiZ09SsrvHZo+tNcjM0aiO
IHsbHl349f4faT39p69kwujUsyh2byyvk9poyJgABXt1XR6HcDV7+0L7Lqo0vO04mOz7oNJGB/Db
+jioyQgsomWI4kZWOEp85popsIyXvf4fUQiTtR7B9brwCS+85GRig2DwhYcPYbCiP70HlFMsoMRB
4nyUysQJd0umxh89FdA2jQhUdaLCrMDjTceIx0h6w64C+LIDfewZYiwuqHJt0kivFtzrZu6Bo5Iq
kek3gwH/tJeRE6oEx1JSfxoDxIV5ySblCPJAHlmXfwxRPvt9pOmGm6PRPpm3mGQj+7cehJSmY9Fc
aVN5AsKtQnk/l0SHyxrh0aNFlMJWZ5q0Hop+JQIV29gRbU1M6e4sRgxQKhNrZqtR5TYJ3qA1XDY8
HD8dRJ9URYMVKyOzOJ9D5V6DCLMGjyncuNdWJV5lDXNO5b3Sww9hJCONrPL/E6jDE4aO8ybHwphK
NJ7tdgKAuEbfCGX4b8fuNaEVLx5thNuyQH+OO1FkwV86yM+vp+/lYA5uc61KAJ3zDzmzhYoff6CH
dGUDIBOclz6h8GpcGMSN4GJ9L8pjelYauTYu5M7QuE9dCHe/LyV8WOMl1ynyYVZVNaJIn6npGeXi
T6UF3T5YCAdajIl+T+u4vMrk3O1YFT3ElBbkp8iY7p7KF5NRbToXmSJCxG74K58FKnAdENyUV1cB
lcPm7CrCNm8zWPN7IbdjyimgZPDDi4vvJHs04cWuRce7qUWset0rmy0+mWj3HSPGOk1VXziKaoo6
x8xOAWRuf/wp49L9xtaL006f1oyw/DdBLm55Kx/kmQV7OySYl0gFRr3OIZJ6Am/maIx+0UyyBgGs
QzlFtkc8bsY7V4A6Wb3iVQQ7ae0goPLO+2OwoT+ducbjDuZU/85+b4+K8l/YbsxrHT1DSECzXPpH
1HmrPlaIW2cM/YtQlpCkIkP2OUEWAtagrTDMwU+hL/Fsl9kUbHJaIPfMkSwXuLlbMvWgMlj9RtBH
kIpMOusWVzKz+K91p1/dD9fIhnd4BsMzu4bB1vTOyr9VJI6Pw2DTIci+nvWDK/BmmUmReIExC2uR
uLEjiHLxIkv1dZ0y6//wpTp3slk93RU9mxAMwyYX0cMA9ZH41+9xV9fdIF2uvUf98zeyVxXKF44O
6KoOGutSc/a0RfLObTJHeVOiIPunXkRdCeg0Za9/zfY2/xxUqy08rWotmRKP/1xzRG1v3YWUD0PI
t8xj6+6jyqysD/dwrLg1cBLoRGmlXUF+MFK3B2Lggb9JYryeWDekfwo5jcjzcElesMPrvv5dLF3L
UW48x6gKuc7zc7enaHj7ZRXUBWpT/fihhHHWCCvLI/PHY955cEyxiNsQcSdXNpOZV4BPlenbHruE
EzTLhYSKYsbbfg4I3cbGVih4/yCtpmZ8O7uiKmJjdW24pzNvz4c+fuvmFxFbr2ZmY10ChNE9XlpB
qawDl2fLl0HQC6nmHRi5fCP9jJrRoKd9N8Mx1kZN9V+wakUhYlnQQQPf2V0fDq7L/I6jmhtLJIqS
vHC6Bs0XWlGL9dxrxXiEhhnyJEfrq/HRXLghJB271Qc66WN1yZSxS2dzsKLxObKKklpHb24FCKJ1
v8yYqwQs+Au3vK/QcJkur77GyDtN0EidYUGJ4robmhKOS7YXql+W7kc38fTP+IpIQ8tht8Fc5tDG
TVrSGoMpEB6RnjGynyQ/qEKBTWfTmDQ7f430rwREaul5hAUU9T2G61kSF8JIDGe9+foaa30o4wVb
7UdpIWFj79NQ2mJMta0cT6eow33Knra3XEBl3ZD2PZE1Vjy34IV+W+ZMsspNEUND29RQtvsUxX9Z
PqnUuvVKVxHyM3tXkBse1zv8MoNvseYWPGXYI3ejLu+wxBlqh6/lF0k2lW5VTNyZ3qw3wzlXUfTM
R1Of5uMximSEvnkb5aPNAL50Gy4RRJbWgL0V4T/j/SbqKuuZHwVNhrj3MNsKKMWWW+EdN/SWyew5
5QDphdBG+phstHKCTyyMJ1IT3i/vKsZIk/M50WFLrvfYcnlDm5Bxqeo1b0w3YIDqXvTsKcH23VLI
F+4TAKXtQakp1fBEs8r3v11MA+RrQjgfKMXAXJGlljSOIABUvHXZ70Ni2DDoQg5F8SBT1qu4MYN8
O+yFvLwHDP7CSyFzdZSTIOGA93Ea5rGWSScIxHfXvKac3yswCzpd52ffWuqCMWeulOEE5gq+KpX6
QkEZH6B/srRZoSPgiEdgZQA0b/1CH+Sqq1Z8SL6G+P+kfL+voYIapAeEWci5TJOvggXfpi+wjmFC
MjzaN5VL/YZn1ot//vfOwE65fTAkwCqHu4/OOqRZzgeW0StQU2PkvsSwlNLsqaiJ1JjI0UJ91GVt
OwWbATGFzOQ7Lpb2ZHjgcAoLDvo8SMtLNDi4+B/ua4ssDQ699szAuTHuRVLKYxzOQy/3quAVdLO3
sJJ7eWwHnqsVTouLC8mmfgsg9gsHQ6zBMAm9iAuA66KIN+OjRS5IFG3E6O/UhDSxAUD7K09emi/H
sK3ngTPjJ5PJ3zKbEYbJPszx7tvY3vhGYfVxheucoIhY+FJuOSrITWUkWnYwrzdJYicfi922LeHg
BKZoRsZaUHcdPMog2v0gD9dlg56nnLKSmTFE9fWcFsE/SYdf/LZhZ41AEle4M7W/kv4zZFSW+jRm
nK68QyHjL0rDSOYudvI77P7cF3VzylbOT5aYcTF11xclueUYA2xwx9Zi+XwWVPzDrCnJGgoB6HZy
jWvihWrxpplNQlUFrCMzJLX/8U2N6u2oro5JX6OJ01g0wNVPzmJ2aXOlHIrdqDi483A6J0MVsa7c
e08zWDUAalL6IufcvvhAbONn91NDT7+27e1f76JvbmoxWoc46622zmySfGWFuoyztdi/6LHAiFwX
Y1WYGdWeIbRT6enpumT01yXQr1Lnthbxolu5mDRMzLdds+ip40SreQe02Rz6wH3/BH8f/vi/FCdJ
v8s9gr3aqx34B16v2V1CykYmORh/XTiLDpbi4zeZVu3ZYEIxjoYepil8QdblMo1T+oDU3WyGWyts
giTdsCS4p0grw+N3r5cB6Q0ngXU/yh9gzXk0aHGMc40NIP7GVd0k3Qq4xlfo+r/DIYOszoGE0dgw
wSWSGCB6sGnBIyJmiwxqJsomehrS5KRAm+o83PjsumUYgVA/p0PUVp/f+Y0vBmf2qloJ0ZVcJxB8
mCvPJSyjjBlglHYoE3h5/6J799ZJpSFn2mtSXFm8I5jo8VRN7/9Li9v1F07BKpRfVInifpFdBNr+
/Npw//PyTZKt+QRk0IUYxudbcwxBbFzLB7ge7ton5MNDlmXw2HPA+PfOwzOlTCfukb81DrInbdY3
ufkRnxKOCoRpZyw8KeNKX18Do98Oy6i2z9Zrt2AYYvqw5+G96ESkV2WkY1LEc8tiFSAhYOFUOhQn
OB3OYPvim4VTYX4XJ7RXB/uhqome6sTRzaEv4TN2tv7Eu8K9ZBLdJcrjatuLO9RxLQ/gq1e6yq1R
6afxE9MB5tNX/2OHXKXEe3tt5IBa4yZQS/HdrU+OiEBAQ1NK9iPeLuT+s3VFM6gUP3AA7jcOzbtt
tmNAi0MBwOa9pAaCFRQSqo+L/SxcWgkSHCoQIcZE/fvRPCJJ+Nv/DrH6vytTFZWlKr3WeTeeDJ/6
z8CUgLSuFjjxVC6Ty9moLILlOKyIMj8Qy36PBVTxVk6UCQt+Ec7jw0gprAd1sexMM5hYSua3hgvM
xTCoI347f4Q39dAQYaYiEouVF/LVTvf/9VmsHTmhFJXxlVhnumrGqw+X7z6ziK7nFCnXUQzaIKXu
x7j8sypJ9PDK7skICa+iUz4T0dZPuDKghsse/jmH1roEHF/NoCMwPvkRqky3P4p74TEd+qs2Ze52
t1NGlumlwsqd1kwTeFLcfnKTEWpesHQMXaDwAhto8SpHw80pzAF8MoyWPV99c6sHIhFaoCVHyqoY
iQDLGPgNyk3uljhs/YAYmM8fBBvAtXh2wxTqo1ydZjqX57P9PI9Ai0AEPgyBhuJggNjYBXxiltNi
nmf8bEUdgfLl+CEyNeWURtT2j3giyiyM8uDEIaRWE7LkKIK3ktDqxRFkpKMRBeq1bvqJMghWUqOo
PWWV7F55K/oN4rc4GsWiZEF3lgRUw9wjLrkvsVOl95hd79B4VRs6p99uw8Kv+E+7x/HUU8q2uc5t
75QsJ8l4ZyyoMTBF5x5Xj4d36DhEW5MWgyLBdnK8t2KmJZEw5HSp3TbYSFwR62/nwFgqitNHRP3C
0naEYfZfi7DQm7LJg2yHxYtlUUqjtBKshp6VYdUkXmoemetkzpc8Jq2gD4NKOdJoq3g30bxuVtlK
4EVPZocvzWgbm78Rm6E0Rt+JSigOp6FVIIHuSrc3uRqMLhjh9Z42Ek2/tfuIz4adT8C6ZawlmsUK
MFaZC91REQrC/rzUo9+uT1Kg+Rd/8GMebmqFLzXI1qsUEfDpa8ZHDSQW5ehXQmAJlLaHSiQ1UUfy
/Xio7UboBcAbNZCJczZTaJVQ2H4CO3hxrcucSWT3vz5rcRu3z2zAdQcxrAlJ5xXyZcAtIy2ulX9/
wYl+QHxyoIWqIrb22yoCi8G40CgHt4vsq3qUMDkDzzVhRfQTEUkuoYEcp+4YdEYTkrEloVWgG+hk
4aNgnM3GwRX7+cjJo2NhlJzRXfT/qwz0S7x7e3TOKIhtjFUgf6dvy4UkNSwTprQU9k4dIr8REt0e
LVZSUm8QvSQMtrxpe/UCURNHcyL+gvC1LfX/u37QfzaNp3hqVOvu849zYf5EEekd5B0k1lcTHGvb
7Kzw+aEhnQ8oy/o/V/x2/35lMV9qTtbYMhlvAk8R+Z5CIDslhOm6/8ozgSKK/IGh9UhaqDliOaTA
15GBym6EovB/e0igyiwK6uzOe7b0TaCegdJcCxLm5Kk/bZSRdB+sYxMqOvvpl5BL+gtcqvhnTcfE
k+1a3IHlSG/37kpaly/t4IeIvZotifqi8jkK0eO18AhZsPhp7xYh9QFgcb0jq+1M3mDo3jrL1zMC
GdUXeUAga8vel+JkKyxagdSRMsqjpBxtQFP3smO5546QbFLi6t9TmKI2Fw83MVRtO+XcX5AFnhLJ
mON3hJlBzH152sQ/Z0PH8VTnVr/f79v9GjCDUoex2Z0rTVoDn2D5vX+1AdKi60yODlpk2QRU7p9O
6QZpdT26LiYayI6qEXU+E9IeQNpCi/NzCFhUiEaO9ZdSz7ea8ojLb/3FWLcSFS+tj4ZxW7WNh5Wn
5ir6CioagR/02skrkRMoKCtbUQ/bQZ6h4LqtZ9AgNryXfT3Z8bPOS0WUrUxg3hKEjif5DTAw8XNK
SO8o/N+svoHOiwARrN+ZGvrdBaNfOEd8XENw/fNWlB2AzGA7hkr8+tDsVIybzLsEq7CmKmft/96f
oELPwScSjbJWXJK9GA1G+8Jyjl1qMBBmKkWfM76YTH4pu8QKwE8su2MjzmNvK5b/A5uG1pvLIWEn
JEc1KMxOvUgWK5wHIHlW2CKEJLSr3wmBxeieDeTIU0/O6FnJY+otNGPEQbq81zhtAdVLNfgp23/d
pgVblfPtAPstVB+KWn8+K8k626r643NL0xYUFUwcXVo9VVUILO5VHmdKHBPw7M9k/WHNhuic5ZbX
8tqgqV+XwWe5VGm+kXrbsGH2EtFX18yw7nPKbyFrs25U7yqei8h+X3BmZJ9HSgOXInkGDX1d/gdg
+KRbfNOT/UIegbdux/RR7BGmshevxEhITpJ6F6u19mZCDMLHlBWcPmmixBAJyyVPy6VUQd8Zs15P
DyJ9i1hVkfk+scMJD0q9hJLfspgrzoCf9llVNRjl0NgA2jStFVOjNGO05b8aSitnAH0PBwjG1guR
cTQKfmZIylSHyW1H2Dw6Arjknkh1rH9tXYw+CMM0nv6YaHagaAfRqkS0YD3+oZIU8SreOUD94JhR
E9pSgsYJW1opuntezuE6ot6Oe2VRy7s7WiGZosAiuULPQT35on7H/61HzfJQ7eXOg1jkcfcN7Jhj
lyjFo+5V0+OvlF2f9+WUdnf0DSSJ0fyuO8XkSLd34Ln10M1zmM6sbyvVtQjuG6wL4EgoFDAuEzqo
/EBqfaue9wYspxbgvlqzoKvqweDWMfJ3Q3a70b46IJb89T7YKnXPEQbd4SJEWHPZSH/tsIaQkWfK
IHfI8dFspGK/kSiHjYcEYz1vYjJ11HMYJPaG7IgmVjChQawgQkQnKaftyB7smL1xshnQFO6nrJ//
hw1lSEopXP6yeVbMcfDPiWtutwALuqZ1recKsBhX9r/5iwNE1qXsa8eAyG/q3vXf9gZwERspmrMS
7BINol8yWDVdzYp7ZPxnkF9xpNAbMfhpPCpB/pQdQkqbPVQkSKS6hBS6Fj+ndz4/JV3uhg9dbs6E
7P8ux3l6dXXFsH4ZxRy6rVANcBUkoPxfqFUpJwPhSNZ5RHx1PPIiAPtauRSdysi89DGh7s2jiSP4
+IeD6bWI+QCAoGrgPpL+QfFBhKPtxa42MiTc55t3F+eA7mFHZTMYkahIV3Mk7qSwK5Nzvw3Nvt4e
S+yexeL5mPSP/APAM59IZBHYkg0Wgla2u4fvjI2isLRJcAGV2nwCRCqRA8DJt40rWfsUv0OGh51+
YQ1gG/j6LRN/+w2xGseK94Ny0L7f7ce/2pQohX8y8CIqsnr2fX4a4XgEO6V4n+J/+30aEWplZvH0
thLNJ429L6XkaVrmJ4XfCTkmcw72SuxxB/L/Mqal17P9YFbEE1UuZTHcbZ8fDTvLEGvVl14rWYaD
G5zTVFAnvSfZ6CPwMGehHBf1kRksRppQsVhVGCEaeHzjnVilmDTkW5s79d3CQ9iGqbnls2WSZZgl
j2fspci48lVZVcM9lnoX2yl+auNxX8Gp+Sjb4FKNlY5cBgG0GbwBmPHgef2c97vb9ozIPjLb142M
HRY/EcXOSWHOO1CbGZxSsHlIkP+uSLtb9eTKDgzDmOVQuj4rYk4eG7ErMqdqaiCwHaB7hEtz2WhI
FF00LMtFuO7Qhemcl1xFQWuT6DohV2Aa/jU0VbPX1hFgjbirnNDBYUmosK95c9lqe7lBjdw/5TBd
2GjcNuZWJZP/92fp1g5D1NY+iQIL5+p2syjHfbSAPcEX1Yl6sQNA4sXA9+TU8WFYPW/XQhiAiHsI
N1CjsxMs57dfN8YLUqyU5VnqFbz6naUdl2IHX8ghWRjBy7xctdLkXX/SEeS2UUQjYnGYofve6RSB
tAmaoAlCm/8djTnwtxivbGWvcGdIksA7TG87e0zkAXN2CKJ5MarIKEmRc9bYPI2+IWzDOU5dj+s1
ehTiDeUNE6g1uAjS8VWMxWcanC9vcDCjC4ozQz5o8AcpIDfMJI4e+naUhONJGSt9Mwu1CQ8XBj0N
uXRPRylLvXzz3BPxyiilqhZTP2liCdO8qWk1hsUSN1uIcICkUmECWOOQj5MMkTOljlkoyrCazvVt
xTYhRETKVabTPDQXa8f1cAoYvgu6n84Gg0hh1KO80lJSTw5vJapPntZVdCNSSgQ4MD1ndhed9tCu
5DbiGdaPUyeKM/QLJAsXrbFc8Zr7EhTm5goRQRahfxQWAtr/LKFs4bQdDRCsCTkOeEeQEqeiKjom
vVtkq3xz3uYOSkc80gigtfbIGLVFHB1XC648JpyWJNxvefsa6hhvtikS7+Qife3rruu6EPGc2gGa
eXAVtf58l0/S7XV2kw6TSwPhOeOIERrpaMnO459ZIck5Wgx67q1NQ3mDa5PBWAbdVm3Dq2dYn3a2
XjHlNf9TY4dT1ODAOU3y0Xtt4O6ygMc5pOp9m9COrrWYSrJBX7H8TjL9ZVk1xep/g8WDXk1cpiYc
Iel2L/iLFmm/k3hEKEuiMHLCIqDQZ2ZH4wSSrhn3oB9CB7XQw9qJOGHeE6o4YmsyXbhIriinh2Zn
pKQCbadem8sQB6ysTxbJgmcW++egw+BPRLur8CgwrGxbNf3AO9SR80XDqBRNDdm61r0mdbf/FUpx
Rl4iSpjN4swER+x+wvNCFbFoqwTCO0S/AHZ8Cm2OQJ3ckAmBPhm29IGOp6Te8XS2ivrz4ShWn73v
CSRUI0OWxp2WhAxw35WGSTkoSb/1nOpU5PVPoGSGKGmME1jyl6m2mNGomQRlOXRdAnj/uaO48bJa
sWY6TtCtgGvmObvyYun8H/CDVf8lQpbSol5cO5qYozF4egW2X1VCO76l71ga8XsZEL1OVecBCzxn
KhCgFzpvjFNVkTMdSlfe2dmBzFbFudidVRe5iwfZkHFDF8x1GzwBr2SuDwTVVINo0imggZNdR/Z6
uoRh1z7Vt9z49K9D2POzw8+ZB3Whq7ual2aJp8kRuE/b4zCm6bnXfw4sqOabqiIZ3PhpRqAxOqDI
9YdrYatdlALLlhk18/gCHiHpqCvRBjIzuj03sqaH0TB4S4DgvPh0A2JpPGmSwpmTbe1gFUOogYCc
wk4jM9GLyNqEWKWP0gKTFkxJcMFe04U9VTFUeMjFm9xvqJU+2v8PPKLJSu8Mv6JV+SgDxDuaqhy4
9p8kTABqsxMGWgFXOhDVzyzH3pHf+xuKtlfVBNVpkayxymIaNuvAOxOr1lnhrwoW96TeVbhl53IY
x1+U5SgTap1V3qEEeSZQ3Ao00ci+fh+zY/sG73GiDdY4Om1ANqtARd6x2gbwMR02o3M1qnXklpLP
rccLJHEsCkM1oJPyEBEpupeE7mwZt/d5JwEPeILq00lwueq4wUKFCcoy0KNesD4fivuf5BjSVRVN
IWBHnwReUYFsMWcyvBVUQq1LAWzyUmr/DlbOzkac5hm3ZkHMQFLXk8Y4Gp4XPJDZBMG2nlSWSPbd
Io6Eimos03+cRK2a2Nh3heTsazx84pmfie4wjaXdkNevHJ70nHeuPD86ft6zR5Y+apbcuIvAVPL7
ojN6qxRQ5MIrXf3JeAKkbU6C4C+3B/T5MuhAxHUCBd+Ny22EODAURIpgTyFxeb5JKZHuZS3FR8+B
EyYfEX+IxGpYhytAM28lXFDVt8DJvL2c66RWeFahC00ubo9TE6ShL5Rp8Ve/5NJOzMS4Z50MVkUW
En2caIuDRofe0JrLdPBKexKPyP3xppX74eZZYXPGIWzNqfySdBLqtCp4mmxS9Mjx0wNILk+TWUAl
YMD6/PcCauNvCIzsxWKkotrGTsYZQ0YC1ONmREADyEhopVxpcWBix19H0saMWrEJa5DN2uByK0q2
LQjmfoErT/moN+BKBzWtFT30rd5XjXiFi5yc57x5NxrP8+IV83sonQvmV5gnc3W6it+DuVcvWdmJ
LdjezVEUG2ztc7wPNjnGVySefnOgdTP5hoXZB151diR+TS40v8DzGrHylRXgV8FNW3nU05mMeNSR
1xbwHLG+QaalSSQ9WJGfATRp+IxwrPUTCAMvpyec2uL3wKbLLsLwpb+x6NQ+jB8GzAa4K5cOvVzq
o3sNmNoTqF8yT/0kO2u9heVHF+ufIM2wV8HPiY6+2FWT1CLrCNKM+/OcyovfeiBZ9HeZDspgPuCe
yOt4srO9lZVFKh+NEcZjDV9Ux26BVb6AMqfezkVuDswKTxpYDqRft8tCjxPY37Dl4VEpB/OLYxsJ
h7b6zO91SbWOPp3KbbinHom+Az5HRUCbcxyCexmkqaIXZhlwL4JaJ0VUKK8AwzhacaALB+0L+MYk
7t/mwuMcYiRFuWyprlBEuwK6MK+ZNlDJhZEWMVce4fY23Qna+ovYpAgYb9pqo1ucWsQhX4HEc5Xc
cbiyj31+AtEbu0vlMkqroeQWyl3jXRJu2thYdwjviZ527F7rCYkIL4ynZiscVb4w95Qusow2uMln
TobXXHUopYl1IA86g2WtK+2JjBB8fk2f/ldNNYlenuc0lE4yGqyILnpZDaUiacgbynx6fVU9FwBJ
z6vdFEY+3/+B9iUZ7UO2+k1jEFkTgcodRYmuG6NwXNOrVxPzMCdQS+EmaGBCIdheOD2C4D5pVTVg
sB6QwDVMnyEFJ955Et57I0jhEJ8YjeG4XVx4fxFCbsYvMchvCudo5Msy+JsyRb6PTarg5dL6pKZ3
sE9Mdo+UD3Td8BVZi/+xs39W7MdXYB+ce9EQZUzkrF17mowqSTBSXe9SuWgsDGwjMYkUYIuIfXRQ
MA6D6v/bloatn8uxKgFt4AMXZEC2G42fL6yhXqb6V7zCWnRiEpPeIK/eXnxG/80eivohAC4F5gQg
ut9haumUSvPXrIiMeYQNGgjmDt0CwF7MPP3ZBvo/Qw8049yrRW9Ec4KVnNMbZ3K1371jxwloqe6l
bDC7n8XajIXSiogXIZu2bUZMljX7OAlgwZLa6x7T0PFUeeVUukdtYVL7iLVIBWVDTeYtIqUADLz6
GvlAKAenXxFH58IJpz1ZeInKfcJh/H7RRzLZJ/58Gqmh4cDMkr4beXSkle5fhCRSZ3W8bgrcOrm4
HgiWgUCpTDKjXW+qxg2BHsgiGUMA0g2z+72NJpGKxYMU57TuPIF8LJUCckwcOoQyKTwEjy4QSF2G
20762DwhPv68AXsfuJBlXLWIAFQO+Mx5EmC37piS9GMYO/Dwq7bK8Dl9ClJt0re6akz5EykOy/s9
DarBATXgM9UvBu3EGSJy28utUvvGdwVqXKUocV19dPOTWEBOTbYkqIvOYyONE37k+TqWuQbQOC9/
A10gqkNgbU1RIoUA0VsmyBLgHeeN+TTRx0l1RTy50K9HVyLFxUJuMhm39eoW9lDeUCfswkxhtV3+
62Ot4sq+yT7morxh6LmOgtXKHH4g7Hv5WJmfmiBOsCIwDrd5hV3HLjwPsK7te49axVxtcrTAvpGs
eevAzzG0vvMsSRRyXef/Bbt4sVtgVZXh1oPBcgeDHdOnJ+PCLv9HdquDtu3kAG8ypTJEW2i9K4x+
K2SbTV9EtFZu+g4gq4EcSNx2Qmd19cagKGriYJGvdvcBLY/bOYOeMnucJ+mHUjyeK58IBi2L5Cw0
4lQYvzmVyp15sQCWNrI68iRc381psIS0/+XJ6y963daXEmGqN2+Y3WUB/Gt3Vk/Ah0vJZRoVcZ1Z
zouOY5CH2knoKykygabBmBO/g6Guvs/KY4mO4oWc2dyrJbFypriRNA5N+FJmAm0PzxUxtX0xhY5v
+OhGAMNvBG7J67MsOYPBHBw7rQAL2oDqfM/RIWiZkHAYdkebOqOp3Os6zOKYv3NthUN4y+pSa5VX
l4u/Ql7gd/C0Le0uebOo14kv2ukTfNVjLPL908ijWm8uEzkLRFxu9nDXYfqXOE9/MrhJuzEU7dWn
ggAvEG9nmhKoRDKLv0v2JMG0h3kME92nde/UJH25Z24sAzK6lJZIGyh4/7mUSCplDHhUB+4Qxc7E
kqXEAnpXGioJvyYgR2o6JASr7ingbUSVDpJSyn5vL8hUXypiI2wcnizx/1n5+Y3CQEcbH8ju9FYq
A5vUDqVx04A2RzdMjV8cVa1+4zp/Tl6+xVa0mplzeP9ylh/IXeqzxMbbWK13H4znvd/YR433Mybp
O5KLd1tnWnmqgndE8s3OZXx+rhyqSa6HJWsN6VG0CBzeR3fdNYz0WtO2fG0Bofkc92hiMkyP92bH
0oc+3kzhEXP2iWbvckiFGYuPw3IffKz2eDdhcFcaayUK3nsUhIt5ABjVttjtuMSWo49K6ANaNsfC
x9PNUaOIXmeeNOuVpY+zXf0U2boqJA3qNIFIssuRinWsY3X2Sf8jSmfc62dhPfk9sUzzewRYdPQf
wJc5utaK3pOXEwYVWZOzGWDEUqg1eevjw3+6pYmbbfRYd36vZlPVETnx4UJ7MB81ismHLIU/h2eT
QWrP0XZ+rewR0OHJnPaZVNozEEz5M9qDg18NnFMZKH9rhf3HeKvJ7w0cQ/u8TctAhS5WEZYGdIcX
DnopktMVHbulbid555zMCQxrjdJxbqfVx8PwpGzU8LL0LP2gO3LY7to0zG8v/KoTinp1PEDCzBn8
O0M60u9Xqek9RWedvpZKM0SO9vahcjRIre+9N9q/AWOcSb3ia94EKynrsXAI2apGVZC1dVoRKSn0
RfS+9dMRXi3S8EUKUC0wRNOJEWEUagKqWh8vUhphDNCEdcqIG20jKB9ulhVz9cwLvATwmmY9H55P
HJfL41GG+x/9crnRhMi04AeeqqlHJwzPV9HSe1E5tfGwXiwzm1E8mxuAV9Q5OfSqf6lu9wm2Gsc+
JKGMEhnKyNRt2AwBS69E0xAVDaowNeENZfv9DaEll4PuXuAb/JNRbq/Zw/MtBXTNY4BCFiQtiaVx
LWxfh2SalxntQv18g0q0nJa8mb/1tL+6y36uG2AUmne8yWbJLQcck7MiJgvw15qJmxcNUUAbTlS6
8XufSsmmmzmOTATfCD9f+PoTmqbQyLDLZ7F0UvnGxp53rjavXe0JFCOB6wahiENQ635omhF7+pbE
HOOvbw+iex5+MHU4JwUQDdNS1HCFDAXPnffqquB37mpkIND0gKH83f1CCKOTndKSu2bgNtX+A5FV
4azdGXfnkuZ/MVCw1tfx/3rgNJ78gXzBqVptx8+1fLwtvvSU5+2VHZVUlI5Y4QXexDvW/FjcuMEl
GZr5F2P6eJVJXwQVlhnFDxm0jIYhnYmInIfLANjecAmHJHGCvhYgs2U6c34ZnR8CzEtKjiECtixB
G+HlOQKk0vM6W5zEz/9NwAhUK8Xj4yjGSSg+Gc3DgiViQOzeWy5mgrSH9vCji/syzNzGksoffuU4
CglATTXDzPOn9mB4M6Hl8BbNMoFRYSv+BMDretKduqWI/4KBD3i/YhryOFbhgvpU9xRcEFUtHRQt
FIIjN1Uyl54jaa+FJlXVwZh30SQ002vV8WVDqps7O97v+q2cgGRHzfGMZN7coX3Z44j74teNZuuG
KoYIyeJcGqcI9l5qSVE8YCO/Om59+9fTSn+pK/mpxQs9wn1CGMnZX0aCSAAzFkHUD/BfkSl+IfFv
Q/SQknU9wmeRIrKzdhlYPOGgPsvMK9j1CpQsn51/aW0qwmhHfiubDiJpi/IxYpR+14yf22O4GcZ+
YhgQ+AG0NkXaLhvmqBrvRWmscBH4rDecdtGbzX92kupvlF+3hDCqG1gfClYi4wVlrccdH03JRj2P
uiKt5hqVrV6ubUgubSWthbPdh562HY//ED3V2b5NK0OtUHIC+8bzkyETkT0u812pl/F9Yd9ytazx
oyuonw+r4Virur37CfV5JTPDv5vQifpFlwUQzkfffC9OeCz6sjpvOGZfF0LAsOxSUy6F1wVwH8BZ
Kv5Q04W0BVXWGdzg4O+VFfuvx/Hkurw2MksbJ0OFUunQVGaXbwzVNn4Im05yeXN8kuxhWcqFnATy
adywCujIeeg5GYq5kTK5Lrzq8HRcdjUOhLLxi+Dll5uxqxztRw6KVK8DMTQLiJdrlUrwDk3nKBAV
KZaJ42DVn/yshvACapyqcI232oc23Bceeh2r5qf+L9q9RIa7ywGTVd5FhQj3Z2ccHdl3t98lMjT+
xbu6HJuMG0SIZ2OWKrZI4pHbyLD82exElPs0FCTKzpVSaeOD5T4E27abLzwHDbk1yZxaR5uWVF/r
JP8bDCUh8To8bZEND5nOYAP37rXkycay3YJx7GFw2OALCGbq7fuYWvJ6FVmkxvjcpeLL1722J+QU
RBlKDOUFGI+fqcm8Obj0Dxj3InNeTRYN54dqQDAXweJJjz93thtCHjcBnRe73LoflsYd2E66xo5m
nc5Yg6jUCqxlxB+qd+ShQW7EVGipIlisyG87/NnUnJxuA30qAoGcKY8BSyoA6gXHJrHc0cXLOCEh
m/qmFLEZ5Gg2WSNQnRdfCVINTOH9o+e0SfANVTVXWhgHN4JEJioRb9PA4sAtkVBwWRwxk1/H4F9R
YN8fBdXUFv9PNe3n4x2iKpy5Mu1YSGRbKELB2nGckxXm+5rSKtciRcFTVNgwQoUu3ptb85Nd6xkc
AWHLhpvzd/bpXkG/AvKGFlwGu0OmbzFRu7Prifbt4ABjlKZXwyJZH7swfrO8Wgx2TK8Lz891ihWW
9qGwNiT1l8CTN/xdSjQAjX+epAS0Lrv/zzzRM6ItIjHomRiv2DyGEB7XtEFT2jM9kUjGNWR1lcAH
MyT2mfSYpVQKyceZCmA19oLymswhlVo8EuzG1onR9FyPk3PdUQb+CcGQ9aqZ0NOfOVVvM5BA2Fvt
baXwKaIHz+KDeeKewHhjeDLMHOivlqXXegqm+t/+RGhjMYw5xsprGE/WOGMA/ENc8mHGlgvxGLVj
QS5DulOvHljRXNmKKCIlKCFE3ELEufeIRmZZs8xKEUrJsRtqbTxJE/LRaxKiLB+T10SxiAakqHyo
H0qw/AxaKNbXWDt88TqVyB03ayDl7mI9MohGLzk0TICDwPS/bd6A/FX+khBRe7s6uK/DfoKFftd9
vJGkh7ftTWd8RyLwXdTD5TNwUS4w55owrr7YzKvE3f1unKZA6URxj6JpQ7t0oghrNEY24VwutXZo
8JPf0529gQ/bClYeaB6sxaiob6CnPIbDKNIcvHlQlmFuzSkwmpzZYpUE8la/lbqFpSvqbn//DXV/
HcoQ1bdk/ApqY37+4NelUOvZpGnp95HNtCTOG5HSzn2XnpvFm6XVOyUf3rgDuAmToLL+9SQbEDL/
YH+wNlopjAHQT+yAIycBCd265FbkupdWfWaGHumErmioAs+G7RcKbWK/3or4ckhaEojhIhKNfAZd
Y3ZtbP/35GHRQ9XGhQ2PjOa4Q+h3Ns2c2xa5g/dYqqzy007vPnAw4zT0GEbWN4ycGyx3VAUvnzJk
FEzzZzZS1vMGkmiiwAJUzOKCNSoxatvBJHPCpHgRA8hQunjtTEvhQRnR4UEFNEERuI5sLJVaQFHE
4YNZXnPrcFO+nnNxxErQRvTA3uQcYEToTgo9lLQVsS+UNazXQXDlgR/F3sk5XFBES9k99wdUNzpQ
d5jqhgU9iuqTxWhVFa9PJDhFnbWTuLXm1YEbD56SkYvzoqDTs1+epqY8IqQGDTF3MPrUqCZpTfGK
yy3N709i/1AidcEfhpPWz8RpVZeMHLtoq3/7hl3hYUV0xDV5rI33fK/tBMZ3EIXEz5QWtvs3tCPO
likOHUM30BNafJzC12yuaudJkGp+AFjkOnX427ZzBAi9GfhR3uEWz6/Cj8A1QKMYoSdowpO92x3p
MqPKYBaPjbvXMFDdabPAIQaZyFEwoGSpraA4uMRKhqpJKNdPAop9P9KFG1OvXZS4zWPF7w53nXTY
JrjNY+JvucHR/q28OZeI9C2LcvzJq6Lcmxyrphyxh0QqHuwmDWB6Mfvbdz51CogONtrPQLBeK0Pc
QSovnjZmoV45Gm+qVstfS7cA1c1Xw3yllcIX3qkStdvliooLDhje3I8v/yk/RYb2UwGspwUWHv9O
WMkhYNiKx93AdV3zET8F/gTnJukL9ZoP9rg9tQbmtCzBbjgEnZW6xTCUN/B66kAQR/GOyu8GGew/
yVPz9WkDiX17XoYSlf09BgSgymKiXeW+a5sjZGh0RIxyt6ai7foCno84VCEZnSkrHcmjzMByVQIm
PhdXjSPXwHGSvw+FYOzqNElGlAqkoAveu3AS7566l4RMkHxnJXjFoKdxYx9W4cO/qtvwUtQws8QN
svfhsdAeawwpSUOe7KE3liHZeRtdhEDDzJ/ZZNAf7+WDvkBBqbC+ULME0K9RsK0RpooPUlqoPjuP
wvc7gOP12tqejN9v4xDxyugLw7trJokBHI/2UIGYkCuI3t8hfkPoQ42k6XP27MvETu/M35qoc8kW
JxEJBTSNiLHEU+ccShqVudvEjRn7PhxaNAybg4xZ0O6E91wct5aCVBhAdE6IsdhMJNn3yBKG4ZKM
5ZZP25x3M9j6fqdztz8EBl6ccouIXv+vqD3tfXF00xxAsmfntsIQ30nvgaj+NkhF6gTLi6+16mw/
dAsFdFJ1V/TPBIp97phneAy77UG+Y5ZHIcObIsNd9O6kgUyqYXYPXOJIejb93a1dt12ExucrIR9K
wGGjj6dZVoojxGOXnNVDN0ryf0PA9Skc55GsWDNFPDv8RTv6tjIoUQWxku/ct3ErlfFJUD4Swuhs
pIaHMs8uTF1dJUUeITlJN6RRsfo9ZSPlO0uVt0r20h4bGJ0kSs3Ut7pt0xHZLwj1w6knEBS8Umxa
QjYwmuzCUbdFAKa88En9qsftyzzPGfSzD3DRSSJnXp1rRKBykrlQt9wC+2m1JDSqkiaGTuyjHNin
ZI0GlVzR7VzZO6hNOZhM8b+g2jSdHyAlwdBTKDXyzgkywTe55q/aWFhWXhjU1Xu1diW/nOnoqLDl
95fy7eqNMo8vbE2BJLvswDiu6ppzBgXknrdyIMvPlc1NWjvz27m9A65fEVzxiYZuNeFQyrUnSv5u
+p0kyg+FD6uD6ogZkBRHnB+UmKZM0k6uWd4yzirdJvYcVPh+eMu7YtbiLknaHIzzN4r3hz9fygrV
+eRKABrXn/fqgnOHHLC8FI4zpD1sWf7RiwnM0P04EPG7St7DDUaZw0XNVew1JwHqgCGKTsIKxEJ/
fQqOrOslUBHjjwhQDhuEG4HatjI04749OH5f/wjkza8Q+dBnxRQ5V9zyu7PAcrlrDzY1wVxMdxwp
BWdaELqlEcIIkS3MS8KxCpyO4xuEBTyxGhwvfI1C9KnmwpLroiFN9J6GN2jDUu6ap1J/f4dNQ+sj
ijK54UVuzGPjo0uMpAw4VJWpxE3ydhO3ELbG32v102zJnelCnjuRz+n+PYTY7zAxJOq3hB33C32M
Z0Azoirhu/W0gH22c4bH+TxoRz9yBwUoAt+Etr18BRaEG7kC/3uT92/2CKOYU8KZuKgV/53gWlD8
LnUTN371A84zzlea/L6CdnF5IAmes6bzsv2vTpuvxTYDJW6cix/EXKR3vaEeoqACqPXnruWerF/w
Xibu3gXtPrxEnkR0sFglvw2G0PaL0ZAw5IlZAfSjGL8QBrTAZ3EMX1NzFJVXR+unJ2Q90Tuu84Wt
rKRSaZvAFnA04x2v+DzW5lkldgrhnGVIHbZSfjjZQUKtRog7Nw3OcTLMjIcDb2cykUZbzjkvQ4qL
gQjg8OaHI1hKQ661EYbS/j87FurIPuL+PL4BT7+LLDE23hTnNrjNy0c375WpYwIeppRxsX50UTP8
7v6iVefPNeHhgT6cJFAPGsxWtTYEaD4cXI7+0buWu84wz3rANynZX46REYS56jq3So0SthAkMSnm
OEoCDwmKx9L0XvBDzn976BYVAXoL5xy+TfjbJqkyOQudCRMdpJZuMB54ihxzCQtkVckEJJoTsyMo
vCDWMuuBNfEQWtYtXhB4sNJYfVyqbAivUtKswybSV0036oXlWcFHmA/FvXtVofrvWbjhJEZ14Zrd
XhkGJ+d30/RfqUizqSnWhbEuEOoyM/C691CB8CO1vsraF5pgWqIoocpJ61WEmYxUFANP7xHfu8ht
n7Gob3SKZfYHyfJ/RI6/Yghrc6w8wQOFwqAIV8AXjNzgNnEPpPpjtz+Izxqr3lGY5/qMg09Zt4f5
1SaK9phfZUuu+zzZlXggDY31v0fTO8C2mR//hvDBdHYeH+1PGE7rWCddXTT8leZv48dNI9om+XKx
HWSTUl402qGexLB7AjdQQadrbC055/5+QiPdcVrxbSiXShIfARUXs+hmfPs3FTmuGaA5OcV41mVV
2K35i4iHiIB0liifrVtbeuz7/dSWJSuTL0KFRSbH8ynN0XGyzz2Yhl8ijHs6RuipnSlLpmRklCUj
WJy+0nhEiDXFwpgfEdAyzSz5P/zyGoopETpLRi7E4aC4xPeoPSZmzOQcf8eOTqzUoURJYHly/05z
9hJd7ZbPE/wMYKiOLOOC7XwZpmQT6LY/hLAnSGrVSczns77KqvtidFu1PnA5ae3DyCqiKR1V+Jji
YCQcpFf8VuVV+u1W+L5L4ccGj5XYW7FFVHAneVqIvmXHjViKZcysxbl/ECJeIdONuf3uhWKZSAms
2UGNuywGde6KVdnVf+zVzQR62fiJNofvgHmn0gG2aFKEPYj00v2GbvdYDazFnL16UrjxD0tU9Qbp
tH9S9BqSWVTFh0UpMCQPD/qSSURcjH7R92AtFfblNLkoRbU1aBSuuTReKu57woC4+GZGUc34/dsT
KA8RhMdjLot7TNDYvgbpH+0utjronTSKSi8Li0X2Ybxi1aD9lZ0YWdyvrVi0wgJo1QlmSy3ukFZY
3uhbKzTi08OTSS+cmkJBiDSOqcfogLiSw+hcbbOXKB1m77qrLUpB5v2DiXPDVmOgXWVNyS5VirkA
xiN1ir5GFKOShyJM60Mbl2WapvOu1tOefwEdgAQFkv+0av1UPShQIrmUhucp6a3cSBJRT1JHPbBR
YnZw3XRxuuPFrdMHaSKjpUa4O2VLfi/4sjKkAWpZIsq3EgE0WTnRdFY5v3+2Zr1iCutEp3rKAeRi
d4RDnOHeYvu+3h+xPJpvPnoo5tmnHV10t72aQlSCPCvsr8IEEGL3djJGw5v0sQM2Xuf2wNj1Zh/1
PGmw7Nc4LrZE8PQkWNwmDccjrL0/2RIBY0ddwXeHSxJs9ckpJehdm2dY24pTvokhixIOykNUgIU2
OvQQkfTzKJBwsudkfJP/Id9FSGOXlHBbW97J+mBa3uXTS8WwLxJSvEnU29F/n9R8SdAZyThTejZF
ULfE4nWuMvtqwU97MiIktUxHPsu4voIR5d8ElGNTurPQfAMgJPuK1AhIPSVrFQomu1PlODLKLRN+
Q+bHfkmu90LO+sHoqR741WRWBFfZ0jgudJ+6tDtte2YcdoguVKKxmM4z6fwHNJzfurLUbSrl+vPn
nE2m6/brWyUdo3cDTNS3PjKde7VQg3Qgzs1JMOls9pUods3+YtrQnFIDnuZQAj8Vqv4lZqX/iGSp
DslK459eOWesehFIDETR6DZZ3xE7XDGVTrSlJDlu+p84BviG40aS/xVLfBUYmJa4q5wDbEc6VrQJ
3oLtDSdXwPMyeh2qFKTTbzlQl9EusjAJrgoHXh1jQK44X/eKo92zRCLNFU4LVUga+YyCvAYPjuXw
/SRFeakK+YXFAahFg+zJXmoUeVp9d80LlVi48J+TgRICy0MgGojJ+0SWRfxRSWYkMXNZd0dKKw6v
GkJ4l98kluROh0mqI9gI80rZ0qMlsag/w3TBZXEodUvwZgA/jMR6sQxYGo/vjyDg92P/LZL0n8J0
63G7baIbm70ZUPFUQMWWyMGdAw9CHUSBj0ARYWfF3hzvnv6d/q8gOclsRsHdfnbIJ1Q9pNhsA2Ki
XC/a/cpdS3YULTqB1duzAHBQsGt0xYs8g+rHBZ2IecIYkHHlmBJasKTWGyMloSMtOhjWeYh0EQ70
HBj4NZeB+r43TCkZYorzdwV6S2J7F/8uk0dikPQdtzrjbNFYqTlFGCIIQ6CSKPhqYz0FtnR1XgPm
oQPGIaJ4DbxkdnxOVnWZ00diiCEY359V7uH4BuaSSFpl0Czy87ITCvST038hi3BlESW3ig7Le0zC
yDIT1hdnap7vEdy7hh0tzwpPocxJc4GSXd1SQ34EGtqrD8XlU1eQb8jnR7OPDada1r4JpQ+WA6nx
3n22g/GubOBFNiQyhIKezlbDknNRs3DftDWwC+okDcUtMcK7x8jtEbYkSn64RFE4FqQ2GY95h10B
uVhFSGDAHEEuzoi6MlEvFTfU+iAqkGGnFmmoKyan3kozFnrF9WUYrA1EbRi5mA2G9JAn67pBwiEX
ArEm5cdtrELWc3V4VIgMel2yL4tCUXSSo8zRg6cpV149fo5ZZ1VLeVYGXoHxOrpVVWnFkzqX/QRo
2LMh2ylRJgLUKJKZjP9r/GYpKNTT3v8Ft4agRFODKipFdr7TIJRBDO3XmRaox4WIJptHoObLHsWI
zlhzcXUkNTDWNTeiENCoPD5yW08V9fJ8QZ/cxg6A2/aCcCYcCnHaQRa5NEa5fq35p9eZq9eO5Mn4
7Wbr2bL1CGROEQGTPqJSLW5NSHMM/bZU45dcG8BA9RPtQNBagIP/8h3Be7iwPCYhq9odibOJIN+i
mNvBI1apxqHD2H8nXsKpfTLm8N3gNTwU+wRRWkB2v3HaJg8kKC/xsuLCMzQiCWm+6hb4xzDDJ5lP
7yQBd0Run6TKlNN3OzDgwtUz/MfHLuwSh6fBZvBe53ZBA1HU+lGRu6W44WUS7LMt478eUSB2bBrx
8ZO771OeBrhg1flTgAcrc5Io1nGyxDR2/Y2yTNDi8XfKzr8YyJLY9mrxstOuBHsu3ng4/GonwZVW
1dbI9In80lkraVJvFfcrydVdtkJdg8GMaPbK5kn3ry6jwE3LiI1Ebrqq7eQbB/j3y0KXKqXhuzek
PfqgNcoF1+C9Y3oY6sqk6Wg0kAZvuShWIdBkBSKbi6bwydXgaGd6NzpvrZQOg4N63wLvI0YkRQsb
D/Z+JMSi6A2xXavbCHid4Vlvjwym8nBFi9IoH5UT38hGnJg7NjM/9EppPmY/1GC++LfDEI4lPV0Y
wrGWYZ7XVH9Vpbq2wTU9N6bx3bIVDU5lG/2BvuLRFTgc0uWfZw9go93H3TmFoSy0D7saNHbZha0I
r2bI988XMjwJORoXls2m3v9VCWO53F9t+JoGcruwffV70IdENKVNGOpcwwOwN1FNcG9rMevk+tAr
UDPL0pyFStSGj1nzkz1Y+QoQ9Mlc15tgO8DnKJ8XZjtmi4KRmAtJJqL0GgDIdeGagLcCQNuejKdU
TusQnN3sIeMAuDp7lzIkmXwz1Fdt3VfDgmPtV0rmfYAZEcU7KlyCUHK7BIl8Juh0Ve9hrWhoKSR/
Ufui3fkOJuXU7Tfz+KkYcyizWaLWtIAPZgvzSSI5c/Ett8GTKBLqoznQ9qGnJrHp95M6uo5ShaPL
VH2tBSGUnq1Px/m82pFxm7bn7+t1RDKZR+iLChJ1YlafvzOwO51gg8tTYvbLLbPqFPshP11bDWIj
WepqCm6DVcvZcSbYkOAQlw+GLnCNg8jriZkk41m6rH4GIIemrnAP4EbW6gkLZCtPtjem5PxJUwJD
HKuwXOD6PqJs3hvnTixHuqnFG2MHYgkeKhdQthXUSzykINdeUga8j9ZLoc5T1HACCPzQTtw41FJe
m2xTB6jTaFV6Aq+y8k9y9wFaN4dcyz1GEhuqSzFldgfONiefQ7tExjIsVw3a07tUplmDklT4WDgJ
9TQIJP4xTIH50Wrow0gLmZIT7YPf2KCgRYNUSkKL64G2DV+nj30dTlsOOHqdQzCdgT/d+SlFgpXw
qf7NbrFMMAtog4k1NHQ48gLGHutsbd6y8i0iXIbS/2wmlHWZnnvn+LFwFCJIopkPfZCoXFBuU4bs
DYfkdpOsiyUZLA/hooOvIWuRwM4UjtV1y/wOvi3b85cvSQfQDNlkMrKNAEO9l6ZKfh9PcB1yb1Oo
7pftv0th3iDFRt3I9pWHg6I/BZf+DmiMUHFHXrpXr9NWQNbsG5doSEPQnKr/tRPDONnENrElgdlh
LWx5L9So9UnVonJoYQD+jvtlQ8rTq5Tnx279ec/0+moEemYgeQdSSZSZSSnERgWKH+A4PtH6wyth
pxk2X7mXcZspqrzw1+Ym0W1jgiPLfPfZ7Lo+T6PPIZp0njZTusQ7ixYYeGL5c40vC2dCRSJztr4x
hlXKK2rPuyk0pYgxG9sGClHPcLlXEQRSTCsBYFeOw9M0sCze1uE3DE0LXK14DWmCjnmNkpSEClRD
lazowG04RPwhcls4j6TfJn4pVtMNKkzAJtRoZwDJnEbVqpN7JHujp7wmC26XKQBddsSbQEoXzNsq
nQKLEMvzxyFQjkzk+hloZ79ByY/ykmgeBIDsId5fqjO3590doIwegJZWwAKZ96airNRQYFhuNcun
YwpVb7uLVWZ2O1MQAOMnUj7k42bSZagJaElIQk6c5waGwDyotlaLGpf8uVZSsMZnn8KmsiUEq8jK
bbZYdtOs5JlqW7vOhKECKNLzaaBmeojXbN8F38wtfmSZmV7OwjxUGPikzhXaYgCNSpifho+FmYgq
Vi04jfNfXe6ZTmeCpNAkV52uG28jx1G0NpC0uBZwTARBs9qoW6tnGYJ9jz+aDZPdj8Cd3mDR3QOJ
J5QBhWoW0fY3aheWaDniXYrt6j4DXshRqIh6n2zXD8YNJbJvkqXlyUr5N6Mh8BZNM+XcpOCSykA3
YsZJi7pyuLHOb3SSK8krjC8IzotX2M9pjQeGyGryF+5KIC/5msn/FyMJTcg37u5sPKCTclNpSiwF
pi12Jy5Rxc/hBOjETMM4Pd2uvK12DA4ZnFTS6wchiXDWEnTxTBBYJqB/RC+iAies6GjxczwaxLlR
i6qHB6kiFdiq0ASbx50pZ6dAir+5yRdoIgBj9cVORPH5wOCg6DaBG549ug2xGa3WS48w96mrXecD
OSn55zZBin7W6skUq2TU2ZHSRTL64tj7gItB97jxTd7PS/IpgcVcV8KDQa1PmiS0iwRMtZBHKrfe
oMVQR/nvot6P9d+FT0jw1mUu+sIpYXdL50Sb5lVlUJuc4SjlLyLz4BVLiK5udLa+CMvL9zpWNefL
tFesNvtsP+kLP1781eMX57cp+C2XTTUTkaSez8AJaOyyjEOwc4FR9e4X1Xa+qOzk+yyDblCNOuez
aRMkWii5n3Hg+gi/qCeYEGqiCZPs8S+icsk0LHDA5C6p/LLQoN77+r+yxIaiLTfaDQvbEDbZPG2x
B89tJhkwKAODoCFAb3up1Q7jnDRNoqt8V7bzjkjSnJH9/vk5W8s4IDYmI+pMGx5gm2XE1KviIQVJ
nO+le/XYAyfnknLwU+SmLRHrbaf8ff3+d6wzEu9J9Zbc6xyEC0TgN2rE2O6Lc5Y2OXqAKOoiKWjy
A1MN4ZGUmnZuHill7E0PtmjnV74QkJjdpDywWhdV/3kmab3O7fR0zXI0BaJZ7DD4mkwkGynHbytO
6pk0BErXGmm2jXanma6YdN1IbHEjuOKB2iTYWFtLW9xayV0Ikm8ujpWswlya2l9BUwjFAXJ3B2Sy
QL4MaZrKToo2c3LD1I4N9HJW7180FNk+udz4UfrveXC86Cjyu4ejN7k6rLCAY8Tn39wQt6opYZB8
CROZuBAiuld/vcYWFIOPfAMmmUSzWF4t8Loa9ES1TwxXyMl22iLhHcMTXB5hjgctO0x/GJ+yXoOY
G63DRlHRB1dNpG8D9vZrm9gf4bmVZaXil+ql/j1o36raLQ0srdV+Ui7SGQb4gEE0y9LTIBsGY938
ojtiOWOc3vC+CJ5SH6om+szEYNpAYBOXDUbdIj6d/I4b3S358hC1rgeWQ/AlFZeLAZQrmQb02kZL
kAA6vatX+qp05FIsYUwlkBJGCUG09hUu+ZMLclcOeBWN+eavDC3NuA9jdcTd6U86lrZuztsHgkQX
wWeob6UgQVk6neHDFADHUE4KHLcasezK0k0Q9gOqhfJsXjrFb8wNq5jaBauUjVUxYtkAznl+Ay9z
C9QfqG8MBNtj56FwA4ljDJDnpUyv4WDQALhkLmHpkM9dK3g8Cu9b1/n5+d6b1RhVbSQkv385mpOu
bGdSHF6cWdV4MC1ZJh5KMnP+LcrQwTMFaz4SY0OW1smd3LFyN/i6N/n94iC4DzZkbUp04JXkPQVF
zNOOG6phIn0tO/0zssTDoRWxhB4sCOlgHGgD0jmEmtlq1HQL/x7mcZhWZyPcNjy7FXT2Am/R3bLQ
qgRvnY/Zshj7tJdKW5Wk7f3FU5xauX1/hz1sGAHwXk8So+ukSgQJWGIsqQBgoUSbH+/PhrIRlVUk
T2V4n0446ccXJPMyYjzJty8jLiyAJl6Opy5u4fQXysULFQCp/36tLVqN9BVcpaz808zbUzdOEDm5
FW+oh514isk4o9BerzFIKPVxTiYkgBjo4RcNdr9eU9ejxVWsOpvXG5jnlljpMZbD95GiNwyxtq7n
Kj9ZTXsJtitbf5x8UXnnbNODQsxbhOrULFOp6TTrXTbfgG5WF7Nkw4zeVWv5KSejVyJSLCqWQ4QF
NcOGDT+HXZC6n6mx9HE3FLugWM/oXABuFg88IVbt36Gmw/q7tCQE9g6H+lZshrL22bwgfeUkB4Bh
NVdCbR0JZdd6zS+90deiYkpuN+nielK2gho8VNheIw2U9BnKHBFqbwGrwdnFLQv+7AeT/YGzjoT7
pg8baF+BsnZdR8PGN6mfdSKQzLHGST6M4OHF0puNdx59IryHQhNmoqmcGcxRHAgNhP6BF0A/dzyJ
OoWtS4Utvd1gZpG7M5o0CV8VpewnXdptB9I26dDIif3PrcLDD0f9y/oTQKN+AvXFv+y66Xe7MXld
lzueuKxGWFluPz+ZrKjTR5KE3OQ6sxqmBGJHzmnT7qSQ3i76baQ6k3HHF8cn1Sa5OFpZf92yVwOR
Jn6LyEo/8CtpEaeSNlmvyTydZZMIBsnsDZe916kLWg/2NZ7uxr7hRl2WBmnuFRlyh9UY5egh9/pG
CgFL+pwYS4+W5C2/GcliI2r1KOKlZl9TuAypEkRtXy1hrciOEfDA0Y+uBTYXqnJBCsTHkgT4zvV5
4qtx0aeMTIVQXFDi6Wyq12BW5khuDXE+zQIu+S/owqAqbI6UkCcJwniWabWmDJIxToJ5Sfflfj/a
aLZFgOh5XEDguX6MBpeXFGxp5A7/pMj55Fcj+L6M8MRrNzaXcXU31voXgzzkpRhoXrZTZhcgSeGC
3j4rWrRNgpIa6UnvYj8QglEzE+J+g0/5XTRfB74BF4To2XO/i9t6YgRYC2Hdp2W1QfoJ0TAQBWMg
RCNbK1OPooQrVYAtGpfsRa6z1TVjkx+c7csGsDPpUM54uWXGU+5HXIyyF/qnq/RCkAtPeG6Frk3G
fe6tTKalDoa/jc+kNS/yi9quynlhhui0CH13GsJORVv/L2Br0X7hXjM0KBBc5OgA2OWA+qb0breF
gLa2bofH0fC0ERXr7hD3XKivAg6X+zowaZE5uXZQGHdkKvQum7sJn2aubaKTkpQo65RSIWsM+hH0
H6bbjo0KKQbQfu6nkk0frVjzObmSVVRXevXDqH+vrB5abbCFFCSM8jlnevS58UNx+ks6YxfXugdZ
weBqyfuuQtnKyZ+QCnzIzjhob7u0F2Q1IkIKRolt9gRLGivrk2HcggrcyLzqP0PjVcx+4kTJ21x6
5IflfBOLLzJKp/v7KVojHIFHiJPInQC617Zvs5JQYxdiTqjYN6Jsbhip3u2OOgC3cHxD3VIOBp1v
zF0obw3bpZaCllk02MmjIEOOOZj27K9nUj7FONUoEgI3+h2LrD0rHHTynfRaOXPhjKnOu0BOJu1b
zqNbjB5H9ySIK6YP5B29WTO2vL8Fu5OpIG09c+7yP/N1jvbBOEkAhwyTqa7KhA6ZLYN5+9cX9akb
RENEd/hyQ5M1Afs5i/ap0KOLgbQiS1Z1G1vzt43qKTJJjO4kvC0BaDUKzzvAdVVy63VqfHJF4vP/
uBrgIguY3mf1xYTcQsIK1Ad1ca8gXwuJCvAg9co0Kky/DXwDH3jEcyoae4HmFwUfgkTR/aMNVQlO
PNhxenSqjPQCpCOAEPfaGwf01OXzmvE8Q1pqz5kqMJvwUk32ITrP/LN9YZtxXyVoZjXh980EZHsG
Dzr2cAt6PsALIDIc5IuJm6BuZS9oNAECCLnFsEjTNHNXd4f6G6dXTN0pArsbloGEae+9FzfhCOg4
+yuVxdd82bBToyVWa/qFEmgH7SHr0o4KTKnFKcCyof2PtZ9e7wTyh15QG/dv0QXpk1O+hbhofpvM
v38ti26ZEXrqoylbabImmSVbORE5ipJSwNFAz+yvYO6LXkVNnLymjJBolwPBQA2w4OgVDzgeJeSD
mO8iFnF31R/8Q+sr98SeFIIak9zlyCncsWFchwTJMLSXx+Ucynz8/wGNEywI5d8Ze6Gsi/mxIvhH
weo/PLndv6O5serpyvjJyadaFpjDaE+nalNMEAqyNwY/XPGwb3qm3fdeeXYYxuM2740JP08N4XL/
qExaS08IE+5g/DD0F3xbvLNGNWCpjRhaALB0Ebj5WpoFC1w5cL5oGGjv/xqewwX8tctfNSBhXKnD
TUDagMEwXLTtMPeakbjxWS0q8YrKRxzrFAfE0XDudyiPfDf8eCi0hUbGckragRF6JigdXJXlBw6P
2oXa4oIorn/4xW7bVPiCarZwAkxEWfifm+92ISjmh0ulfAYtJ06I3bO0veguQsekjy6mtvHq3s1M
g1+1zYZ0Vf9B98zaSVihhzDLm20dqJwb/dpWi5tZvgKTm7mgvGSVX9h2va4jIP0pf0o/u0iG2dLE
WdvCn4pHXmYxbuSFWEM3rR+leZkvrFjO+NIlpl2fMuNxiBL9wn3ZiV4HQ6u/Q72eKuXlhC+CHo7I
IYDZo0JiJFuCi/SPJBxdgBJUHRA2uSQ8fusCDJgWQhYVlzwGi4CYjEXXCPs9d20qnxh9OjLU+i8k
kW07+H+sIpFIysO9+6mLnQDjINfXc0hmqU5K5UbCiKt58XYqrDk2UC+MDKk14cwZxuEwaZhOLTCn
MBiDa88O1xlopwfLyiX3zBTQvxvYlYsn7SLm05rlSc7wlNdgcy4xS2DNWU2JajBBkIjPc8M83nXl
BLEtb5m4L/mgsRxEOg8DOPf3dsssgXpEht/ltKSeQg6P6kFD/mhTbO25GLt3T6EKxTOXPzIQHdeP
Ct9FE9PdhsiSqymgeuUyx2cBQjsWsvlY2ukTUVTKAX4KK+kN7GzFuToLyQ8JALcUB5LFiBUS+qzO
2q2yhV10Jyvwyc8WQdCUEwdiIgplVxI5sCeomsDTG9DmQEYUfvNwABR+CpS7QdYLYDX0xOrMW1++
7VG9ydDLW0NDKJwIyDGz3MO6Xt5YP+GCoIREjEixcjJdDdmoUVxUjmaoBV3fYUnB0FLS8TjdJV5c
ClJs6ydL1lQr6+z5eMZive3HaZk5u0y0u+hLr8zseHxEKDqBdAojPCND/sJZidiG7kkf738h/+Ym
zg2p0BuwsStrEz1BB2fVjtrIIE+3MVPL4PUyDBKyO3hNSkUiZGUHMsdDXwxYfVsbWuKyjPrhjJe3
Ps0Xqfs22mC72/by2il3Y8NWF8ypgoVVpHH+P3uDiWDSONrZI56KA4Pti4iuyZg1oN/V7yYz1IIH
T8FEO4FCiW4CcPIQ0FsVDti0yKAowcbDUD3pOAZ11dSmYe6ds4eLM7SJyXERgj0mTq3ZMoU4mapd
927GygrQldglvm7Yy2IyZj4+cdfgYE5o+eEh5QF0ffuwprRDVwVilp03DOhV6f+nUGu0QA0Ivsr4
tLaYrMUi+QypxB1XcT1VHZDi+Hhr1/WcwiTpXCavJXeDP1h0W4UnSMLrTcEJe7u9mNJ9OmumqW+S
5HsWfhNBDuZclvpKcRgbRBEbUbYVZIPVr7piu5foTyVQaoeGuKV6jm5y0gsT6dWxy+uroEd7bo5h
7wXCyGl7sU+IjbEKKIpZzyxJUwzZYIgegg+TimhT5qeGNFpBERvg5JRiH+h+Pkxt6zGbSXzEvPsf
Us+WLoYebCBZfaSVjCO7Cs3r7qbY2vJIFJHqGHn7Ci9wiSeGcLp4yZCFeK0YIKGngkRj6aPqfyxw
U/jZWtIRTSfCtg4+yaoq7QJgJHC1PF2hPdZ18kksO1iGpiJAp8qWHr3gYUVFPIWq8Vji8tQeA5nx
r5c1TwtMId0AmkFfSRCZzZKRmwpDib9y0xlgIxGScDvCZ/4UkCOe5uWdoumSm/jEKMG9LvkQcRme
OJFTeGJh6ldKMmjuTCTB3IXi0iUiuh5MvOR09mfTuZs3eN5Ag9oQOrDui3jTNvCJGDm8Eu2o5PwD
9zEdByGXN99sbj/oBvJV27R/w2vqBZpCB3aGRpsUrFtwC4oUYx325Sua9OAxLyzQNfGLTRqyG6XI
gC7W5vadOXZyOwtXQ25kVbrBFrrs6R/wt9IUTj+TcekP8niMnjdfKZ+NP38gzyAQNLh1EC6X5WqI
qsyCNStFGovXd435Ub33B0FZ+FmB7tENZi4OC8mzZzkT3t9bueoxwvKGjetIuPwzSUbV/+bZwVWz
EEEXepMYiVI4y+se7a3Ento1wnv1pMRAgoAhbIvf9YXg7Ru3Wtn3NUQPhd3sRy7MGJ/FL8tqyIED
LGV4XDcwueO6SAu5leNICxSlFv8VK6eTil58aqlURE1+Pmjx8WZh0uRaGd7OqrKlzV0nzDp07uEI
Ub7vkW4lShozmGkYUkYXJoFR7EIgo7oaSyNCY7mqGFeFpeOvxjqynsa7laUCxcPZMX2kdbX131zr
ukP5wfiliDadKMqXeI7+QJzkBxw9fQ5l4y+Cj/Ue4keR4LgGDJ3SPG1PU8wp8G8wVcuN+zJcnYZ9
iwI84ck7+Qvi5l11eWIkfbDrCHS1MVNdfeAXr9JKOmR44HvcmZtm2XzMzEGh2dj1++PbHPzy6AQX
OuRwPmGGqpnGwSzBPon4UR0YTx6N9GaSuKmSocvFO/9sviMK0gP+VVzJyq5xDfIdJdNQ2ex2yA9J
HQBnbDLJFTbiWe90NP3DarsFdaLPlYrPOJU51FlfC10sqdNWNKcesbcizcUbpa9xCwXOGdyH/JXX
M1OwtEtL8o88OAhpMcFsJ7EwVvMdh67gRYrQegYXzgFoQRGzvgYYPgSFS8BAN3MEJDoiLOqx4iWM
yS4GilKa1j4EvxvmPNrb36T36YzWR71OMA/iuCKAGz8OezvAEIbF9po3N6n2DQrLMmyFpbZeuSQD
Vx2olvroJJvlSaBl1sTIlBkfPEhtK6QLaBQMP/sh9xwNqIRxQYrxdYVSIDFMUg2BjvndX11JL5RA
64mgFvU5a4yL4qv66avNRbKii0DGvLr4pQ2qRwRNGo4L2Zhix0AyK6pnJdb0ms3KQj14voQpAcHN
HJ6W8bjimVpyjps0+DqGEZkvYW6hk2SA5L5o96dS0lEhVF9d8PTCSmSz5rw64TiwQs+7ae/4Updb
tQ2NXBPJeB0EhmGSeIFSoD0iqp5NXiHoshPW6QJ0tfW1DMcLboEi9nmmdaqxjLt3lGCYKuw5fPpE
palNnGusMzErePyJOcY738u1k1+pmxayVogpiOgYS3wvMKOTxuwD4QmAyTSJO3Mn1d66P/SbzdTr
a3yZh1gtXabsb1RXMCp9aMEqBmW/uM5meV/CVIM5Z8FSFkDwchoVAaSrevGxrpRHoeb1lQT4Oe1z
FR8AcEGlGsQQEWzarno1DdtYdyUo0BLLNIpoptZVK2m3wWPvYY1TVoAteaKZuJvYuP2hUnzZeBtL
iHFO/C92mZg82OX5Pudi6VcOpV4yu81RbbqUWHOU82YdXIF9CNJW5LQctxaiIdfX/hajvSoBFgMv
h1NUYdzrBv//ZcIyIRfiQYSqnYFMB7qrQuDgSd/stKBKd+21RlE2CcXpyZKJcnwCe4b81VPmCqNs
frkzd3YuRUJwnmW6ya07oONI0PBJBNe/6CKUXXdUlBVONe37zYCETY+sitXjxv9/UTw2YKQ/DOKv
4QLw0ZJGFj7q6TOYDerZ4FpXSM9qbs4rebQj/2xuh57T0vkjBqTbjlx65trHmR3oxvcJbkTtmdDo
Wcmp8Zpt1L9fwD0eNHHNpgij/9aMaq8U/viDpQ+B0dkeoaKje93FmyHf7lcLb97XF/jJ3g9xVw4h
9P3f9tNiA7yZn7+563L15+UwZrNAO1GA+Wajsq211Aen+YrGLX7HFF3C0urGPHooDEKzS9wqfgFI
VWWYmQeDGxBuyl6MU1Q5mImzK3RFbsWjR9VbkDu/vHFCopZASO2iuTjz4ckWxT/JaVPAWWWVEV+k
s3GRMJNe4klSCWdxO255lCXNHAE36zwzQC04YQIDXbUJjQ+gOgeBuXxPGMduVFJcn+WRlvFzvfXA
5dz2hgpuKxWpnbqEpQgooNjuCTSeBe2PtKmZiprpZzAXaTzF4RpyA5Na/hk15NSmAUZ8JO+zA1B8
NPffdhbaCIzBWiSAGmQa1RVhbepbF533+F/OnChX9W7C0YsRIl2Y0mKJZEtmsRXFAUSkUbP8WqON
9MipebmsqPC4sJlNI/ArtilpWQZ+LpFqhMub0LjCFM0WcrwfPDCPGHV0AlaZzSutl5VYmqk4ymPh
Jg4MA/WBYvMzC6/BMWzHx5xNv8KJwgygcXTO1U97J3QHe4d64Oqb9f9w+Ob98KEzOQsLvwS5Jbov
0sRfJWDswkhzknB+ZFko0WCm2hX68OG4pvYgYEXuNeVaxgCl3PZAz7yn7E7H7bPrjytY3HbweMk3
igkG7TmBsmrXP2GUycPQw7wMbQmZgURPmd2jY93PPYYet+giIoNa1EOLLuK0nt5npJ93Vh8mNFQI
0OTqIT5MKIrQK/8d75vildEyypBStGGNnXQhXupSdzkna3tiI1t6bSQzoEa7pFVlgmPhUkmmgaZo
3kVW1owT/rkzVKAtfbg1JTWzhMcjnoFiJcmaHj1wsT7ccZL4ICncvgP8iTXhtHtD47Q0mDAiMdmR
cNiUCvhO5XCxsY3BoQ5XfETCuKwGhAx73ZiE2k8V6I3I/gN62J2qb5hJSgBfZklq7MU5wqP1/CCS
W/Fnn7TxtiPSazMWOo81gjp+6lBkUmnPhzod4o1LPU9CXOX46u7ki8OzeMBaDetfQrJR/oYe+xI/
0rdvX6HYlmQQgXZfzf888e8lu8LsktcwMZKlffQp7GESS/LbwFOGNc9Ro+YbAOX2pWjSeH/2iYgd
su/OaFw7JxSaHuFgn3tGLt/C8Bm1XyQOCu+MPzk6jggETw2TmFcuoQ1xrI2QggCA62OpfoCBkrGD
vsKAeSKis1OWJysfYIIokch4ZpDlvQJFX90DvhuoVhIZPWpJC+TpzeJEN97NQG2p93rrbfgLRq+a
sTXUd45mUnbl8wO0dcSH7uevqY5POO+wi1Z6TGY9LGWZkuYF/yNOgfXBQieIMLi3f2NYxPx2hObV
F6OXjiFZ11tkL5kKxGjGiQnJ7WLxurunnXVRovWWCFhAdbJSj+FbmG1we/itgqFQigON3My4+qMd
cCmrcgxC+krsvBY2S2WNHfFHgcNcs0Qj1xRqzKZB9RO5W2+S0T7583uVTcJ3Rt5riwodqw3YqQsq
zgMAPTgY1rlVn/LPD4U33ICz1g7N7pEefHnkz+2S8191z04Z07Ej5b3RG8/kIPrdBpdbSfmiZg2w
E8YSGrkFcCvL/ABv+kSKrGfd6sV6MyNxkDGuUWisXQRsb9Fo4929SYqz7aZPc/XWoKKxz3hVblUS
mtjTCNI1QRUBA7tYhf6O7gbh/uoiWaxteSJFIKz6MlwumNZ5UTkblJzR/b/8c4ZKy8VVqc5RUDZK
7ot6ktNIFc+oqPgqasu6LEddWD63+4UpoaiOpnSIFZxxbiRTMY/dCXiweZwfil5TnQjMc3DcM8ED
xvxCQmoQRD+555+miZuGUmrR+6Y5YDpmFUAAh/fvp9h7nLNvSpZ4aYWxztrlCPqvHk7nKd54/bsW
c6B3WMsiv9xrKkN+5U76z1i29hcVpjhh9H5NDM8QOdVlHl7EokmDtdvm9GHMIT7Lv32mV1fheOJz
Wdp5OxImD/tfLTCoVEHy/BYoqZcN1RxwZp5cg0x6/zcPsjJGpEQNf1MUsgJg0vnY4zH5JMpoBoCk
Aza9SWi95RQpcja5mm24A9rv0XOMvVNQupGPsW3SMl4RMt3/R+kJqS1NpfJg8S4oPh+0YIEmuWIZ
+YQcgs7nCVNuDhbdcDJK+ogwCPOcfTgxkrSh9XhnMRLZwZx3bJ56qPToHjIwx6TrNl6wEQ28zVR6
p/62dDjHTHDGHLH2joUnUotaS+awbHkt+JaU6Z6Jh0OKb6wC0v/rjCPsr/AUibMud2Vgy6WvtZBk
/sqkRN5SW3gBUdgNhetXkoRDYqy9t65LxNxvaPYvu9bwRCK3eya7BZY3T4h2VBo+H9UZ7sX0kfoE
4lxQy9k4ZO7YRvAEOjzN4OwOUXJyNILaIbXWz4YSdSmu0yCvKGjcAN+iFfJx2GI0NpG7yZB3qwlQ
W5wK+/oUCBWK/17fPdkmRk2DxhpPP7xJCQ9oCxMriQEUgnUzFXKEHgsBk0mF/WTZ7UqWgMjVk41I
1NvwXANoTWA1yulYi7nyytA6qz6S8/U1rokY/5eeiKEpNGDK86I0fV6vXwigUOiV7Z2wKCO1ItsZ
VZjhi+ucGRLtlC1nhEU/UtvOzwH+E8g+9EqgvExxXG9Bz1FqDs+28AZj4lzkm6McYcAsGpI1JXqI
zAvXoG/kIuYa5eMULUd4Blnk38E+lxhuD6fX7kTpxJTf92u+HXebMbW5X0Eu6qH+Ej8wIWyKEMQR
GxasBSTuNLVizLYy4KlUeY13/dkyLGRzrsSwAhy2mQs2CuiSNoyZkscooW2mRX2W5phlVYboa7WH
9wgBzhxWQ8Zzh9pqPOp4r2P9WAhqWNZ8ME2Nz9w0VQlZ+G4UxotSaKr7CCNBZsscHsHrMFE+jV2Y
oQR0iwX1UW0HvHjoWsKffUUxo0mIQh3acsoVfWU2xcxmxm6cAixoLm6jmYWMmp3QB4pRZbpzsv8w
10TTZWGSF6kyW3dSzL+NFtLOo3p+7EqBkdboU9no/veJ9+xJ38x0IM/v4dRmLMTggo5PuiTiT9GT
p/X++bGk2KOOJ1FKH8YwFvsFDStufjQp91KxAQOACSsJh+HtPJC9RpsSljAhCepKUiJcZuJBBaQf
n/6ISAJS/lR+bHAypPAeg09dmEW4+ESn5bJVi3/vJLRtvTtxXYiIlL8L4ftWZOb+AKkexnRkSEdO
dsB0/AUBiLrLikBLSBb122lgSsjgmuY+Nj1sx5KokOS1S0GJ65fdhwGxFMq8IvVwsuGySHTWlwJe
6yLbaxk9JEFTU02uM9badlk/yIB3Ow8b75mAy7gQRtVkT08WyTQMvrhpaGEEF9cjLPXSEy4rCJrz
3TsmFmIWinLKVu7p0bLR5t6QxPlL2nuasu5dg9vLtTP710fehuHx2L7AvAdu55Mq0XWi/JVKia1X
A/PC8TOKulonqxPGLKURtPEOUIYCOGXFCNxBRnij6Rf9p8GxUNcOF6iyE1IbaiexQFlOX8ygfUCG
yUavYF24TTBN4ylXxnTLRciy8TQYYycZa8BBqHHiCEgEkZmPnUE2s/4Sp5IuvjsOfkOv33Z3wiur
TDQC/+au0aolf9t5vzkKB50wsEX4O+QsmIlCrBCMZs0jKQ6m7f6H9LI86/vZKTKW80ZYvptXJfm/
bmQGcwuvzTGcwjbPGWb9xk+czeBaDKVOqKn5jN37FKwCMtceqNjDNnIVb+Xe6iJqUup98JhC1O/c
Kof2sBGzRFkTO19GfqprdodyiwRuQ5EEh/pD3yrnWBFJQqnFV1yVbL/b59PcT1TL9WrrogK8/6hL
IfmHJubCjonAyvGatIe3sC+oaSGv0d9V7ZggbLrCdmZFGBS+urvOEtA1PILom8GwolkeTTgkRtlZ
PTznSuhn5lFVH/TF97vJNmfT7lHY08iEpCunJyiLKX6JpZdhhy2Yr5vxI8InTFkAoooJHrPGrwld
T4t1nxQEDMnS8leLPBw5y8AKyqIbTB3KRbYf284hvHDnDNj4z+4NOIjMIXx6G5LuboIx+uLcGZVg
PYAn3tZtcdDGUKFhgKVuqZYQ5deLD4mSu460e9/5sy7bfPFd2jR9dJoWTyBSpNsvX2C0JMg7PuMs
nD3nyRYbjdPRYiSOnvc0eQhmUGlLSiLolOQESNdH1buHwqgFYZ3vehZWhy4L1WURKre2Og5Ub2Jk
pc6J4BJUpA3LaAPENwodpqac8F/yn0cAgudjLoimnM8RWcMXiS8xRobxlvNfV2f0IuQBQ4MOz0bv
E56iJj8KW4+AtJUB4LS58XFVul/fzMyihKK+DbVTH5nn21SUe72H4CEiSBvVKMLxfAcDPQSe3cTW
HnFgBPa+OegmICz0PJhDO59kFHrO1qulGmP+SJXrEupvubhz7uERDYHlAzV4q2a+yKaifbU6LCQD
fKaSC9USB/ejwp1S2+bP/TvH5hVGqURoNCPEhX6JsAxDNDXNjpUzhrkVB8dWXKGRA5rM7vnoltei
J/YnuXZBE0LmbWc1z9C79Mz6mwOz1hG4fJ3C9XUVf/J8zKHhhbtHOO8EbkxuEFMS8Ncv8pNm/cs6
AyvLdhKL5e+wmW0le1V6PCXFCXCiBUNSniWJOS34Vc14763+r0yUjN6Xca5vxVTHbXK1L0/yggB+
/IAKEaYqE2E+kceyfLS8aeA/I4EUzytSQz8eXwFFwmmuTJzlkdlMH6Hyq2pWcgOnL4G2utcdh6Wh
om4Fd5sIAc8/V1FvwkGBLcxze8PvAIenrpbM+wYhHhD46LnvxWI4MHFYCJxLPVrA4ZjTBeJy1+Xw
NmbmPalUU5ph1oB3BEkC20zMsPLdyLqwyrl9cwiwdIZYQtuBJVLcI02ZMUUUeB/TnhCV3i9x2XAb
YBGlvYmYWCyHzPEDu9hgzbxjV7nv/u32w02jGEXwx11lnMSCxyDcwG/HWeH/H7umdvxOj7/MmU4k
9WVOZAZM5lgyVcE3qwzYxFQySl1m2/M1Ds4IA+UtE9KDlqOCUOvMcDriakxIpv8ygVMvb3/loU1O
QjB0ZiavKl0oe1VdjaioAqeFOoBEDEOYy4mf1mnYcEUZxqcwX+7Ek+kahFEghTg8aHJiP5IdvKMB
4Z0VFeHctC1XvM5GDQjBMJyMJRGnZ732JjgKvphrryNZIe45bmKuVPwwEYy0KUn4j6ybGDjutyMY
RRxd5xntAmaKT9VSdFSSpoDIIVgj9zBax7G1OQju37bUMluPKdYfPo4+A5no3CzxlTMWIx5VoYCK
4OzoRnXZ/p+NZjoMT269u/flIY7qpw+1gMitFm6lF4pRCfUKH4ND86rLs3LYfD9mI+HtvnLdiK1N
52to/zvTewbZ1BoVyhotyl/GiwmTGkWHMz9SlEKerNv2khj/4ZEXG11vuMcsdIkg2I9fhAKo49lA
7gYQTZWwnDUe9gwGU7lrkZDX6cHTqgstA5Y/qcRQF4YQXzjaAlVKhl07EySDTSlCiREsIxbZJtqN
K3I1tx9ZGjEHcD2PJhTf8awoGfUjVARoXG7/HXuVrqUASSRZgGPHhdTDehLp/nti+QYS4zNFvQeZ
w+hs8LKOIy8KXlcg44r3Hq+VKE62vfBUsjKNTey4yOvgQKfzzDW3Ko4S1J+CrllDt2f0//WV6hd6
w5MUib2g/ZMEScCLkFUBZmy9ib9ECivFJnNObSv3CFNjfdRM5woySiqU251pkx/mJx+IEyLEqboW
9g2BHR63Afa4e+lzD/ZtXmVs1LkaSBriMk54MGbtkX1havtMgyRA8uCC+/l9pQiaHhXwsX9IyE9W
wOOZDKY0cWSfYxircSLGZgz3sdSwjHOSVWD6Q2UDMp5QdKqGuE8QnVL3Oj0C2juOATy0b50kEsDR
GW3fzfs77lpTsFPqtM3Izn280fcly8Is220JgD58ETVjmeqGJgy3HJKuzUecihhSVJX1CwLRdIgH
/GXc76eLnhJR0e1mWkOLdao7j3J7Qu2e3AZF6wcCP61GDAiAJz3KrNlUQmz0LpyORBSD0/wL7v2B
v6Klp9IMd8aUCzPqoYc1tvojWmy+8nuwMTz19tb1Nw52cDeqshInRJYPSg/aywzhxr0t0uVkuz90
ESbiKxJux4B0Ta9BoXt9yNtQBTMzz3p7s3LptN44fCdnvBwtRuy1QaD1LtndaESbdmlcW5GS9RRu
zsbAo/Z6RS5VDLZXMxPjYYh6VkrXJE4BHbDVSchdhpaOKsWbVWF9bs9pLjkJgKzgAFyal3Mk9bKy
OEJ1bJp4vodr6MYIIxvFAhnFEy+CAmhgUYLs/eocByfvRldzb3yLrriwpG9T9ORW0KNWTnG+DnlI
KAflN7wjl+uiTuaO/zhxI7inhLaoYhixOG7Rvd20aTtrTKEDSYeQw6moVEn5K5A8PSMG0ZxH2N18
ushisD42D+tTJHyct4uGz6s6nmWLUYiUFT3MHSS0k1YL7LIU/Y61korfTiLVAZL1tKQlFla6DWwZ
Hgy4sysDsmo3dA3Q54LXKkFOghS9MZv8fzIuBeMJfNglCdP9ZVvqWoUputvAVfHKgOc/t588/iti
0qEg9y/fG2K/n9Ht+k5uINxHj841os9QSdIJIiD3vQSmjXGQkSd8D384xNQFRsrLsLtFC22Uuqlx
qhAhI8PrlOahYfu+tUGB5nFOs+M9hyemPQ013E9RSq9XMzkBAqxDcANYipmSa6iMj16N8/ZjEPck
WahiVG6Vr71+hj45S14HRBrB1PpYkuCzOCU+iRwIL8+94ZOumP8EhGXnv/RZp3oA5/dU8XkBtEMA
LSfmlVPBX3RAqThvycYUex3ERoA7/9nXuUOVHmj58/o4gNbWOA4rEHoFY3GaTeUV3Az/HlLAPx3N
/C1N8jqRHsEFSaZekFQfX6GTNs4eXwGJdLvYRADPSGDU2fPLsR7yDgudre23+fqDcxBODivV/st6
ElGDA/k+1YPQzq5okqGvdO3dUC6Sjpce1AK6eVrWBVQ8ob+K1Wadm+1ybiBSYUGYs9ce5kM9EAqK
6YXO+BcP+OO7UY1Ml4wfUI1en9M0o44uMkTv4sbh+EdlOPHTkKt1gN9Ti9vNW9V8ssenva1Rdv/x
9pfRItBTnyD7s1AWarvLeT5TdL+2DT7fi6iqT1EE2qRoceszzkhSNYn4kkgmDrY7FSD4ET2MvzSX
2E8N/jGlU6ueE2g2Mhu1KmaF/2+0QjjQb4pXASLWnZ09OUKrx55JjfwDBvIHi990A6CAmhjbZD/c
jvm+xp5fmXWZLITC6MdWlwbA/eK+dHr0hQN3HEJDhchSmvgx1BSpMHgClcF0vZp01DrqOLRLHotc
e40vBHR01vaYWC4/+cwrjL6Wn9FjMjWjAPw+8cBouYcDnQxDmtWXQ6mYpDaBsoT2nXNUQ3UuGSMQ
bd5z3/qGEkVGviuxPyCMk6bR04KP/b8yuxUTjkT18PqTH+rZ/cHZF8A5rKw9ae0UFB9nJ6qzPM4h
8bLFRmfYhrzyM99tysvtsE2NkX3uOzZs3051VMjhgnsDwdIrW/GiJSYyRlpC2uZKzZy+ioznjLtu
va0d2bSt/S7dS2vLSAnuxt+tKZq9x34KbtlijPdtZNkX0YRNHQ8HRddZw6grO91AjKVSiAn0iBei
IfcmQGvOfhDplT2JcamtTdP0dqlaESk2Fz1IwZenWoAYTdO64LGswq1mx8O6wpNqLqD23+ZG71xY
MAKj5RmpjQptDz7FPL4Hyw1bM7Sbqmo7MgLlAzDWdZPfS7YHgkdB2Vz4CSsN+NJAhKbq2hGivtA8
e5qJrDoXlH771hWlD46AR3Nvb25FM4FmUBrDNK4wfxG9BqnEduuGaAttNjyS2FotyP4olfpo71zu
SI3H/KNrdblNhqpuPcV+98uNnanlE+gnxxTPpYprcRaieXUChAnN1xZ6n0Mke8Eij8BLfWkrvsmh
zRV5Ogn6+GDQjKXvdpyzmIXjMT/E6wirzGkEr7AI+aTs4s0n8G0doyfaZn8SIsbZYSIEgPDuZko4
ydRww9fhv4MLt/AHL2LWbXDPhodsvX2yM2nm2nA/rJZGxlS+sMMPERRdgcXQuGPBJ/FI+DLI2n7c
RMMGmejTzhzrjJ/7ekzL7vcV0TKaNiv8mQ880LNxWD/UTgWOxQ5/aj/sQMm2urSVUMelyfMzIdM2
pbwXoQWtmnSCVf0lS3d2+HUqbyGz5EGLALdPRFlrWEQ+6cEwHn455f1eQYdAE3ENlvdcuRrfoIgM
ZntvGPpmybql54ykbTPI1HFEznBAa38eZcRh2YH+x/ky8GNBjTqYrAwbBxossevBPR1EPvVu4olo
eo5F63AuyJg1vLN9+N4ryqOZbEUkr2lPs2JoEFn0qPaLCDr//UwH1oJF+UuB81dtwwZnAt0lSvsU
w0/PuYbpLP5Sae6XjBJURutspVUOeyEZbR7boBZGQrxATqOv7vhgwKYHTUcCrItQyN3wutSy+6KH
HkRIA/nE8o68oSxKk5QeiFRKIcmvga6yXpR0dMmuL0Uvtr98/b2pjVCyois/RVNTtDPUR0YXnI2w
Nk5T7Rr70Rn4QM6cIJ/Md5ettICeNV1JEijd/sg7CK2g0LdLuEghofnUJ1oAutG9qEXikpMIltdy
dC3p81ZxyaE1tWkwR07MNOpN5zG1KBiR5Wok2K80pJO7sUMEo//3oAEBEcmDmwHIQcTkBHLfv2ak
LudcInMOlq7UcWMcdaQ6PRTv0V8wDX5YJf7t5sgzbBAFq+CY2tMmOlJyGGjQKBT48gY1h4+3vjq2
q5bqXsDXW8g/HzwiGPlzaT7ISB5yKLOpZ1g147xhp+yDkHhxTa3ej1TkCV+gs3usPC3PNwGnYbb6
XCysH14Sp1YeQzen14U8Cz2rZ/d9eYylPkj+kN0jMm5fzSDSMqDckvdXxJswDTB/LOILqVDkEBBA
HgKeJmARAP4xLWI7kj2RdMgjggAGiEIccLlGA9CjVS1w3Nz7EiDhmz+LfkhW7sJCgg4FfqDF50G8
v2jD9nG2gbmFT1bU+RuyRgjIxLywadRUBIqN7ihq7VccH9N9oIBbzB5KvWM3eDO9WyaPVyNgO3Qp
uDo8PhHZXNX14gRk7uE+az9XHB3Y5Ljvr0a+7YJMhUTFdt5NpKma/4+LMhOS49QvxerpU7vOLt7J
WaDueKsfXNt3lbZWgGrGTBJ7gXhxhlIhrjCD7Y50crFFVCd7D1rHUSiGtxm9jclSZF75bqP4SowM
PUyA0xGe3uszx3nJ+aMkmEd60oj7GmNbSWj2bKN4/uWWbBxJQzhPh2zBxT9NIbXdQIVyNSQMUtMl
RerT427tqfRxk1ystW4JDCZsj2nOOM2gDZnHPk730XiIiyNZrHNBOrtMb5Raed9TYYQY/0ZsrpwS
p34K+4MkvKfluE9nAu0IUrhV1sJH7pruhyBbNPTcSbljGa9Ca97Zn83sLJ+M0SGmgjNCNQvoNPSG
wyhSozr1KLbHqt0++xIiBDo4fLese9KDDMBa3ANXYZOK7uHf6oknnB9pQ/Isn0sVfaOVv0s0T99V
ysF0DvUKIHHVcfHOfqSgFtobulNa8GuZebjg+V+G0wBNtl0BDFA5VlZKRdneQyIIjIrCXD2LN6AK
zeYgfye1PKVSRmcA+fkC1GjWzJ/T9WKT/u8gfQxBWcO6D+JoHDyXmXzlxiu5fMKkUGj7ambG53AV
SCUvgJjbSj5cOO5UKLskqRV7wHjpfSC5zQ/QLyHYTuUyJYQcizMW0MJMpHxS540oZ8GPcyO1siqq
2WXHXDr2kxGB21Kbf/PC9z2bppVcp6XDoDSQxN5VGDdnfpY6ZmQUUHBcDlk23UXYn8X+KEoSxQpc
oDSDXMvo7YM/JStbSx0xdQHkFSq0eiRq1GXfN96mzSoBPTfsOdWmYsJECsYFf9/zErSMcdp0l1o6
C2rrOYccDZrsdlg2R3fV5AtMFf8Bd3Zk0VEkwGtBNCctl9c0kD5gmgLmeqrFTlZVQv71UMEzogyX
wcrGqsGMeWDTadyP4UM03BAoOPAdUYhSnWPt0ErsqNYssHLzsTbXnfQe7xESAbDCOjXthCtZLvKg
7H3j/9CtG8q5/0rQmPdmxgro08p2BGqbdR4AuaIjQej4Tfh9Eb18yYn3KOpD794PE8KDlizDKcFe
ZzYIlNxPgGfmCiq2eF9V80d+DwT6UX1wyB/5DZCgyXHCxJFbkajFIBD2c9+gUCENo7OpR/1cTNhZ
DaNVMnu0cXC7RlelLzNxaSF08ThARB/i89nPH+UgjY9462MVfl7LP5xzhGHYQk8xV2nN/mh3ffvS
v7hZ5Knx8ZQzGE4tGLw5d+WxhfFj/8XEAGWR0Mi+xxeT3Cqumx+V5dwE/EdXqjsydkphMu3/4sUG
aVGa8fXjKHKbd6drfVkG+vA/k9/XI+d20RE2WQEDXRVXP5odpv4e1e8n8bUHJ6z++NSfvpOQVNEZ
42Fh4ierwV74pHVjYY+vxwHzLf7YMRd4r/uVLMovQBuHJnqnrUHLO4W8eVctNc/sPkxy2nhWHBdQ
uceSqqhdLXp10XHv6Dype3Qbh925KjggEL8uU5RajZvB0bj0zUIf8B5bjrDp37bg15iNB9KIriQI
oVsPhMN1yxs0c8GfF3UM7Qa2JEMXBdll+oE0/Ehh/EUaKCn7k5AulVg4gZEt/whW4fPgJv0Jo/KM
PPf39nxKaezKYhcTuppmY6D0B6KkSq5rIhMoxfao/gVf6FVLFRzJz56CU1nbmk7k4G1a66z3hMJQ
5Ei9HNUFOGH340FJ5VraCMKPYBEnD5F+8boFWOf0fvri90C4GEk6k/iDW+ILz0iJCZrX9dp95dD7
ZEvoDB+OKE0ircw40ZutAlAoh7YrnFv8VjnWJ8mmtAlK8JKOXJsWjXvQUjiL4h0Q7y5vCZ7UVIQD
DLsc8bowNV4ufPTE+YF2SSzT/1GahY2wh8JxQnkBxfEgQtjOMweJykMNzpqz5/zjjkq1yhINMeq5
qqtbDnR1F5D8BYmmvoLRo3thnpTa03HONntGV/L+jca+MVpqHOf9KWpNLPGGy1k9CNje6pl1Z2N8
eM+GFuEqHA7fEQ6AYec3BNDOliRpp9f+gsYQsvTEeliyUqHe873JbrZHN/+AVojui3ilnAaSA3oo
ajoDiwg6NlLtDKUNZ2pnZOfoqNbVbEZIbX3beWL3P0i3GudQ24gccZKny5rBY1hRCjqiVysIBuE/
NHxf3beJ1XoEgLspxU25xlKOBgSxQhrML5IMkop82PqZ75xiIuaJH7AcH91o/g+vtZPHXRG4NZRY
Vpef+0N+TUgcnF36CSqrh92lkofDPhKarJOglnGTYXiSRYpUoUZdi2WV2tsr9YLZGttykj7yeCKF
1GGISj+D4tmGNu5VnVA4x4+eruH5qyxkwkdgdO148qiSweB5qf+wwLXRk0i0fyaerZlIhaM+0kah
gjl4DOg+kG2zWxyrcWYH5B8h3oJePjXuf3D33XTG898wo0JMIqVUb+zAhSAXL5oDOP4uDaKp1eeO
HsbruJRgBtubDjO0KL9YlHdZhBsPAKaTSwk84zwsTkY+6SSaB/4pCAZ2Ghq5Kj1BSjFjZGsupwEP
PidAvd+xmLpJn+F4WRHjJFkSSIWsUNJn5iW8s4ekS4pzVity6JjoAFwOmZ4JM3+TXSUq8719AMlK
jAHa9CQ/WRh8nBIfllPp/vGeamM9Jty3RqHkbHoU1DPMVnkbRaYoPLyBfhqUkgzsneJp+TwgYjWm
fRptA4OJUWL6lKjSd9ZfbpkNOF9ebPdjgrBs5xlcI2c6Kujs+YJZPUtCHBRd00KyKQxCh3hyFSSs
N4ovvgTTYCN1lne18STRaT5Ktj+IisZtcZkuuyijDQFKO/OuZql4gpOekJJzBIpS+57xTQPG+Geb
kUHv1EenTIuvxBCUhPl4pUFVcfb++K5yqvnKtZ+oWAYIJcoSyESGkhCYdte83T/OU6cxmT6/AbP4
GNd1gKYl+A2ClnRZ2nISsbnsliGfyWOnMlCwcgMN4ktvvI+UtLF6MAeNNtaRUEvwZA7wWuFTmS7a
iiVoMNI03Gyx8MBUVe/6Vm6xMDrG+nMpRI1rrsXCgsqm6vXJBrH5tP148X+gqLw5UVEcqnpESkY9
TBm+txwvoKoNWTaOGUUgAAqHGiIEE+6e0mYxxJRLZt/oi0npxuSL3pPDxprwR4sm6VJ02A1Swr5t
NDt4klnmuaTTk+3EXjgmcOFKjOnf7reXbtK/IizvfIovWMy5vDrt9Xg6f44eubP8idS6i45n4Lmb
PCm4kBfltZDPHbrrVqohjjDpg5Elx7LSsr42Am7Mcdn7YoS2DsTRP6YgVCb/sR+Wo61x/BQUeXDe
pYM0uChUwZDngTleXqk+P4bMD2q8cbwUfuYqn4rop1+g/nU6Na4lgHZ+urXQtchVvJLCJwYr1QeV
4uwR9kklXqc8mBfaGKMEpOIwQG0Wk+bYgWN8KS54uyR/5x5ucX94rO3MGDJY3FDL7jptXIJy7tip
aalQKoCufhHj+TFYG6k8X8bOC9mCjpqiWokEATV/SM+7Of/YrtAoCF1oHinFFFIrmW3/tXnstI8l
yJ7YSL4aCURp99Lg7mVfMNB6V72/+4X1hJsFzSzcIWGv78npd+2WcSvDylXAGL/NHbxFO/3ghmu2
qEp/vzNut0AVNtjkwHIMAYEV0Xwg1WrOA7XDeF//7q2m1yQhFNYeFg7AUKdTilPKanb0XtRBNZE3
OPdrDqygRjLIJfhnF+xjCiBSg6cXgJMEEmohG6vc5qieFATDfMPdaw5VZFdugKYg3AWeOuu7tPIT
vdt6zu27UK9F57RkPCDMVaLjkxxn/ww6UggbY2WmT6yuQj4OYZ+HOn0gt3NlPjQi/g5ijhDCfDRT
8PFcNHoxSUEdr4vUWk+DN2zRrkUKO6iZe8sPzE6Svulr89o3itHshd2CyzZ7QLpb39/8I3Gh3/1W
LnaNXepCRMPqWHZMOe/7+ztJzhP4/CTrnPOLv1fN670+Wyl1Q3Fq53vHiTv0eGWI5EKSgEjjMwqg
qEIxnnAvQN45pLmlgZqaIB/FG4/Waob5bTzutYXD8pEsZ+uQaKO6mrt44RZjeJI3TWTB849xdLYb
9nUhCHDSjgeveSFHlQO+LbiEZ1ab91y2avJ68I3D/0gIUyI+UUkLAQsCSTtDNwCwK3FI6Yez0HA8
9KQ/bSceOugtiyzb3ZsdsyiEah4j8tL3Pi3L2x/JNHC82goJhJK8FJjdoz8kM1fb0Be8q3jEDimi
AKVpGMIly3+iFkWaiVIM2YkSChNRPeohTIFsPFXHjc1BK0u9AxQGoA4xLaV6/T1TP+FIevD13Fgm
GPMOhmoPA2gjpCjTucPKNnf1GS0uLmL18ZO/Tcp7CRmK3w2hxEjVb/QZqmTpTW0Q11xa4Td1Jkfh
Z+jg/2Lzvyua3fWGSv62/jd26/iUlYqkZjSDmkNwJrmm5PsjEFCdaiB7iKGGk1zpLY6bIQxH1cYl
jpjavGoyu1dH61fxHqDjnJneZlZJIWAJqoz0aL2Vz5dCojvMjx6GwlPYgoSfOcSfTa1w9KjHxmGP
pkhyngrDpd91FxFtc3KvLhQxOYqqUP0UUG0pK0+N14XWquMyyxBQIh5XIt8TFKtOB9Uuo+DftxD9
XR2E3G/Ae/sJtdeL2HLh4gTakHMverZ75Q8hAt4vl3NnYQw4E5x2bXY41Q2waIYLjvTrdlxerNOi
ZLvqqcvmxhqjqWZqo1HtkdHhcqGGBPpelokfXpIzGQp+LmqHkO5dgt5JD1xEdo6a575bv3a9rLJW
Uu+vppKN1pHoihouv5SzJwOFatXASMl5LAA4odMFHjmCyXwMv0G08AnWn2tu6GquOZKFBcgjT6Z/
eIZ0NGqp/qjMs/TPCwENoiyLTsETD8gEzfcC1ey74BP1NnmoYcdoMMjyMGVg95O/9NNlZ9lA+8sZ
a/6ppsHpxycoUgc6/uj7OAO+xa1c4UtNneCcV4rQ+BjUH8RN3Kc/Uh0w5OC5pf49kZs7kTsJcnTr
4Bre+kueTnPee2GSeqH+Bxo7y4b/YZe2xeNiNMuuWurLAyUYV/IiYo0h65/VtDN6LPldg7gHDf36
4oA2c/iIUJPu8yY010Wr37WE5x1jyqdPj82OK7E7iNmZJB2oumWAAZkbUEkR1hKnIcQiKOK6BHO7
LIvrPVvDZy1bS+AWQxR68IOWkkqitA9PW4JL9TLhlBhgP9mx9obk2ltQV96udcGhOX8i1mN83seB
MFUKU/MlqTW8aq4iUQnYAzGPSPkxVV7cBBL4qYY6nnEhhzmy5tL77BOpmNfbH/sgU+5i/qO22RBg
S+aMQ4WG0bYFJZeNJc443vtATL5aDmMpVP+/GtAjZaUcb6+ABcNtZh2i6YLaWQ3Z2hlxFno3xVr7
+CRYB0lGBTkLcfzsfSIYoUiO5RRC15r5koMARKCFbJK5u+CzBkkh1XoPIuDkWn6XyLA38RsMbqKK
j4Tf3lC/ytlRL6L7/bzNovaseD7Wms3kJf4VzsO/z6USJIL4ifRsP5WbNX90ADzWx0sjj+aw24Xd
7ABJ1mHDLnyTT9NkMBvhJnOP8/it0rX2otGCEjX7CS5Jj+ssJqYdOeSEPIyDHMp5sXyZg3pr3oAs
wOdibHm6g2m+WFOIlvxCZIPrduJlIFxAL2F8pekzMJh8+EKW8+LpMVyycvz6qDggA6jlpJMt+2AZ
0aoU0vor+1FQiaZZMUDQNOjLPOZEll+PC4A3E6s5gcyWV6uyutd+otEe9HvNjXNQmqrQzkHdk+Nq
xNFEMVYUip3THD9vc4FOQwEPdghwri4Nb3s7MkBOYX/D6YPRb/WnPP8MAOwGq1YhOWIgCXvjRoLa
IbG4zWeUA7qK4NCYacz3pEv28H59MfaLOl7CH8sFkGLRzIh0CTmeRAwrhMEkwP8PEo/TaqVarAIu
QYGaUWqVB9mcxwN54wPbwZfahG8C4TsDIPMFa1BBSRelbWmcuiES6jFvXpS7XmhHPXQG2+doe3N/
vftFyvwiwjycOmu8azcCQhY5hn2VUQqM6uSkyVNE8ZJ+VzAonFJ2uB3pKOkCr4xs5b6O8y3tLDfU
kYPQZtK700XrBssskwIhbf7+uroSC1p6khnvluuBIqFtAPTSAP1/EqeEU32WYTFPxXPVgAVkn1DF
D2azhN6jOcLuJUgLqe+NozDCca5++Ub7TT0V/hnZkePFrDrx1Sv98EAH9M53LkTIU9U7Q97zFTrM
wmnsXczYoZtST9Dpq5YKfjNlbIYeHqTfOjHuNJ8+H0NazZi0JRfIxr8O8A9WpNkIF8f31b9bLsA4
IM2qnRwUuelXEVKrPQhEGQ7ZuA/lqeMjmKKEWW/Se49W/eQfMDXxWV6kRoSSNwhfnJPpslgo0/Y7
DSW8df6v38ZMU0/+5jl/jhveZ5JRaSEey1Y9AVBU3gxz9W8JNa6nEXo//Pef3t6zfb4ny9hyh0/e
kMzj+uKKQdHwGV4R41Pv1xkdn8kXSEmatK3MeJdk4WZ+x7a4H0tdKToUoeSWA4GDHO5MyXgpk5jc
CiwDBnYa9GklauMxLlSpNoUAtlwxX2AMbkTrLIRhnalO9YXGCP5mWyXn+xTF6AW89WmLpYjCv7Z4
oVucRN5B3+yfclTjPXBVaMO+sJd37mreHprc9vKaPTeULc03CH0QxngT7vz0GcnOwzPT8Yl21b2C
uWJTaCpDRNR81YgmbfeaR1QW2PmRrZRzJjtBdXTtk/m1p6anIvuQiRQokxXuI/CDTWEiJycU2Zp+
bn8F6m63Ni1+11vz4aymA9v/3b+tPlWxmC0HGzqz+mrxxWM+3ZN25VTEeE2cDzA8hYjI5EoRg2Li
yDO/q8tsNJN6thXGTwD5wJyGK+ejxqUCOsCi9eH17kEz3yzLNI/fGZCpn2ifA5QkKes1GIjuCoZe
8xMY4xXoM/SmQjw6hxTp9xtctXh8lkqUGYdsA3u6NYUnV99YqmJ2wJ1hM0BaJcwY8G93PnfEMT6p
eC3IduvH3DCnlTw6zuYcypEkLSfHlqZLosjEwxoMyufMp56xP0xeHNfw4Ux3Bcmp/LkPUIDbRl5y
fWdlYHX6i1oLcCWA5XGCiWMvQfEScnztLPCKoQYX4jW/o3TSxmQKF/K3TSfg8zud7VYjVs9XsTZ1
cESGGkTyofMdwH/vK4/ecBoGgI2OcyfbmVJpW8Us5NcxtuDlYcip0BEsozaDHlFKlyWTr1AqUKk2
RQ+BuE127DK1pUocsRxP4BTaFJ2BZ5Gi/+Z4LavsiupYqOEQylJBMCOlctFjwqyEnkb6WewEjaAa
kdV9vnrVwVRF86pZkLwlGItPqp0GxQZM5QypIzQ2mO2eLh4/w+t76e9Vg/baG8gzk6dF7I3hVJb+
Q6OQJ+guc/TLURWUMBzS76x/AucpyahYeVPk2cXai3KfmOUSuu0YEnSjPN10IfO54hvI0Nw+DVO7
+9OXhINNMCf959yQuepYG+fUZgTNYkwhENlbu7hZXlHhzSvsVRAddJAyJXIFs0eX+6fib0j5zRs3
FTyov16NS5cHc4Ynwei0aEa0MUgdgwkXWE8Fk6vhzxNn+TVJanvFcq5NIaJHAkEtrDsP8qj0GDS9
ijS1FFpMq27dM2Ew6ysX61qGg1THjXg0j6yxVg3lcfNcFzISfgeDjvr05i1hyAjx1pMZvXxXjAtY
9sbM7PMw8jdmGP5EpTS+Q2pIXktnRbfKMmf3GFWVPuG6M+9C6tf/MKSTyQmGz0LU2GG8aeSntePd
Gw2vwX2snWOu/QmdzQKbJ7ubiIPnZHWb6u+I3q/Pu8ggNtSd7hhARLzfspRJZSA6wZChyYn4vNUT
R09ZK8763jD0rlEBBdh7LrwNw1Hl/jcdrV2ne/EMSgPml5dXYDgRRuLkNhBhLBSuv4C4RZcPVrJu
CJDdjTEJsgOe7qMae4WC4LbeyS8PVApL7vhadaP83STaC+2R8mLA9pbO5USbxxSv5F3/YfqaxXVB
/1Z10+KRdkyNuGjhcNeCgcqtLi622YR/gXjz51mxFFKac+NQv0X9dxpKskhpfRzvrHnNoaY+ENDw
fdWt+1dMBusuL0mZ22H9QQJuzY0PbbqZmP7WEZjnSUlQvcIT3YtP64lShlYjQ/cn6TaR3YVFgrVz
6SUdXDUgO4zcmJOZoOvhLYSV6TGU4zFFThqeAz5n82iRrE6qXMytqNtJ2aXAfK2UUju75ZDkvh2a
1s1pz6/do5Q3JvOlTDmMgWD/PRLdh7uqfBNrexudRiSXgf65ECrtjf7h/QFwAVO5P8kav9E8Du2O
812/d9mOoMRZcjLTvosLlU+i6CUNXdY7x2EXKsng7mFE/JvXAKon1ym6BglPLyxtwUeUTuvYpzJF
ZlnYh/rKafUri86Gk7YMTYJOJcw4Y+DDbu/I7oVqIviUc4BDhcVSLOK9RwBnxZLgFZB9Y9FPtAPg
HniE+YiXdRTJQXZ0qluPPjcTS2C3cXi72/r/ePvrXu5fHplb4hV2nB6gjwe7mXQCjY3PBGTcuXi+
kLU6bnScV0rS4XvrY3lBvbM8cohSyqT0/MDTv1dHhjZIwvUPQ8NxDnf0J3a4LyDnuMQYqgGtkhCP
hlbWytiKg8Q40pE4XEzKx47gXoxieZYYeFF2CBEako9tWxYPf9wx3vXk22cGTKvadeyOtMMZXack
2vXp1eGT62YyuL8/Hy+h6zT2fXrE0BQTqOXVi6DzuebrpX2xAxo76/E1PwCtyK9HAwG6NHDF8byl
lSipSRe+4IiT/kueVi39A6sKUN68MZ4JKsIHGdsn7Y6eoG7WY8BDHFqUpwXMiylK2u5Y0NdPinGZ
yT1PiHbGvZO0MhRog5F4zjzs5jf2WQvTmz4EJuTWs+JH+Iqi2VE5Oul9o073rCV6Z5Abv2X53AeS
VfcybKZMxhMZZvTpPW1DDPqKfhNl18jet/KwfQTAoXf4XqOQLrcxLcrCRu4nxtGzMPYPZEYldSla
M2d7In5qfF6KeyK2XYV6Sc6BHnk3LW+SFD0Qxv2VWYeISK0P4iMLkIEHBmJjn/T1LrYc3IIHzNqk
Pni25jP9UBhnA4GL0nHHINOlpdQlczXXHGCok+3e/dGs0OtGyWlITjqp5TqOp9fq5KaWbWmJQ7an
N1vNrjzUY8+TAVXWBHXmhDUf4p8ky2JWugTgpX4WeS5/BTjkqgdguknw4weXefowThUwQP/jZ7Bl
Mq3lS2XaQa7qLenDtfACb/zldlTCHw+B4D5UXOx1u+41gChATHrBM6pSGauu42LBIQvyBEWrQ8nv
9ZnYZxVoIoyiCURWRx5iUnqk7z25sIDDz1xIS9dTAt5v/2I2WNTE5O6M9NH4SEKugw4pavHfaSgh
ABgilCcHydznokGFIEBFssofwVpciK7wW8F+/R/42FvGtbPByTuRaMIR3XRsfflFd699dcwJ6O+T
TnblO6THocNUP8O3Bv2boWhM9ACPFVahBqcP+HQgPOlmgI5PYcBUBTSG8MfZFBboA5KoeWsJ/tjC
JieXnQaiWic8IFusmC+4uIwXpwzOTmoiJZx7VJ28cCQpQ8us0BYUFb1WFxH3ZPOshvguGG9MNZn6
aLYt4Lbm7ooB72K4PbB/0kUuE5Isc5d1ub447ceGirR/xmjzjrpTbGgwlw8zrrNniXxpS/e3KUb+
o3+bVqulfJZaQi7uB0ILCa4qIyJiZrrnqoZgtDGWUVTImOYeAsIYHheQAorGcVcS+j+aFa3d7A8G
2XNH/BK5TEhjlxAvOxlK4RHJrNe4psUaQWliqsPn/DHBXmNFzL++yOntFD0SHcVlexoyQ7OdObO2
IJrhwNoWJOG8bF2o9LSFoA6t01MZhGBmnEwEfomwuS2AgSR+PS26NXmTV/otmKU9YVI0FKvaXDfu
7T0e0+tXn20RtYkS+9k0fWG1zbh9E3dH0Z3OSCSsmBFsq75TYsJjpGcP8gekzMhg81/2pTrwXigj
dlXBdW2/F+L2UT++y1UQR4WWN6vGSMCvonho65cCgvjZJsvne8eXEqKk4bZO1EVU1Yaj5fgo4DAp
If0MjB0KpK14wrC3d8g+u03itTe7aWdMJWfoYG2/Qm/Rt4aUDlBrVJRDQKpw3XbumxWiL51nvdEV
zXIPifvjfgo4kaPlnNdzKb6SlvpLJKReQApVtmWCtIU+051oZsb2TfxOMJcECj5FWA0lkQUR7aDn
NH/j1hsT+6KrhJYpXbRydxzJTmqePp+hi0dGIEghwa2Kmgn4VoE6ZbGEduGnAOLBciAyhBakzJwN
1pLYYdphM9uuynmGaXXuUlgp+w8V/uYQckc9cZc5RQk1d2hNOjFVqvPlx++nPSKfhB3vSVCPcrxL
KpAGzfSTyV2mUN9l92qFQdVo/C9a3tetvV/xhfL8t1QTl3EZkg/muDKWx82Hgv3twFQglugAacjD
NSHIcQEV4QpXeT9wfKcD9a9L50R2uFuH2muDhFeiLl2JiWTpgAyTtvVp9X1AoMKXw5IdQC7eOxCP
3FV3fxuewynkhq/DYm6ODx1KGAhtKaCP2oYchnP3M/bisv0FfEEkU1Ao57pU8/5/iIVsMm/mNTmD
8txjHJNEju3DR6UeIlfW2IHAXrdUA0fe4N9I0simoeVKcbry8zTMzpnpbqB0UxUDAJxlsn0BnQWd
gv4PQkeBelbV7ppR+McXbG0vj9ZrejIzBVzw8l0Ky+tPbup9AgxLnEvy3cneqfTUTAyrFmnBDCji
5JVoK+cVhNZ0KvDrtWZD1uhBwU9tn7mZeJ67l81nZrce6IgMHrWzKrBc9hcjgyHp3m3GQfvMiLbp
V27xhIz6cN86XQsflYbmVUaDwd2NYbFcBeW2d30m4THAoy3YG7/7hrhyrQKaNPsiBzUm74R4uBSe
75IEda74aLqNs9Zp4fwyi8IwSDzJIQE8RkDzvfTXyHDIPgmgbsCj53jd/zv3mXSYN8yzAAlIJGoV
OcG/qVBObrYOtEYdbV8Zrz0b0XT7I0Lm5V45ikVat3ZMDWrZndAAGL3caHJhfII3ilS0knXxWRkJ
Epod8lsZ7yWfP1JFC2mGvrUjrzL4/4n7ObxeEaCoXhWUDWE3nvfdITXorfeKLXOqphWvXi9xhoSL
36rS+oqmnolgcz30YOKIZO199OF178Efy8fLkaSUVErQpUqL4yRPRfHtzWO48Ivv+U5j3M0Wepva
8dyQziSCjT4T8byHwE2rB9+D7dM2H356xzOmqrB3G/5Khf+SwVNkFBL9ysIEWOt/xxRaZi4MyltV
0kL+Jo6owt5RGLLRI2kAJQyRMRhKHkrRd5fqa3+Ii1061G7dazrfIfaoLKqCpX+0QJnuYPntoXGY
QRFsKX/nGQuX79fACR0P4NHSqeGGbD1SH4ABdOTsyoMWbqDJjkYVS/aOp2xLGVDuZ04DDluVNtHg
LMrtCbUV2+z69LANXPO2jRlkXcqnQNMzFRzug8zIepSVHTW87qDUwvHua0vWY+LSX2kAhyZESzVb
AukGC3jPx2nU0k5GrAhaoMK37/ctgZBEuBeigSAwh6DrHnYGNMe3TTRXSZGV2sFMrI4eziLlGtbx
DU+hrkBoA2AZ8atXVFZ113qAhmvIqcCcjhHnLNTc7+SfzKQWbQOAL8psQS50mwL9CG5WBEEK7Rou
opGl6157GtudFIS1nL1BA2WH9rTlWi6IY5a6v3hi9Z3q0RDYlkCeIHIY09LcvETQ4Zjptqrxt+gw
l+WndFqSr+v+3JK+x5cqIz+H1CAobE1gk61TQv8tMs0L0h/tHQTqBCancJ9mLDalxRHTPp61XMN3
ZcaRfIVfVlBBExzTqo/cGKjlgRwY0MjF9IKgT77TiGxMCIi0jBnu7Gf1xL8ekql8zbTI01d6yGMY
4UQdNy74opIPLl7SN0PxL5XB1f1wfBjMKTUSTgGudBU55U3gFEoFLs8HA19ng4e04VZaVTo4lAOH
0Pc6/lFyODnSH6FOdjO8bBs8kUGgct/RHDWPN9/3HNA9SFYkrSe6U+fSJdk3mSXdlGt2BhIo6se8
DZmOh34vLKDYTcJPxDqALR+RoAUL5ScIb3HK8WRk9EOymhq7rXUgrRPS2iojpLFBszsYkIETBifU
VqNxGG3pZb2+jh0TTwaVz7Vd6IqTLJkDl377v8d+RDIt5KoryjVmkTC0a0ThXdrtBy2MbjWI/cck
qDGaJzIIa6BEc17aI99ZEYfbxjTpFRNIucBC4POlRniAA7ghtwD4Wu4e640577VMRZ9VPIoWPj55
0RLPuqma67OkB8aPzgomvEanC4F/tO9AMTVS6SCS/SYpqYPHFvcc+bOXUpHH8OIlp1VATCHAhLz7
0Zx4kf7oBICPQi1CsZ6IenxuoeN+Uz2YMbm4gD/sVPkE6HcNUCma+elSDaIwP1kmi1bUfb1DEa4a
Gjxcd5WKV7+kEgPF0h8wkTYmHz7BvQQtb9/+LmgmxeRAf2N4wZjXLp+3Mce3UQCafh0VsOZ7dpkW
T4TBrlODxemTbizxQoaDXtm82cMhKo2kfK+2C9529havpcGwXN2SJZBypnYw2T6x6i+GbDv5CjZK
nntbyecgR36ZwOy77tC3zWqdQ10k3jbZUQtNpY+ODwNjZRd0cLu8KGMrcamnlcp6OaICQrzm8Rkg
FD8vZRzUtqzV3FOyq0uDWxkyfoLULG83su4LBbr9pL34rIz3rjO3q3oM2i292ehj2gZ5ViIqKBX8
bwsE1diwsqcRxtOV8/Nt7ASbyD/9RF+NS2xEa0klL9BTmVh4sn2rVxY5DU3joH0yMEb6ti4LVCB5
m9YcvRYSVRKyYuMgRGErjxLUFIyGXJls/q1jlsc+jqSUYelNJYGPRtp+IHNFf4K5zqBDgttZHyJ6
VYDRd2mprNO16TMq0CR4zKVxsFirrQ6LpG0BbLmBC6bz1QguLpZSCG/fJo2a+qDzvuAdmkEL1sYD
DS2rTqMwOmLkYMINmHS31LzZNKqVk+RBariQT3wXRtKfxCkK83uhSPFPresVn+Bj12ZhryA/icqj
YPs2dTBbFzPQYs/08me7Cs0cq9gVe3wsWFQX+Ln954Pl/TJ8kSiTZLPfu4wtr7aQmA0ck1fSUmEY
tj6d4zMWVkbAN2WgRehMVrMZqv3qZnOiGKX2otDEyF2gGQOslaEyleOCKkR/4rBXOjsDbG/DOpta
K8lt67ilHMduyZpYxOIrEW58scZzG5Y25AGQ/29jakONA//TdtEXeN44ni+9dkff8hGosybxhWHp
ktRcU01WvAxWPLs6quvPkT5LRF8tvOXEjgW0xnIgwseY9TL/nHktPc1TNjSysRjmM+IU8UNGrFck
ezITp8gbzaaxOxW646zhOkwxERmhaOzgrHU0LqdnuwzlDHC4abkGPOSz2QvCjW1Be/piz5mkYK6v
YkLy6U5VFYwd6Mwh5mDBP6lQ6OFAHuCjVi6rGNcN1zKWk4oZG+SAzsYzwzUL/GhRUf7hzWgdvBtp
aIVxbvRE2tj6dexZrPAA3ngLv/Vd/Wlf+ud9GNBHvEJMKdj5+DDLrx9VBBdUVVM6gzdFnwJ0XWYB
qNPsM9+zKY3pWXotqAcB7MAolBM2metOTFM4szA+c61RL5rge0lLwQNqWZ55KDl9r22GgNq1JRmH
phD0ODyfqkSxE8VIn9Tg30bwb7sRqnse4/8mrsOwpsB6yvAYiG4sxQMgNbcOagKQqi1t6DXlnzPR
bxDcdxZgLWGJ/ILKargPncWpdUbNpDoD2fBXpO5xDpn0e1ZPWKv8HSx1TeLtFLZ+4G9GluFz+i44
DScgTouwPBXYarOgvKxLCzujuiP5u9LhlcTLCBJn8tzkQ0/ErWTVJLKFKjByffinpvb8ZFNsq00f
Zohyv/thN7QBgYSONF2JPOd/7ITHiyOq/QsZ6yooRj5e86PGJ05bJoZiRdmQxQZW4oqgXyePWjh/
bQzNmzr5rgCAemWQI7ITVX7gwh1eaxcA29uvyIEma1FUTGk6wRZiiGefxbfmv+xFYfhPlyKE0ZbX
KDiLbF6eLa5Gd4ZNOkGisumdF3OqgC/8P7gPvyE8REbmCR5CNxcpMTEtFxfAUfLI//V11Q9smoVZ
+pXEilUAVyblIPpmZMSQ1GQkRMV9/2F0OHioxGdbSAQalI8o0DnBy/6wr1NnLlVCiEy/BXfRR2L4
BSTE3QMqIRGGFpxvGWvENuGIPBNiQTP/M4cshw0XJ3cbjVnvWH5O2ZSzqVv78TV3RiBS1IsiAzw+
UrnxddGjRAQMSSwKI+KJx8uf2UkGtInw24F6ttvrJEd6hxcuh5iMuzrVY1K3IbqOfg4DuS4c01Gs
SOZD6c08bKHXpjH4LneB1+1xdvKKE69plZCSom7GfLZmb/tmPEMGDHGaDcFRwMy8UZiKvWUSKzwS
8JXjdb7lJ9ohRAhGUkd/dOd98SnsLFti2UQWeDqrpL9NA6RSd1/WlALij386H6b3VMSPp8xHZvZM
U34OTwld3wveTCLtwXogUAs9TkZK8KQ94MSYW4/Dznb7f0h1YtITnTgTc2wesfYo5nO8D06RsEeS
awGS1L0fg4+FEr3rFDxOQTZZ1MmGsTBzgsHPrb3y7CYwjRYSSkykr5Mw0XRLh4qsU/+Y/G0Dyo78
BtPegE+eiHUa1mJywAXBi7uUqeksi0tOkrHo9/qoMF7pfhic3hq+j2qkTxJqu/CjBVAetPdCheHM
EDYUXDzKNu6CYw/4P+pRqvr7OF6YjOT2O4bEEOfXtiFqi2kjHr0izgg8DZ2DdaKDbvfxYk3A7V4g
rNFrdT0QVhaP0bSp20PpK7JXFqbfjA77iyVDJiS3h6wSYFJCtJmB1hGIuv6bl3haFocUn5ld4ftb
WAb822b4sAPiBjfkUfrqBb7ja5dejG3C89AIt582DO8F42NgftFJpFZ5NEDpVob2rzyDO+pQ39kK
L01VQ3ADaDH6gAA2ioLbI4qOIeC8wVDQmNNI3/s/0EeckH7OBsV9kS2te0B02Nd0tUlqGpf3LiOL
1X6ScqZuGAs5jPqn0SnaUri3TUmDM03ahLoKZAuFtBH/4sp7vF2YV28qctly3OQ/bynWPRNDm1s7
edi0aeoA0cd6aS2ymSG4YvH6cq+NX1RVrNUYS7YJGPUu+cld29E0JP7aKq+wooM3qJdrB0Um4CD9
xbCP5/aYX52OHac9yWYa2UKCIvzNYGNga4Ts/evt2ceqAvvZIdnks8yHVFZCcSqv1vAPMtQyRbOC
03askrNwJaknvPIm8wYOh0GF3d9fRhBI6q0+k+8QEgyNlKM4RJ+Klj1y4+FnH8umoLlwqpfzd0m3
8GCeTVsrFu6iVw4wDQurH3usJm4gxos9ALyp8kGeBISAG9vtu7ORp2Mdg5JqmEY+FVZMulbINvNA
BoLruBoOlzzxrXl5rtgRKmJVzWvF3+KPUPVkMRn0qsVv0BDrZYh4OJ3M2M5aN+gHhUoMNTiruE6O
dYjASSv6/8VlGgHt8REIqzIcGuudZgjPdCyW4Va4NrCiMd94JxJlVbVksJX+5zLsvaQDMPd4v/UQ
TFppFtR1iuQ017AolV7LaxhSVAPGxxjMmizaOn5qSHZoy5OCQieNBMzhUaSt2x7m3oWpv4eCqUgm
3Zp2D/AJPJRj1eAjmZujV6SZBkzJAhIdqrgu0+ilSjylOZpkCZUdFFAzpV7RlLU7PDkrULM6F9+b
VIbBxpzXCCOu8UyVRJh6qza6exOdbL1dkmLdIXxFCtQ2SvEXNrwEo+gTZk1PEoTLsBJW+3+AIIUL
dLR4QeLz+bhNmKdTt6vZrz9vrsbB8Nf/FXWURmzd4LnDAldRWEUZSPykqc11nZfklH8FPj6tiIUO
kSAGTyxaKR5N5vAsXUgkJ1ADwkQ/Ya4fppaL1SJb6zoKFDRS7dCq/um/ZZl+4WqjUqBnhxXx4XTK
RTGCjbQ+lBxJTsTgKQg+phrfHQ7tWXDfhEwCGg2J4sreNSTnNAHrCVQFVSMtG4lt5ved+CS2Mam5
9LbgPhQcCG1ligmAe8/xvvYhlH/mbzy4nb+FeASrjwNGcyDeg5IiP3db1XQMnd807fI32QNsrK5L
x6EJ7lycUBbazeS7hptTquX3PA4bx1L3J+rnxkHKPbZp7PRXE6FayW6wdDuEo7dRGhrR6JomIS3H
vbkUzHQ5HLIUj4eycPSTlIEogUHzpyPRlN7EgLNG/tLXESQwVHWx2x2RWI/jCNKCTku+uKQYfR3J
LllIaWV/LxupZICQfd7G+gQqFaTxXv3ITji4+OOG+umXPyfp4O5h9dnQ1fgc6Pd7jhCiptkyzFp6
dN79xWPXeR68gisoIacTEAO13BdAToBYURxQGRot5QIuEXXNhF1zJl2xSxpxLfnebA4XEVMHC0pu
j7Z8B1d3aHZfMyRwaUPZhzEBkvFJdFQJO9AIGM2MLHhuHoKSx958QcBncaJPbBUq8F/WDCE0PxFP
T4kDg/wyhxEOIWK6jjzOqOlr2GLlpRH15+yIhA3jsKSB9JgepP8DgBkagUeO6E4Vo4aXvc0KBQ9g
jBfOVE3aB4eF2AoVJ2qNjW23rvEH4VAlzfWtNmA6beLuwIHoto1qkeAx3tONxGxbl1m7lcYVYoDy
jrHV64MnhXsth8FUUwM3mV6zzQYjQ2o9yFEMmGLqi3sN1As7au0KJmTRPxQrF07OYh+LSiRCdJnV
qQlS2jTIIpttR28VkZfNfYhCreWsa84ZXvrgFSZdb+D8FJ/RvsvO3UoectznlpOfg5QYYoYM8GqG
QirY21VT94eYlBffbEAXw3tWmD9ZWneK+PJJ6GhdHkUAIQC2nW0n5X7MH+/G5yXPky37SyTsapTW
pLFcDYtV/AjQTXynEQGixsI0ucQJWqWaOsXOVvr3/9wBLt3QSFKEw2glgLAELm7yi6PXi0v6AOM3
YG1joYzxH6/xKpggl5+KeMvYohsOGmDfNLxM/oZXzInLTZ+062NwOYLbZllxSdE+NWaEaLlfOp2O
R9THX1l5iHn7jJ5LRe9lU3CspO7GBRYEUVZhnLF7Z7XDKGOmJLwBAU9mhfciXT3LKO1GcL+1q2zc
j6rE2zC/QG/nOVNbSMA/NhXPd513XBYKvvxNQJdmUO/6vOrymPKbfTHFao0VEeu3EPHW3jmaxa7Q
upA+yWsgu7/KGWQPoJcOxjhjV1AkkEDoVQyaqueD94ErFFLgioqELzR4uqSxeoz98v4ksv8Y/NQv
hJszDcNcMeaDf1wFu0twp/7dRCaHRdtlIQIuw0I636i1LIqhU2ul3XPQlcyrD4Lnv51bsACVstFd
tUd5YSPx3CojXOoLuDznDui/UfpirIWEqjMI58AVC24bWpIcMtRZycj8fq7EmN7QzYwG6AvjKsfY
FIjL2AyVqRm8PTVBVEVasbEiyW1BUDJlCjR62sRthQUHbs4d9tHtiq1yPIy2aVeMU5bZ8VH8tvzF
ede8B1eDvAfSOJCMqmXJV1w+F16fYhXujzAY/XL64QjXPnFSwVFJQdKwz0ncGcVrQDPP1s9vVlSb
bRn0Ou7ykWcSlmYJmGOeT+ouaMnli9k5brT0qckEHDyXLpN4qecEyXzpYXOTM/z0ySTuAOE1xTCh
eHOgyu7nYexty+MztVxOI3g8YJtvuGTzwUfQEa5oSoCXcGHnd2K3zJsEdMcFdYygOFTRXCIUyk3z
4GJnRkM82x8vC/zljPOcQTpE5IipbRW6RY5dR6F1JXzGPTOHnc87/6eVY0+flwQl96jp4rqdlZj8
fdQTw8AZdpUMgRRsBJF96+2YeNO2q0JSOFFw/H+m9m+r/kaZ67Dn68/5BBiqGlnhbTN6MYh4mlmm
BbhiPPEgNXcKdLkqNTFbUkiv3D9x/RwypXvs6OX43yzgMxU1YvtECn8WUbSN8jm9p9dAfeLBd8dQ
iopOzpjYLCQzfBZY7FISRYq/ULYIbJQ7wT9uSgi9VEuPWZUMge4aSRsZdBH0WDIpNTpIpmuK30E5
sqLp/fU+uZYYwwU7umtNMOh+NNCWfCxbVyxYPvp2d0zhp5Ttbm1z0Xb42Pxr0y7LLkE4SP4gKDgW
ZVym/KVbqDY9XpXr0W9OYL2kXglPSQx/OEj3OitRXhgGBdTT/8AYqpU5WilfqzK1n9G8gAiPDONl
2k3qM9svUDiY9S4TI0U9oxMZOqLZ6MwyoJIt0AqWcfT6Y9uo1+KZpQenE3uHPsHZi+eiNTGlqLyQ
vhOS4h8I2g4QfG6Se0PEhjcuy8H+NqpQ8PsDKjwUtEyGFqnXTBurBOSR7QeNYnm//HFsg9c2yayY
C87nKUFqBAuTYypCu0kBsJ+kqOazVTa2GAwLhuVRYsXKaQMqeb6LxUYNA3mXipqbYr/blgcLLhH8
CCFUVLx7Q8fPDmFWnZWtGK2MgAQYQirS+8y1nta+zKIdYilPK5G5lZzPo0+gAXPNMbaJOovBzCWI
z+2cwcKoj5HIiHksRzurhTlUgNqcaw4De3Rcr0XMOavZIW44GHwf2I+5qjrJM6LOMTE6fnmFqnHM
GT8ScEd2cfofzDm2vZqHDIl5w/JbRNMAJSduieOrFd0BBLoQ7+1oQUOjNlo5CKul+LrMtLFbmzWd
KGSZR8iG6Qm/Q3wrr27unH87FH/J9OCG/1aMIhJwG5TvdyxHbPv1CnREHZC1uLfRtKgjx2dmUpMs
acclcP/K0lhoEZ2tHuJkdGFYGz+9RbmZW/CScBWPNbN21rV6HEP1Yf3ZFN2SxaXz8FRy/uMp1Ba4
xuASiZOfWpT0RLMlsYCB0EE/+ch8E6bPYmaBIDk+zed7WNg+UY23Z4Ch4GPPh6oidBPGhNBmspdv
/Hfs3bujv9pfWbp0BAwFB03eTarwweP8KzwnhHbAOs4jSOzK92Z9sUBN+l3mAZ6VdqhXdAJFMuG6
N6V1OHcC82eXEnss+9xA/hvrUaAQnWyxe6FKMT3+DW0Js5nn+zmxJA1cGNNsIS/1w8WvRpSZqTpt
Y79drTZ8EV0dx8KhDTwC09ZpEK4ydocJ6TZKnQgC7siFQM5zBp2fEZTNBCbzdwJKG2osJYjVDr8c
QqpMc355y+4jcHk85p4MdHVczKM+RDgoDwtBgZtajQnbfKFnLSOanwmNySDJCM6HEarRTSOIi+7i
r82dCs6wC0RF1xce2pti5iGbGd9T+O879bTCI4Zzequu7sO0wtwBSjZYR54xvbJRf4/7m2/mFKK8
Zv/oAp5k8fFSsEKHEftUU79lP2tl8uell3rw6/avcPaNgu84U4nLWfO/YsfRhbLlr/HZ1MhJ3YBD
pj/shzXwCyxWhelQ/U2uJHyDBREH4tSkZ3tHGlZCkKzTFb7dgkQDDcjmc3RjuBfM1Ci4Z7oQKBf6
YoJ6j1HkMlIgHD8NY6ghQLRzBvq0j8Lh8U/6GuZb1m+oF3NMQyPDdIaw6lecN0VMfaZI1Tji45xA
6pq3jCcEctkIjT6rAAyqDrnvVwDxIZtfiLf64B8oYIGLqhlwSnNHLWAaSgRNjwhD3MR0E2LLrOId
69FJRjRCP/mV8rUNbtfpTN1qfHTYqf2DHx3/xLbTA8moH4tGOk0zhBCRVKUBXvFdIDU5nIEPYqKo
D3dpGRVbnMMmSrqu34Nk+rumo7yAesHEK0/EVfcxVWT5nUjcWANgKzilXta+fBeUg/me7gQZpCIR
3O9hsjqhW/b/4GnRbMcdx02CgA5eI5TW5mexKsoFeFBpfjKrTEeIXdrUnU/tHJ1GqOZ4ZH5Xd8Wf
fxVOBulM5aPIfuOsXfgjJ+rc8C+yepprSROHdVIjsvxFw/ixHtyAFYKatipxWnLqFOdQKlRIlOrA
JNGBOoN5odHwaoAqXqclz2NwGGYB0zfHrCLCCZhXbyJdWkvKt1OAeolVCHDtBD7b3B1WX5/15SDP
MpWXzWMk99c4hRPd3A+0NmOtXuelxvrSASwKF+R+p4cHTFtBQxJpAwdOFNrP+Mk5o7q2gWuwTGuw
6o12R/fEszSQmnxZVZ+KbYuNFOuTWdtKc4TjDhZ/NxtWa3/SW/wHU17FBfZxrCRkgo4VpW+y9PMW
tqAHd1NLwvmOFaoKe4ck8YgO9Lj50EMVbfUsKM87y3sYtt/Y+IzfV0O0Avts2jfaSPWpWlw296qZ
eCT6n7inX6eGtZ3jO8D6uCx5vO85K+oGfmXjqu3rlz3BALgGoC0LW3KC64RU4HS34YW+okIt4CJ9
PsybjBldUQcWzYplEEvJKpPj6g6ENvWWJ0W86Btq/ymdmJ4ih1BBJ9OgUwrbNe5+OAdB7c9RaAoV
ECy4vWubVhLq5dwL7ADgVc1TFHB8sh4j3M+jTxOGUadc5ylMkz++GO750lUk2TD45G0CTwQfvgG/
ezjHLYn7/S0+IcRNVXTk6PcNK1PSmORqwrjB/pkS1UpJxn628bf8d5p5Kw32RSlRy//DBF+czgjv
1er9vBqVH4kVFyxKCyzO5shzLtwfObmos9S/xNrOnPA3UrKaSI1bhvCDdnjmSCOEcLKhjvrED2DD
3kIQf2IU5SX9qiKnEZrmoXk1LmqYnlu3jpSVlO58p1BM+sm97AZuuOaPoHN7BJ2G8ox1eTtJP1BQ
mUpwkdnsqkk7NocBkAy48ZFq0zNPsYsCuBFmwUyhsAeViN+Z7j/GdRTUDgRz2fNUd+B2HI0qi0cL
3d0NQn75vqiUegk4p0MJWEuHp34doW1GLSW8UY+Mg5auh4PRHLClVvFjQTzHfl6NzpuDfdVl/yPE
8ZO4lTezO11fQ3tsJ38N9W73VDBtpzchki/fwrPYbvgz3MAWp35wkMt5CoYlJOI18AerqPpGRY8Q
zwzNZn9hrNj2Wr9y28veMLyCfkIIxV5Wp3gHmUP3QH8AQuvzw8Wa9WmczN1Nwv0AAKEFmnKtgWNB
TDYGvwhTNkpcO59VsvwAVddWIQXyeuw+rPD5l5HzHJfhNa2y+GS7ssI5wB0UAfHS617LDimkQdep
yqQn8XMJNYoAQLKqLNkMxQyd3lLJUtS3gwqvYKxnxk/Cfp3rBDaX8VDugx73lMZvehNNlEV/t84z
Xa+ySFa9bQNIMez09OFtxpbenYS0Vn/FQ3HUKCrpk54rO3XmCpG5lmmPBBa7KRm0KyUlygYSdPvT
KRoU7BmGox9ozicBciFWSFh/sR+mmzY8f8r67dmr2dC2f4EphTBOdskxDuto6gQAMxzkLN/7z1b1
oIPJicGhPSpCan0TwV3uwJhGzqgcTZC6L+jERpvOAMBsgkKqGMabKIuFV5qfT+Yvo7TadWQvEJh4
GtYxMHqFkg+rPm2o5rT6PWxlbUrzGskM3Q+Wlyn/FY/HKhTr4Jj4nlebJN4QlZyI7S5QGDsl4PSa
r0Vb0b4kQoGWLk7ci9GT+YX2mB6cJHTlwGOlGxWc25KNW1U1XMLDJNnlJmNEOxD3efjz1IaKlB2k
VHgirvwdxm8wDjYeF+VQpL0bQ4nMOU057iVotjIy/9wNTMuPDJHIrLGR8PHlNu6Fptm0mhg06u/j
A5TBGuoYUL3YVYabSdJSbGhyV1Fq9a87Ym6cCFlQ6/sng7USM4hp7cIEb8BpFryDWzb9Rp5uRBeX
7KJlNxMLNGOcQJTHHbCe0aWGKde2eXbYxD8EvWgNJ0UNjS5Oqq7bhAVZfrc++nQW5LPXRi+bmHvr
R9xNZCcIsZFmGyYUGjys9HnEL9t1uOnrSvm++qnG5h8A1aBB0rbPDLJxQ51zDLGNmLFUcQzq1lkH
zTwZ/htTizNXWGJV+ArlW7GhoZMQxXDh/Stf8+OWn5GmjR6IZ3jNP1nc3hTREeAwcPezmbFGkVDx
pbyhGT29Bp2OFxbKP6FFMOdRuW1HbRaT9FQuJWMWNs6doOrMaSvVkkAydlpxTexKDjqpGn3K2u5p
5QgYU5gtipQpFgA8JYJKI4x7xS71Vqa1qVfevdBICWC6RJjJbsUqcbaZTXbBvjgC4IgJHSXUGJcG
xV8YTqTcsb4i29r7ob/8pnKdqtHLsZdqKR06Wkk8jzD/PeD6agLA/APbuU1+OxptoR+VgZvEJNyM
pZW0g6Y74tRpLt8aMBQmrJwFxBeeTiHLE0qKjVGml47b9Y5eFnYPzy4uBXFpRB/DxL4cqSshyTiI
0VA6Fdv83jWIjHS96rBO+1LvXk6PDHvedY8vuKMdN0WgCiDD3JtqSbUMpj5XXyNu/J2FnR48u/OT
AMf79xHPXRjG2I0BpTP29CEwGyaDJw2gPEJoY3ybUusYDRC26isjZSVXgakIYs01ypCMBKos00ib
zCD5RhDzuQKi1tB72FWLNbXqh3sOlIxW+4vayorJl/F9SJzBCBcL/pLgQXJhg9gkCB3/eF5U9Abu
82ObH+/+ToDaQGajNVJ1jXvvREdCs6YhJW9gSvN0o7TBIQw4xBXQu6XgRFJShtewg/WLyGWEindx
3aitNoOwLnf9+lVZ1qG9ScaDYHr6g8TTsGbBDUKn7pXgRb3Qr8vktcY/KeHXuIShBxXFE5ekGwc5
dccKmQrQ3o1yPeIIfiHEotuFqSsiDT+GGhS88SCOl5LXnPMm6s7zSwrszKthDmq3VaYv6YmcORdc
HPg4QDYi21X4GtBSkqhHe1SruIXaPL40mCPInGVr16V8wJesUFbk5XqbVz23JBfYTbRcSiRq6Hvb
APmIGrG7pvBLMBKMD0x1KoPYJG0Ul88igKzchbxs+XzpynxEWBCzA3LFDXPMB/Wm7Ru65QT3CF4t
mIsiPfVW6CSwThtqseMVLMytbeLcYroL6S0n7cUGdY4i/z237UBeUl32NFBqkDiVXsE+lPt9mOBx
zh1/QYDIXHdKVdJ0tOg2j13TB30DWrjsE05G33sRayVr1EC8b8cDUSWhuN6YR3VCNZ9VXMeT5/z9
U/Mhxm1wBh7zR2hNEEn+XfR1qn5YozrkOwZMWl5pqWSkgdSw4tT7xagKM5KfOQNWBAbsf/i0oknG
MlqaOlzJPIq1uS22++UkRaLjrjQQSh9heG29IuVuDynEnZ9VFMd4b8s3uPUNA5y81pAc1vjuQSCt
aj8NneKj2ao4bnl1Zj6K+AGNtfquypSGvwOiJbBBvS/NkaUtVhR5XPrPYkmA4BlFW7gyURxbZyQ6
ba5g5hZr3o7vi90ev4wUegnsFUq2o60zQHq/RZSriTHOe3zfdPXbDNSI/cpbixrhE+TfpCAMAsQ7
RYs5HOUeE0fcz6/yrnIPAM8+OgCQYE2TiF/7vERlXHWSptMa2+Rpi2wVEHnPo16woESQcvUj7CwJ
SBV2qd83s3EgtbUKSmx5CIC1MRyrVRx4iQZZzT4j/zy+4wlSy0PixmENXK3V07D8CDMIhHVUKDyD
oTx1qLLSOsELReNJTjeSNoHEK6xS50BjdmlSsMQdhzptz4xc/KNk7FILQGyCyiY2Jl+eX7utIBqt
6uzXdn8tToW/SNpFcsXstGhw2Mln/rkqKaqnDZEXJUuum0VXsESwKGCXJsxGiYI1IdXixLbUGUP9
OX9La2MZzrGxWroJRXS5lXIkGI+qlN1PZfk9X9ojGd0bYem0Mv0IDU6tsc5G6JBjabHOtDIl3RI+
6BRjq7S4xHcWOi1n4hfnECwRAWkRukDiy0NRSMCah7vSzYH5fml1mF2aP6120dR70XqYu7fodRsQ
4RmW8u+9yiBTFZtGyc9mFv/jTR3bCDCLfa3qTR0XVFehQkSEBjqgoJ0rnaeC/a5ZOkZ2ad6p9yKZ
t+mIoC85XS3HWzqKkZT+RYj1CvMR3QirSTV3X0E6jVNS0lL2+kNnqYsWASIn0XIKVu0hc/fU3fKs
+bK+LjYwUCOR7dU5rpa77WoBiqZJk/WMfablZ4YYAsrr6RjmdoMc2nJkSJUE4EFH3oLqTDFhN2V6
8uHm3rXYQm5VQvQNvsRs0XwBOH0yhNuSHVpQlmBwThpawcPgI5Dmuec4MgXtq7GKUZfYXOE9TrdP
X6JG9D0jZN0IlbwUl2P9cBh5vqEHtH+r56RtoC15Jk8cSE6OSUbcappWN/MiJI7qfGLDXEoqXFIH
7+otWXVFhiN3lVopalI0gckeE0jWG5fvHO8rTs+fhLl5pyZC5QVY71IV6myX6inizsUwQ6J4owEm
uD081x66i0jtoKOwJAko2EuhHh269wxMRKZ5VbAyctLdz2mTWJayu6+4U4jBbFkV019WUJ3W0gqK
u4E/+bQRqusoiRPVVrkS2Eyo89XdGOxcSrilNKJWpZYxJmxu6NQPEIEMDazCIss2kg7ZcgzZsh/l
92s1hJyymx5uVP79vKcA8DTBJd4HfHjZVf5yI7SmlF/vqoJ/VczqYWFL2RIt5t4wD4jsYBvQFPol
s1nAiUVrUdMDzhjB4uBmHkUmQP+IvPAmnxP/AKCp6cgyfNUGaBp5MiRD8v+1uN08GcNS5a3CtKHi
hz8vddBxaQyVlupa5KZ1RSuPTMPLKJ/GyrKmHB9fv58B8SrOcqRdh7jHCrb0FmG1VuIeCvNjLOze
AaCDBmoW3S0tJsT4RtKhgvGirgpiVqVi3OE4cd7jemyDqUvjM+Mpj1Ky86w416iYdXqKTTL+QxHV
+KyucvTWVDr+6O1QNLE2DcGeREg8T36kjKBaxpAwWzTAAI3LDl+uhBpSmeU+Aq37WxLtsAGN4OVc
OEXkMAIt6m5AkLuIlUKdakjTaBLsz87lRgHu299lVhvB55GwDvy/vWFI2l9ZKnQDTfhA93aRfj4x
N5bi0bu6gFNVLEqLBvzCl9ED1xkEF+y3aylAY6n3hCfZDCF1dMTyMTt8yoPmtKfydaOmgr/+5TzA
CYU6e1nG9t3GusxOkGLwJmZn5GRtAd0WVU3iyKHxXbU61++edByPLXshlhf7JDoGWMP80w3u2pWQ
e48+7y9RmCD5j0dEGHCH+tS85j0+KxypH3lZarO+vCL4YPbE4RwjOTWfn+qVLIKN/9fwlI4KNSUv
FcDEXW40JMzYML6btIQPC8/RG1xlU+TKHfuJVgQ/cCnEHgIL9LMgORCKYuG6B3HclTniLUr6fMFz
n3CiS46Kazfbnb2t2gggCIdf/1aHaz+9iG3BcKN5XOBVJl35jXndQmDK8OjoD4CAQd7ZQV9sCC2g
byDoAGZlqH/K1fGDM3qRAPX9h1P3QvvxZj8Iwah5ZF50AM7MxzfqamgHjbECWPP0NSVyK97xePO6
WC1Pu7kkQBJMuvtmoyZH6zgeQ9pPLjKk/mKtmDheb1GE4fRb9/ODW2WWxUAtVTtH8WWvkBwWoGS7
YvPVtdugUev/Dgh6TxnMoaKwzxwTu1Oo5T1uBRubj1UxoqSM5yPloIhl+I88k3p9x2i5Ay+0IXLd
gQhvcSsAwAiCTysxbQfWO1wTzIan/WZKmwSYSoGQ57Zs5AAmmJLtjKVvPMaIvleylvXGFrfp42Bw
1p57d3rkTqL0U2Y6EL2bTfld160ZHfWeC05PK4iT4uGBfFA2LATyGFg/anvdQYZc55I0pDNEsn7N
6lJEWaF+TAo7v8ZXI824LsDirm4sUAIWfMt94m/RN80lE84SjI7jFdMxJslJwmzklV69GjUlAoTl
42PerdAQszBR6T0pDOsdw68s3pZQ6jL9bdELd0gb2RN7Zy9UPXH5xfGaHhL4AaJ6bztEcwXA7nXD
DwMZN6qvbwkdr3n84sGDCb5BrGXFP0glCvElG9DaOgYROlvPcgyAMdSiqkKiQuUMnSd2fmVL4bFI
P4SYP9Dyzy3OglFeC6a6t8ZzZyoej6X6n5zVixU9FLPBlUC7Uy9AdnFGS65rrs1iCzEXQMN6LgK7
4CvKqRcMZArEu8iUXGPYOu6i7aK8faGJLVrnfHkqruR/jnlGlG0Mmx/bBgBAU2NUWnRHgh/13k46
hvgK4bL8uuyWX+bqawlO+8k+cWJjFm362uqVJKI08iC3jezkeUS48G5PNmGES8BUdgFcSUue5veR
J0/x5clAVtaAr7D2ebwUhwCh1bXTVZSY/5eKdzypaq8UugALzXUqj681SXUpMlHSorfx7Rdd05DR
caACFYhBRJRQV/91qOnr9kFiFaDXIcwpJ7BGqordy01CExuOjmCsy2H810+FMtXLWUuu3M3HgUhN
RUHcheT0vLkwlQVGO8LsDsTh/CNiGtJfPB9G//3Hr062RQahOzTqhFO9Q17KEdmnNpfzV86vYIeN
luwuAvh92TjiIcQaLHT0iiaWqFGvBlIRxdMFGVEetJFSt38Lxd36SV2sJKSN/CE021bK70CGflcA
7Yv54hwurPRCrKeWvCWDgNw3/AwWYQfl7J2oXRDKXvVVnwLTXEF8aZTrcCwCArR+Kb6Bjd04W4aO
14mZMzpensFWLO9eSMjoUEE9QTVyqVeeKfEUAKoVjCB08KqYrWP/3TkqaTxVI2K14fFannwZx0XR
9bun0Iwk+KG0Quoqw1YP5by3AgusbHEOgkCeI0mOZ4mZAhR1plltv6/Q+8fzWDIrm15k/mk++krw
eLWoPfFM0j/RFPqS56R49qB7nNYdBSxkiNl0XqEn+uRA1Clpitn41n54mqZ+buh4JpVa63Gy8TdF
dzyacF7LkkYANQaSfXfgb5257dMpttUmanwPQvE2Lotx4fhm7Pv+vqMlJf4qJMjb2QA/xJlkFgiY
XBYXA0/ZOcenwF8y9+FFVGqmemRx1Q0AdJVfR9cnlBNHfbGJU2WwSbCysQXCroeR1utBtmUNuBDP
xRpZXr6UTvXRFTVMZMCN2S8QsC8sHt15U5JbBmT5H9J27+cdMugBy9VqUsNHaYJ+5owe+epgnohf
5jXMpre4qrJ+lTB/kd8Jpdxl9MxH3ch/gKeZv4ErS5OE+hccI7UKj0m3bkS8iOxDrI3mpYGtTJOs
bjqSN9hcytoFyslpOvmoN+xQ5HU8UbyxN4dnnH/AuIQtmzWYLIB/Bj+uwp0h/mQsWzZ5tWx0ZITs
RTMMATJiY8UZ3KciIftBqrfC5tIrvdsjwZBbWsPCG9rBuAL5008/Qm/x9bpbgSkJKyAdMBHdCadM
wRhMw9Ja3V9Cq3q84WGVzcAFRyVgxeBiGDeeuFnkgdTenKMTKf8zadtJhD0xrhKKiRwz+smrSQcZ
HRs+urAKkpANztQNmOu8evPTmIQTme5taBXAESIN6b7F2N1K47slXEe1dYu/Wa1xfj4ZnaXeRGau
zvlKLdVHI8ctYTcn8RT+xXCTxfgYsON2opO/6wCvpn7gNhWNwEYl+cvVej2SAbYO1MyrwIsE8NgM
kGGHoaKNikWzt1WidvbAMT6xaJz1yTnQq2QJcchoTwnPh9op+hgjVvEdZqWOHr3AObl9ItsGDewa
aCPoG9xOvpMRlqDDTxHclGwbWCNhknJQB8ADWVcWVl6Td2mGEfLx3U3/MbGP5mtsX7VmUJ80hWf4
cbwnn8PO8JWm2kXtNUS1rL9KxZVTIgJHoIk5NIb01z8STvAzw3oqQqyk4BfCMg7lIeNcXNAAD9XV
3Tp3Sg9ZbXzfTJSYggbdPrxZtHBpsPvvZsi10C6/Zq4S2Uf4xw9yEm+/ytlUOMO8I7U8ffmb9gsR
ujDo6ry4lFBSsO3dn7YOyBb2AN9gUh4lo0mrMsTP6YLClbsLiDKJjVm9MsIBEbQcj3BsuGw/kCu5
dvlarNTOIHbbBA81N6SM/jA5535/knvWppTVu/KU4I7HzqF6M4dDQJc9YrC5bD9e1KXJ565+32O8
yEdJ4gbohcO+ql91Z6ro+taXk6IpHVrmeqTnIaQyQy234MAeGYsBOU+0cYtjxeOEPvs2uii88Uwp
34/Q5RT7emJ9zvPf+zxN+qrNVzf2yhd+6NjZLVBNap1OuYdV9mQBfI3cPk2xyBgC/Bv+Y9fiawUO
7vfpr38JEueE786x1oP+FgfeykWZ7mUTo4/alcGmDCy2bQ2wH38W/X7Yz5VC/e6mRP1WFN6QGAMC
TDIh158ElXH/0+jIjtuMQW4mzDRTj0YOG2Ci5PoLENAa2FNYq4cE0scpuIIfc77Y0mueipCcrlZp
wucma3qgBSqBZCVCryE5ukEmJbay8h+ZLVhrZ23ThvUgckPDJhG0T8sYAPpQ7Omk+DHleQ0pxewx
aCg1SDHrkMZHCugRYoM31DrWZcotMIObUt8BMivh+lP73KnPYPqAprbaYlE4nVGRf0bbYXjPHwBK
V4kUNrFm8dot48dXag0muJcw1QAyQr5jpU+hqoH1rs1m2GGhHWuWdwYt5qfVJP8JLhaHb93Ns+Bz
TBMkk9pk2QABcxdz97icWLqa1zXWvN5TO8nW/TCKR5RaqXlw7e/cKEwLwLr0AvzQmflPmVCdBmSo
WGv7C1EyLC6UxCgB9rhOnofx6HeOBoMfkWNBiamyGxNdL/MAGItfsm06cHVOkov4rfO3TBdO9tMg
XcoAgT+evNYLo4Qukr6EUzv00Ym5KY4TgDc6KtirrxGp12Z44oUJMZ9kSXQcwBdXdzP5vLBKVQYt
Z26xtGqD8eh0x+RZxus8yoUzKCoOYmJGRr1c3fDMw2iuIxaJQk5kcG1gq24NwTBPiz18G+7QpetI
fx87DP5unJV9PKOYcqh+HW9wxNjHuI/tHGYVuZSB26n8Z/EvI6QV4qJOkremVkNevqAnFpNl59Pj
cql/ojbY8jIe4fkYX4nk9A10tgP2NbDrrIBBpv5BaM840WUDQdMNjvITMkpb1kNCT3e5HSnv1GYi
npoKCYrTwsHmdOR11+MC0wOp4SXjec2CYd7QJEHwPX1rEMxNFV0AV6H7U1289I6jYovN7rAbVbYP
z84fq9p/Z+RNZmi7Yx7Y8hzk+UjMDHZMA6esNz3g+0M79EymLfl8SeyU+m6yOFyeWQI9bH5SYC2q
W7lcGO5EFksSqQJPP6wcbeKyQrL7VmC5ZyZoWsxNXRPtpAL7r8psVSC9Z5uqvtP6+ny+Ce/f277d
VESF5CzRzcL/h75OX61jQDkfpGdnJ0kApB0EfHl4SQBMyfPfwOu6+w+1loUjPrvS/A1AMxIpRT0E
9nWaDSNJH7YCrB41KF3fnEI/1F7UbBmjVetFJPh8N9YK3I+JRzqd2leENTMyIJSaw89FlWVps49p
oMAK44IMfeSV7R9dGU23ThoLUdMUD72vGHqFdNdcU3bUbK8gWtLyQZeuOtAWYminUubiNeD/pIWt
xAMXPgPUWEb6Emlm+0iy0KQ5ZcJeK463yx83J5uypeN1v5fitNPqmdNc/CacFsvwN1Hzu0ELxH9z
FxTml5RkRAv5vNd24YSsdS2zV4lvcHNZkUF+hV7NCQIPUAir7yM43nso2MyUgwFCBulvXkc71Oo2
3EjW/agS3sUi1uPKIwl050C9Iy2yBc3uI8E407PhRT5p6lwAkXEHC2ECuIYoutSHcItMyUBdWItS
w86wshpXkpi3W81fquJi0qwmKE4cz+nhoJyAYx/VuqPskHWcVvYyi6ZcZRGG9znVxA85lZrs44Vg
8KJfp1ZO8KANTOKrtJFigAhBy0ol9JN5+KitWrDT1NhZ3lwHXjzGIIfiEED40Wedt4zpANBlmK2e
8jcI2iFgJw9k0oFIBdWlmbg9PXu6SuuG+soLYb3zBuHDc5IgUqRi0C8Qsz4GE58WjiM3ACr28sJB
xekxoocIdRISvVQnO3wppKr/Ws9BXszBHTPmmArlkrS1XI48vhrRDEIHqMb13bV/yYxY1ol/D59q
uolGEVJzwrsUuSMlICxfe8WduygArbGbNDqBivz/Yo2UJQ9Fw3jDH2ULK8hWGw0PDxIZ60zvAgVr
CoCmRBxF0qQIC7qRuCU8S0bwDKph85hAdNgfhQfWCythMliwYxHzGWqh4cAw4ibGvgNSiZIFtNoT
UTJVdA53KPRBJChfSs8YiUCyiTWLHLP832HLokGO1/3HPcA65U3GhdkTxXDlNg2P+IDY5C/JT1h/
/P5g/Ufr5bHmSF/tqmZMlP5ffB7IiYWl70QMD5hhz2iw0KycyeLid623XEWStCRNd+eEUsr70OGh
Musqg3zwbZB3rh6qb62+cdyRsOYkFwU21fojH1jdwhVP/9EStYno1W4X01wVMe+hRppnPvd6Nr8H
rOKGJgFfgua0y7t4PVG3u8nO0YxLlJFkhzy2XhiZd0oYwx87/hl+/2Nqgf6QtTnPuSuZkU4Liemx
h5bL45xJYXIt+xmj7TkXpS4Yeg1i/AaaKDOxmYImps0X7Bnr04aYxn7tkAlmR7/GS4X1jxFdFVeA
2/i7zJv5P6p1W1Yb9NeOr0V2HFLIMOg3nTUkURL5Jk/ItnNeOwITqOKl2Xvl5lJqOE2wFrHs5l9m
DbEtaeM+w5CoRvGqtVpglc1zQ855dWwNv/rJu6lIzVu0wRlUNrkrYk5yR2sn/q9f/1xJW0Gaiqjm
pBXAli6OPrr4Rht8qXaKKz6QJ6wW3pZU/PSpsZnri+EbTgzd2beHoNFw/vfRhZcG5uPsrPNVfHNl
q+gV8d2VBWpI3rF00SU4eiWLyIXs/rEp9tEDWpUMuw5uE6+EdWjxEGceg1QYHemxyRhEd01174YN
K1FRH2dqQIrEnQxR7nBH098XNUOO5xY/1+a+EIx/JwbH+aW7MFqKpVcE3otpozBgdH7q+HHgjl6h
eWzEzr00UQADxdOKwEiIsc09XC+iATQ4HQF1fhyNAa0ZBBSO1EjuZgm8P5bSa7tvYbd2qIoCPbS1
L9VtCtvUoGSIbvR3fpwidEIomILKc5nInY9Q8emY2BLs0eLiKVnHX7Crrb5JX0b+NAG33QfNO15F
X4y9cvpVx9D7L38oxQvcALzd0Ex0ciuJ6xZwYWD2263Ju8P8+DazY910cIyg0V10ucy2wGAy6aKl
Qfvj1KXkRZebu4gqvOQ700+bzQFNEY7RcpZQPcoGBhbjx6TbQaFWIRciioBNEq3EuXteP7XqxNkY
PmIdu0AbMzbu7XojVvr6RmtX07QqCaMgwihqMOjI7AAMH9uyFpDsUcFR9o5HB8UnRL239hiCBcAM
1Um+hxK/apoiGPYe/HZ0qBOtjMComyBYP6JKu0awhiW/jdxRB08sIAbNca6kwdC7gCdpcqwde1/R
oMIhcieBtrN5rsnC560WDPQ+jAvJqSWWxCR+m7W/qP40VahHL+hqF2qNAvKF8JFNmWg17CgtYK9k
8h1CZ40ImJTgwVR24c8+ubN/N8Peh8Ey7ji7WLsPVt1kIHk9ceerWKsPFuy5il8CNAeGQvl7vuj/
8TsC2lxt4ijbNw9PvJTIuJPGwk230/7mzw+76MhX/Nhv7LJZt6gHdhTxCNYFjtP7hUU61LMNyB+8
lc+CZYmTDLqfsA8VM8RxOw74cHwAYVLUhph55QzQ2U64faBwNl1U2okmzHGUpO07K0o3V352L97T
Zra6FeWLkZXHaQh8fdfBNTa0MVJn9Vt+qUw//qsTreagzR1F8bntuYGqwbgOdKuPqN0MM+aqu6XR
vpuDXaQADxjPJ45vH/aV2yrNnNlg4ljViH1YBB6L2eoopvv6IHM/Ie6Rh4lIrdLIjtDZuydv0j7U
isUomdOgFVkayh/rHesMh7L5Y2xVRNP6hHHedHnsrYbgF3KAbcJjAjLJ5dNkPFUhdg5ZadurEBdc
VnBCH6TO3vxIgaZ9oM4Pk8DkeANum9N3JRjfC4xeEBL++uw4ydyRQpazctnvjhy4wcHIbYyVqXCd
iu5lMcdX0pzW5aBACrfnOGkEwDrf6wKR8U9ZxXzgygQPo13fFKsihU4v3Uoef7Evw/Juc4Uem+kB
WuzTyi6645rlky7Jpkj3hSTPgHX2br2ahnfQM0t0ORoVNmzLwKN82idgE/trlKVvvUsFdLofpevH
i18p5bwTmTkNJM+Q4wgYyNPasmmqqr0gAc5BLur8D03dFiammvrhXFG+2jm8bh+H2u+bmA34uU5T
4zS9dhlF3dWf3NM0GLVcu3nPkBi2Nk4rTlEiTco5NDFPB5BmuznA9EzG9M20XwRYOMwEVX/iTgtH
HxELjesqlW79SWLJf3DWm5/JdfbbdOvb00IsKjySkLmqr43j7YoCvAYvVE5KpKoUr+nSS6WMWTYd
4Ld5F6hG6iBNNe/H+o3/eOHmE0D48Ycz4392LmI25lz9DyVjMvT43KzCsKoQBchqOrhj7v/pRfqo
f0fNpZoJFGZX4rzyjquYy2Sa/6OVn/O4mGts/BGYn9xlfrCBqr6tp1z0LQnQ3U5zmdriEjj5HI6s
g02Gn+CakZl5NQ5bDDus32eTbu6EnUzQ1ooEqwI3Vot4OUCbYkpEV8JWsE3gsI96dhzjDdP/c//E
lmgEJK/9roJD6BG83dd/w1pF41Zt8oY3wivioED4WSge2sepARrKVy/LLe4uoudqKV/w/I4r47PH
oNfMnuSqbrkrR8vPi0vLG25mTUtsaKkMwsvo2TSZLZ5V4JR4/CVW1SocAk0DoW1ZBiSTySSLtQsU
71xahnA0ecN2sc+0kN/cIJ31KLf4jrk2z0CJxUEabudB4bdiYKEC33DhmTajcuf5Ha+xrwvPqkTU
YTNTFdLPq/pFZvLJEyS2dAOWAOsm9fzHc0l6ITIG6awRxcgvn6PafP5k3I/hpwK0VRIlvoCVh6xj
2IA84U1urDNMAyt4HWwTqFqCnYbQMtJWJOiZYigGLRsarb/izAyoJRrWym0LJEIDOcukTh6OypBc
v8BoaH5uwEjFd6QbVSSIHGJrmsEC0EIUBpbnjyuAmcnBcaFgxyABi90X133qoxb558MiJ3qFrm1Y
z1+91hQDKTt2DmdpU0+3iq/bJwMUFK4D8fLLP34Vobbte9kq8cgH2mVGsjLMefXf+Miesr7SSn8p
E+4JNRqyN7HWCWlWFzJLETN6/2uZxEc68nJlQg9cpZNUZgD0cmZczv7cVn8ZV/rVS/FrA16AxMh/
s0e3/4fTwc9fXVYFSaKUQtXAU4scXtWD1alPEmXZiQ8W6haoxZXF579JJj5mZHdn3kU51j7E8/8O
8mCztKk2Utao2Vw3Bo8mqQnxUZ14Jbb6sVyvoS+o0XuPGeQ9ssbq9rVZWUATBf4i1dJvIYLqnYHo
ZFv5HT4UvSeO8ouT/Ds7cGUj/BNkU845AX0+LbaXujXJElAb1dpbRGXRZgZ9MryyNxmdt+tRDNT+
FQahPWi6QMapSozrdR8B1uYWDMYqosIEuaxf8/SPeRWANBqkQPWiE95s6HDw9+IF3IBb0wb5Y0vB
rhOx7fsijWAavRUPO3bsZZY++VMHIrxiq2HpBpwwuKqRWWQNuoZhsqzc3QnCbG7YTiBLlaOoRMTF
8oNYu5RsLVaIjcmEicbgXbGjSyn6oWR8EAoNzCHCQgBbrFr5H4C2/mK1s925+iRn0xKldH+M3B58
7z7Zmuz/u2kOTibrTi1dyiufAgRBfYXzlHoqFw2P8n3mLZ+vmRJ+BBHaKAHj+vRO8r2aAVYpy99T
5KM11+xe2pyKeYwrOCJj90l9qDWfdIqCjuJJ8k+/KXRjSW45YKVWrGdFFwQwzPcf5Nu2Wvs0SnhE
FpIa0BkhET6RPdvWZcQQd9eIc7A/qrCvnEECjCXKQfLNobCaQ3cUg1pQO2V6/hhaJEIhesyAhdbq
rWdN4fCcw2eQ2nTp5Ht3WxddRf/gIAIwqSnMqadqYUoxRl2AaBHwKMdj6oJI1TvIHJaD+o3Kklxq
fpKZshv6dfWAxrcX9ZAqkQ29j0h4wuMSpoq5mIm+JRDgNPKYMYe0sFryY6pIeyxg4R5s+0jRRN+Y
ei/F2brS5QgCUQm/pok28ZGlrGTiXkXXfLvHmW/vsok8JQtyzSy+9NVC2WbDaeukRERzvtbBFbh6
j6yBpPQ8CAGRE0k9WlZG7Mmqhy6ilMJ7rLUS90lPknNDZ0oD99CyT6IGElKJwK+Sp4N79Oq9jbDX
cje8SLHJCqI/Bf7wEGnDnXiFNH0YH7cHIG+i9L6tLwokTtMCBVvFGO8/QZNLi6hHZpOJFaytjmZN
OHOhIEos7qe9Hcsf2a3Xy0p16st4cyXJz2rMNQvJeXf8zw2yP7EPQIl6rCdbPf0WIizdhUOACvrD
wJCZOxKcDToiga6UuKMEBUKkGjin3plJ6FCnFO3X7tC49d5I0aAQlZNFDP22hawJ7KfL7/D1X8Gb
HXENJEBZa067GuM7Ppjp7ttFj/MYmYE0LXV+zeGAkrwQ9ti+vo1QvnBnWLlonmkxdE2JvBqBRXYz
bM5FZ0Xma77Txd8G5pkXJNBqUObRmnEWYgQgu7cG4oasWJH10NiaNco6iF2LWPJaqQ/LK+6en+QB
HzI3D1ajWAS+ZPhw+Zsj+TE/puHdfWrgiANKbL94fJ7dbMqqqEaTtKesE8u9aAzhDqHjVOjN0chF
UW+5E3OjjEkLQiUYnmjFznPClkgn7JcsGSQJYGwujoX/6Jq9MXVuvbHGeHbhA2bUo0O7TrPt2j1w
OLmBpCV7K+l6A07RGQ+7tfMlE1vcC6fmZYdg59bnMgIuonw6QlKNyKqSKTfB5qkWt6EwJawWWGav
bcMpOWbO2RUUqxtTG3cH0vm5TiVAHczxOl14iyREFCK/gF/6zf2nQL0oWyb4SmDwrPleQ3F6ikSZ
SQchL6bkSEt2fFkKHpBfLDWxTwey8d0hC7Vblt0PAzVlP/BqPVXTYBb/pZYCzYW3ibIgSbEQdHXo
8z7NDpKtA/ffJqJUDjoAGicvXGzvkB1WKa7jaivYZ6RD1GNitUQY+amOjSa/eKk19XCpo//Ucf+X
sCq/lxqeVjkglHQVy2pBDYhfsITGKorPhsF/d8J1a28A4NceaI0ju7OP7C0CJmNbvpOg93ucvPUQ
8F4haAoyLVRKwPHknZmuadwpEZDf5oJez9fSFyJ/IzTC0dOc6q5/K7gjSBnUOhKqeKB+4buu/bja
aXMDaqrX5BX1DVfcvdfr8YAk5tafiX3bzmoyFY+DilrjWg72smMNBfj+2Af+8pnMSK5RTQhTBXnl
Nh0fTFX1hsY7tLXTNK7yT2kfofKQEuEQklG2OjmotSdhO79ZAwdzQTVLzJSWmB7WG0kagcCWJ7Q1
aQJW+AMTz4WyMu/Z1tZGnBlgBC1ZdxhiMSR2zV/pfFYlnqV3YLwiWqh13NMDTJG5HS1qFlhIFUrg
K0rFY/0S2eu1cgilxuIWXFhd8HhVjNlBMfOnC5K+CB/l18A9k++2QAWVG6O/qfAQoD5wTNdShEKK
8OuLbQqoUHSr7p/EgIzMJyILQ9HtahMi8peF1azilHV5sjIqKukn+hRKXop4oIZRaEuZdY8lZ1i8
/EXlbrxHUzMRQ+GcgqeNVyyT8YBy1ane21yf789vm39Vp+Xv7PiBrlvPxrgNZihAcCYFIxUV75Xu
jmXFV9Df6KwNB8I/V/7B1zcGt1ekUM1aXTe55VBCz01dqrBh3JnSRYbByDDvCURy7tNhaa5Rzr3w
F+2iy4FnE2BpSjuwXVGJX2FwdQwL0uCp3G+9iB5pGdmqpqSIoez1aU/vHZJcRYc6X/WhyembU2Sd
Jzex3tUvHqYb6u4YYPzoGbyf5vqajFokvBjg0Wrw+oHGSsKnEGmthwGkEi9+BwHRtHvKguN9t+qL
XnF++GBrMiAmqEEEo0zcsaRjmkbZbHWr2VuHUX7P9pcwF9gZIJIuALYJED/cpxqkYCWEss7Et6Io
6RqlxkFNsUUsLZYubzAFZMuzccY95hD9GFuuEelHcG+mV9n8pqK+Y1e3Bn0CK68Q/dBp5UDi22Wq
cKfKTzrRVXPeeZSVKAI/Z4PDp0Deq0d60zQ82AJPDbjTP28v6JDhyP3ws/sXd6MYWOyZNsJBSkWx
LpB8kIU4ZmNC9bNah3T8/UV870gyPHODPWFtgsw4SSSW1+QhFxeQJb6XGv93y3ytjqDeZE3D845P
wL8dDsZSZYGRqag4FLqANPZv6BZLgB+6Uv6HPDo6n0X913tAdhwiJkipqEEr+jZ+RlvjkX5zldWv
zNIIH/dvnSTusiFa3Bx1cWH3nsKTcUdXpnvGiHPl+z9HeU+Xrd/2bfpayVT0H4nWZZaMC06+CGsD
OHbaWY+0WOa2AWzFbLYfVuVA5KyvTw4dKIWz4tJjlCEgY27h1soxY+nxLsFkIUzKds2vpGCYWrBK
2z5U4fTDHp52app3jWePkFZL42V215ypIddtQpQHlmc18UaYcLBs2TDOk0TAEqHcVKIYX/BPy+wK
lD3drLNgOJ/NhZEbMAmL/CG/u6etLAyoC4dgCRdkWp3vAnJq7Bsyd69l4FXfvr/7d+4WkFsUHIa1
PO3MyzPo2h5oqbl92U8yYTSY2x4F+/eelNwaJ6Oci7QbMoGTVjhGquFaLXJWqWInOl0kUH79xR6X
Aq3vf+xIDCFGlZSh13dEbqxVb8gehSjmnztrSM/YlX+xY5CV/VCaSe1VQHEOzpxKPJLjEAw3Um2G
hfrjgFYSLLJEx25jUKc3/T47/Y2U1lfAcUoVbnNyj1w+6fPWStAAd4eYUZNz0uCqv57QYfj6lI4n
QplyjIS5JNm3zRevqdSRjFb+nFrk0e8/ZIQe85JDQPYCEQc65yIa2IUQDNHILp/Iai+D15VPq/TS
6bXFtUIBj/gyMHnTYf7pdRKLqtDCOxKD521KyddnYl4qGH+INrzGBrFvjyM0RT3r8Fb2LWsHHzJQ
LrBNpNQJgTz+u77SxxBREchGOGmxAspTSYhfkc0vucrp26gMyBhBWLAbRFO1GCCSCaS59NG+HioC
tKVTdZ8BZxuqK7fUBetKYN50zUxpOzNnQPFrymaPa/EuvPuQ/pwnCM6orhalOZl+S8CWcSWGWBzz
EeiivdPkRNe+NLTLyddNLIVPeXA4IcDGiPUfpCOFvTNEG9Ayqg4QS6WRHU+oBRZKAT7gUUr9SRdP
L2vomsnfzsik8G2fdX4iLyOfMumIkqODy/9F7TpaRBVb1z8cWLC5hyI2ttLlREFfbjxu1cuO8eNY
LlpVaPStNWIRa9CXomJBjSf96nkB0YGXuvIfJqxtj9MvXzIeL4rpeoFc2NBE+GQe/IGZwrifpY1u
R/MI6kg8tztdcy+Oxo8p3aDT6qc1I4Zv0VJGCf0RB5WPkgjJeP0XgVMIjQ4ozBXmO7Jqu4ki6Kmh
qSYyzOvc8blegHB6DbRMPg3ilH/ELzlHxFDjqh29b4I7HjSWRc7t48xm4Om3PB9AbhODYJVF3qM1
h3uvTetY2sWVKa6vBJtTm8vNPxZLj40JkBJ00LZ7U6OdwMX6JAgba4I0LjCsKRRNNaEeCfbrz4om
kUSQYwtQZ9zFazSSKUmW2ImmYIwVbWBeQDj/8uvRNy5jv0yj0+lnXvErTLTF3rX4gDtZdHgFfNOL
txbacFZlPQMKsHQCaB/6HxeZXsivv4b6RcEqKhQOZspAqIaydgUMUdixUoixtP+m2FzP4dDCwbqV
yqKGhqJ7X6BexjPHla1Nl8iuaocRE+aulj6RBCmx44AqeaQ58fw6DNU33Wedw/JBkjQohmoH3i60
xIsLCOS32+/FOi30EH1ky1NYLQM7JhnIfitr8LyMaIOkprQANgcbzPfy8OfJL10DCg1dIZVO83C5
OCW0EaIV3ssoTFNtuZk7VJc+3CGaQhzVTvFCnDdpwITBa5r1e7m7isH1jEF4B/zJnJVbGhtX7gys
ucR3WHvi6y0EtmyiaedhcQ6R1Rvft0ITtARXCiLGhkegX/M/OoEORk0dewRqCaEyZZ4MkCcY8Lg+
Gg6ldKU/8qSOvFrle3ALm1Kjs2gIM108c+bB5Q278mUw48DzOusqSQtCx9WE/voIKuzBePkaigA2
im6kWTVij2jy/+J4SqFp7iLN3n1pJBj1uJpXwx4N91dPLyu38o4GsrETwewKWbxzgM8zjG7/0g91
EOkixIkYvIbNUJ3JQEK4zK6cApCFFL/zbdbES4+CqDodNrNi542no4uzDVehNBtqSAKB+RFnMvq8
u66z3JT3GTA9eMwMQpsp+CuVAadzb87Ny62eK9vv3V+Xtle/IQ5B7McD0b+e8bnG3iKtDkczMO5h
3rvnP7aiL6u41CHPlqfpKOPdJVnlOFDrkH9D0DagKuTOMdPGpL4sHFEiPKM870rBee8A2kBh4uAE
bh5DiGa6xWFV5OzlK81m/ozPQIQLxPKus3JlFkmGWy+jMPFgnQNlPOHhZ5fSIccvV/31ll5bKTFb
DSrjs3BU698BqpGsQxbC5eYQq+ZFZIdasUX0Wu1OiwBoLwR977mxcMktecPCMO3DGLwMTWyKrXgE
flD3n1BbwG5751QblxVdtzXkBI3zm+b2lUjWQj7lthIdkx3KLj8kSPaGZmAUcs3zPT1+rDKPnG1+
hEKM/OWZ8iHHrwO7tE0p9qLzlN9gTepySISIA3YlVpNaTkPt+W3GajA8ZAZ50XyiXvgaC2MJpenY
Q187GB84WyTI4XtX7d/yWN3KQcAFWPe2KjDFmvCf9aDEKebYf+adsnAK3nMfzy671rSorPEjoqlb
vf85JmXB+0kZiHEuiS0l6NFs8aP2reQwAF12lqUKA0Y+SPSUQCgekHRZe7+hYqCLiXw8hHH8x4A7
fP0cb8u8zP9kqQvMtnoc4KAD0884DVgaD947gchAlAwLuzKA1HiANxpvYx6xt0YPTx+urGNZJWU0
yCSxsyhiy52SDPzXJvqDnPd7ydKigsKyDePq+EjXgHS2kwTmm2rgOPLnVSsqFRcq5nQ9qzu8OB/z
2R1HAP+cz4wMgvoDYhUCH+n0o/Yde7xoZ41U6tBE9C9ZO4LyjrinL8FxORSOipWFQpqtqH6w3vBe
lkT8boLs9/OBFQszG3zo5O26g1FmIYHhWX+5A+Jym6TnhQW+b9R9zbDrXl2KCkYmJB3fY7XP3eIq
LaAucVDaMjF9M9VdWdIAr9JUoN6XoYpZdWvXppxCi60cka+LF64RbsbXLDIfUINdZfYyu6nnbgDO
d6ZxuWxaNvAu+IPSbWONZqwc6cTFhHHwdEsdih8FN5FXQvh1QW9rZUCjb9AE0TGuBSQsRITlBSxb
zU5EpueMrovYoOBY2KEfGO/Tfex2pt+YrvYO1xfd3u+N3ZL8daKzqZ1VOAcvrRAEqcKgeRkD4jX9
29VAEVt+vyhb5eenuMFUYqQtHcwebNaXKyQqPa8qI78Jm1febKpF211XQwWcSh9JwJMcmisPQpyp
X1YH2yypqzddrpN4aBAQvmKyR+4Nepqq636pA7XjMixZImHM6phIM1Qk+y6xbAnaiJnhFWG8tzVI
uNoPejm7/6mTDlCTYrNUX7cgVe0+VzdNBd5OXO0pzIbLvLJypkX3OE/c1v/O8VzTky7Fvhy/rNPM
uTlT8TdqQX1aiDoenWIymk0kTSdbvk+56P9Te/W3QllFG4ikG9ha9EGp5HnR/NSYaGC2QhAweHa+
KNPRwG/zMzVyF7qvtr2nYf8CquupQYZT/MAle63lSFJuJ9y9dhH3ILMyCQrGfF3PJruSWXt7Y6Tc
7+VNbWyYch5SotkXreQ9+VRadM51zcjOFP/ozqYRQD3DwV3lagsbmHZkff6EYO6DuybIZN/QUp2Q
ZsU0Vdx7nxATjnDU9AdlQiPy4p/vY0TDm7FneRbiia9xC+fh9G8/slwCkuNGrAs4XUWZ0QWOCBh2
AgHnWi1hKewcbWCvEqPEIOqUbKAM3cFVd+nKnT5RVx+dYRWuw4INAMwEbH3vBbqAHEztl3HwMbKK
VQFyd6WYOBKbQTdQdVog9j0YMSINydXPFjIx0yD0dsewB2hah5sejjafXPEt2lJTpW0cJVtE6ZUn
P+qxyDSzCKjYAnb4qJastG5cyVclPIjuVQysucyl2LPdbp/1oTMNRZDP6tgNHck5qxg+j10WVgU/
f0m2nPJ4q/9Y2D1yYSNphGk2N1fvrQMF6NoJE+LqGtc8+ncggYjSfZXzUP56ca2lIJOiXb+H+pQo
xqrmkX7pXye67LY3ILQNC1udFN+8bnen8pC5hxoDtVbQdi4CMSBDmwfUmqCbssE7b2LGE0/XCJ+k
9Nk1h1fjmy8FgitSIAGVK/QZ39U1VSrUo2QQwULs6+v+Q8E/r8oEhaAfDcSCfP0HeX+3ypKeCaEp
NAAIQpz0Jr/z42w1dIpZKmqDyX2jz/Imh60pvsdeIpC6VEu5IVRO5ukyrVCyv31QqFIcU5xbzmH0
0U//GiQxVepUu2n5iu2Hdb1zL5+6mJFkUF3HfkkjCa11xQHS6CBijblWqStT79ODsocJVF3+9+FO
wRtCQ8WqnLZfntYMcQ1qC0JwOodLGo4hHflvpjGOGvLdh7qmnZ5VNCr1X8J7MGopF0DGSROtNiMM
OCWGPf4ggC1D6Jvwd0e1iQceIgOaN3zNLpDAVBkBxrjJlp5kb4pHHzaGZVYCIfimSsZxcxLj6Puk
O237hgqBmO1R4vD2P2aG6J0i5JEhPEpbBM2RTDIin+HiqnYQQNbVS3PBIA+LF26X09qRDB15HAMF
5XSOsqZxVWyF5LBHuUKPXzs5T5WxLB0ooTF07nUhmGts/P9a8unaW1T4hMAflP4IK2u4EXzquV5I
xr+k4Bb5w3qHej31PJ01bkLrpAVvA/cXuJM6WeUp68zypwDX+UrIyewYMYExuC5SAO+p5SduxONz
FAJq7bxqmNlFkXq+2Ga0jUg6YassFFqoe4DorQMfNyu2dJN8lgwVAGtoNin6KPiEgS7PQXbmm/I5
1mJlwlzzsUnGcBjEPqCerU59ru/juztgM5ecYFtoOSbKL44NmkyXUVzJNb9GL8e7Ig2zsdOWksbo
B2KcVdDjYCdTBdNdZz+rd1qTT3/lpBUShvJiMlluxYUC2ii5oCbWRUf+JIhzxyfzQ4pKU1Bs2reD
jQ7zXpSn46QiWygRZgfUAaOwbGcNd8SO4wVMJHE3ncenw/Qn42bgACnKXmbk8pqhVBYX5zcxOd1h
2ixpXw3/gtRubMrwYnEfxXpD2j0fWmKdSOzC2BFQrLns12or9u0NJolBqBNReyEdiK1IpsgL0VDP
W2OU8aF7Gst3fRoJvFdZMXHd1WVeM0Bk4j8p2pseySICj9zbTfW/2MKxJZeYB9bUS9Eu8BYP3Ccs
ltwIfsrUzShKvcBzfmh+BhfstHZtmJorj/dZ7xDWxYFSSjClyvyk+IWSQ89sH2efNuKM1QB4ttse
jmt+1lZ4S3ouRgcXbaFm0R/NZFKntWhImcIYJf4mvfGvFFC5hSxyWXVsDWf+ylZaScPQJmXJn4fE
vS0Da4psBHUnH0K9c6hKYMsGAMkNMngEpsbVWM9U9iTzB6Es9rYbNWtMNe//axh9vw+XMaLKFVXI
niiwd26RkMBTRSiYKeZlGA8xdPAUpr1L9SbNRgZtESQaJbvOrhyu3s01KsUoK0S8vJ4lHIubwRD1
VaQCxsShGqYQ+o9/m/VwVYbP6WBZG9MK2LJ6X4DFdWU2spNNnugf2zLp8z0UL6bh3NIXg5oxa+n0
yR7WNnfaQJ/D/QM59QLJj1CHFYfIbfRt9Ccgcy40yRu0DF7+r/3oFNPkn1mBcO4yuj210PYtEGK8
OMpDTRvMi6IZQDHHB2yy5C6KwgRstxLX1hFYokjXHdMcTV7UU9AzXaPTpP3smE+U0/QHX1ZGgD5X
1gcWoBE7+7C1cWJpr6IX3A2UjCiV758HPLckDnDDWiH3rpcjKr1A4YOxa+/icbA4WASJKKyMXnDw
5yal+dKLNybUbJW/IMp7lRmCm60gWBUkbMlTWbq0QcpChL3MNmD4JOT7FraEc8uG+BqfSXi6DGs0
t5vfhRKQko6d27fpxLX1+t0qLnkPl0Zy81i6ZYV/kGCKH9B+Q53b5J8uXj5fDiakJUpLUFmEgUVR
oprOYwyp/kK+uXXR0o8KEZsJrpHxkN9eaBIPrJPBbg/aK95f5Gmyw5SDXXUZ2FLc8E2a8XIASELg
0/QFgXNpZVN+AyThbVVGcPpQzNhr87VMAYsDfIXZs1rDlyc6iO1TOKccJpZXh/+w01xxSiH+k07A
n6sq8V05YImcAit1CiFf7LaPtIHcakjh/vOpZEDQfN5FTrWgRnJvDncnytgv1wvMMqZkJxtqkwtR
vazuqihVZp37NW6KxIhBYHc72EFHt0DPF1PcxeTdIv3vUk8wHd8xV2HyJKr2nA/RRwnjcCCW/BhF
VcPQiBaKI1mcaN2uSdly4mHgvNZ9mXlFv4vBzNnzMeing2uL6sWkkyU9uFgEdsKxKL9O8/SXQZsa
jr4POoE1iyjBY+fMFjHzAsLLpz4WjsOK+sqMX17Q08gARY7ayyvG9OZe6W0B8hyutEYIVh8NrqNL
0Idbx/mro2TsWQRSDwth8KpqPH7hhddjImEqfPtGnuCPSRiWKtlINK7k8nZQPxc5cueOMJ1ZCiEm
cKp0B9DGI+9RBpsjPSMHYEj2cBg9onJftgrAbuvg+Z0vHx8diqHxyWTr7qvhPB4TMpEQfdqPNLw0
hXKLvjie3hYYL3D2grugkIk5II+h8k18MGQalt1r9jrIcQGNc1QZdfQwac4Tfgb3jIN3wnbDBgfR
onPodjudtqSkyzfQRx2PumGQ+Nu1cnf+YxbFbFSInWyJjkTNTJyKwyeMSddJVXZUoeUS+j9mdD6K
vGfcFNyhoKxNYc1ZM5JbV7pnbZLN1Y8xoO0PFpAhl1zzr0zpyzVSlkl9tMVvTOopWubCONwlFy65
aILe3KunpnaAk8bGaplLHRP/mDY8oTHOvwNVgCZYsae9vH3pRKIYEMiAFTv0HbbMHdyd2KRSeDXU
QszQYGSEAhoh8lTgh+LNWGYRcKA2mQIMWBKlBBrgLBcjHczvS26RX/FSljej4vDnvN9rMKpJg4v4
mxy2ouNE8MuLVYAngeLw3wH2B90awJ/IOtZsfN5r5eR3zDPDL+ivSNT3+X4ZNj7DsR5uLCHTw2zB
bkXA5kz6JxZP8GF8wNxNz58zZmeJcJKu3rPmrNgQ574qIwaL374FWMyR1eYGKLym9tUY6d5kkpKp
qmiHaJDCTU2sWaB3C/uZknOdXJPGDBjpc9F60k9nq3YH4ehH8NXi5pypc+/KQbaGaN+1NMqXNAE8
3Q4+LtkVTSXGiqqetkrDLZJBqa7GrJ1pH/ixEAmYGGit6a4JJEmkO7sjnOHbXn25yM+gDBOQ4iKi
HbIiNW+PFu/ckjkf5n08o50IDBTax7vA/G5ABu6PBZGUMEsKHoSwZSmXM7QwSZcaGPG7yxq/kcIQ
igzbPTH1Ng2swXiTyDksNBFNwK5onrBu308Ly3UXuITrlInn+TX+mSHE3UPYfhwd/PtQPYrYugFP
Ka7w1Cyjx6zU78sL/3Jz6gWB4dc8bdfwYkK0c2uz3VsljV25Ts5KMhnm+Mj/4HtL01Rk3UZ/AB6N
+bzAXhMZqsfSO41dy5iJQb431ZH6NwmG/hc+Tr0ybbSvA7VZxaWnBuYqrGMc3JihaiiSA2SNhyBr
ju5AJU3y/7mHkER2LO6P03krGxBAfiJJefcggHvSBpUBr8N/a1UC3bFuvRtnGY17dO0+8K4umExc
2l0jAh5h69nbH4TS2h6dIGmEF4kIRkTLni6Mbwplwz/kfexyumnHGu1zmhrJeKlMdGbvISLi0BtQ
dQJZXr8YBh/gZb4FQ6ZgBbydrU+VZ7hS492Po2WXZj1oFXQYQ93j66ePXc7lNN9+Y70DNlPkLHbX
zcpDtI65V2VWqfSKqX832LrHFn3oyNKCHUiMTlvNHarA8+Jdjx0HNnJWUU3rGjJyiPSBqX1GbSXT
CNlThm24F+EXZCjU5sZeO+YdsmGS1PLBjj0L0u3lRQa54A3kxjfh3VOOKmKJlfKhnSAzyqgSxO9l
wqZQCQMEsHk7Jom4yG06In3pJwj/ZRVPmiSiup0EoIE2fexr4f5cUiMUU5FrdiaUrk7sqTQfdS/2
f6rMIoKKZFsiEuKa/zo6b2rUR76EBG+KX5OVbYQE0+p+8ikY82cn5LXOT3LCB/ioS0jewMG4mLiA
YeXdkuWuzL9hsppxTGdjLCaaj8EoWrWtVM046FzPI1MpvZEHoX97enn0+BkMB/ARa99nuQuv6jZx
jbu9I7/p3C7djuToiS/K1PSkL5I3zKcsq2Figm+aMMgjldT+rlECgKZVG4EyhUZb2PhbzJFo2BRC
7MU0ASfhS4Qm7xz25xkBhCxef334+PrTeRUH1U+nB/Xn5tRvDZjz1bwajAmaefIoZeO/7Fy1+GKP
nM3ObtDBFJWr2PLyZAvXRnZjO9m/Cn0yENLmCY3suKQNfRqHkvnznGaWVPpAhEUBNEMmGBTv4TT/
04oyIXJiANZgQndIprCLEoqSjz+Ula+YYPscDm3Ws/sgmsVPp2oUPCGgcJ65Ko8ctRWQR/VbnJOT
tb0cU+eCL2lFAHJnOEl3hlbQCFJwgtqm2xVLW9Gt44xER1XyywCHJi+bhCBnqY3o8u8MU3gQ9fec
Iz7D624Knu1rS46IWpBU2fmMJ7UPMHyiND2QWoIGE6u9xOBi2NQC13RO6CE3z873ylvFns5wbCvY
5v50l3OoKyLUa1QgNEhvHsvblA8NlsPGby112O4Q40YR5WZujuHYO/Bv0LZVee1I9s5S59MIg6Zh
tMQmD+HU8QAXuGusARUXq1fjCYwyIiHMcwR8hDKjHv4OmAkfYRNhpGRJPpzfy8b+431jzD1u9k1u
gS/Bj73H3Q5koq4ThuGb/b0xRHVf3bRALS4SZYXkXpBMDnwnXocKfghP5BVZrHOFPTUbJ4pzJ9sL
JnvdnlQY9X/jPFB5Q4y4gAD2fLjcTK3vKOhHf92haLFvl7K1tTQQeUN+jy1mgFebRM9pK1T7KfIV
7VodgE73drVEoqA3eBHF3gMpsLqfz6TSLL9dSFfSvAieLylfsSnZlf/f+Mw8uzZZhL1rUcRNhvRJ
XLP8OmxkP9wDSvBkuemD6YAI9+hjeywUmH8kQ/esCqF3RikAWfgH29x1tEjoLWe6BAxhiwbie/RG
Cmk+ysK1kejrfuof7vadKx9Dzfhddn1dGX8tBesxIow/9wof5rdfE0c09Jx/fHm0n7sGqYocZe4p
uDJNVZfBvAqo06N0ADRYMEn5KkkgEE24OWQoptlsLPazpnKJpZvPm3CNsCyUm2EVzoAF/1wKks0V
V/t/+uZTGWASYsHLVmgabHg0T8USHY2chRDCQzhDeyFu5IIX5Xt6xQr328ToV7GUWA0yl0xzPB2T
bi1DuEnyDQCbyk3w/v2XB8PER1GDaYSKj4Mh62pTEC6cZRQ43A7xzhn/xmOVq9MfjqeZKZpUOS0I
V0jyXB9tlkyDNMpoikvRVOnN1gNALuRTp/eIU3pKBDQsExEsPSCufoFOUiM5krz1YQqYWi7DHpP3
f12f0MdsFmHbxOGjSKL/XmESvkJoSHJ2jI46xlmqx1gToq6OSaHoZyeNsBMmvG2F5RyBmhuCVBZT
RjoCUggsw1nX6p44foCb6CPLllqfgu+GSntVKe4+02FoaDD+kzxsdI4zXXLXscE+2yov7056UXd8
wA+tNJpG0iw/yuDwI9OkuAwWm0kmZnBzfbw2MnWOWVibmXvVcGpdbRoW7Cg/MTIsQnmNdoRFQyhG
Oln0s4oR5cDmtFRCbKU9aJl8G+nb8uyMpXNUi0nhj5+wlTjz1BolVn51p1pZybiAOxon7rDzd/RH
tQNuQcTTLMk2IqoCWYvcPdCrRKeNF9tSy4DN16+ZB+SOokBH3OMWr1tz4i6f6ekd4kFPy8h5Z9Bd
mEUeh1f33eDTfqh9DHzkhQzjqlT7bW0QdRP0g4y900lwvtgVvudtabsCfrR9pq3SGhEmoVnGOG9E
O4dm+axxZ4A3+gV0XHvefAcjXzkOTA3jnOfUcYDusoh+ZL56lOXJNp29ScIqyup5GMchSIYCqJ2K
WmmoEcbXABmcz/VklPPMxbYBBA77uA8BiFMxh9Yx/ZSuRhZe8Tr/83Sdz5LxCuFVMO+R3agSasvX
T6p2K/l+suTWaQf0gCztnd4FMMZPv5v5vaYGGjW2kkVnwwK6FmKgLcxB+N8De/So3dnFCZekbpZ5
WjDOFpdhE50iSLU+SEJTlSoP+2wZc9E6k2+0mef4LzbqlLlkuFOhyUx85xwKf4I7wYVPGShEefSQ
OFNhwR5IQ7tz5GDUGFB84ngym2YyTmB8hOEQWLeKLbNl9/TZrX+HYown9WyBB0T3y6VZmtdEOBIF
mvCl4pqheNeSug8JmZ/ym4T6HFIvqjz9LgxbBFnIM4yI+vnjvF7HCqfOBLo6weOuR4kIJYzzPwuO
h6HtgyzQ5L6yH3shZMfgfeha8fhbNZedXStis6fr7P5X3HopwfYLHzlFXiKiHLI9MCCEdUqwxjkK
fPMel0bMzM0OrOy2+1uQgV+DDH2aoWWpBOotb6wp3qJTTkgm7cS+xb+BN/Dm/GxgXa0T12tDK/ln
JCy8cRPSpl8BTOEkXgx+LQXaWSZQSRxuNS1z7FJt0/ndzvSjZjaq3rFVIXYuQcJcT14EPJRP2TwO
3MWJ80f6ntAkKAWoGUNvpYFByvtA+IFzYzOnWkyACQD8qHhi3rb3U+bE1QJSmIEI8siDmbsFg2Zw
UVblpKBHLBWfrDOQ4hJMbeJUCpR1kiRhM/iwVk8He6a5Sr8nearA9bkjDtSFMmVrGlqndT2vrawM
2ET5JIhj9t4wE3Lx/xWSRX+W77dfyRJibqSvplnSTJrsa5jE6NMaMpq7F5AFoAeW+Piztl4hFDwH
NbkXDaen5sq2UgTwNlEYEsmiLxycUZ/HyqKjqw81V3r4sCCQm3EaPDMHNVOuRuBeoQyQIDpPkcT6
RPt5ZX7nc9M/p/HcjkTM6//DW+7dvWRVQrkIPsFC7EHhDLUrdPl+eOPj5Is0e5gPSc/b7BYlbl0W
Iyqbv/3d0X2PLJ5zv6cKoksTnvNkam3MSRWaluY9oZ+pbkBk1hmZYlKTrKx3lVeEIyTP9MKAM14C
KSwFQvViQ030rDodz+aiNaa4WA//TbQMH4tYRoXt9025wagkWxTkySahGh8/7JpuLW0I6smB8T2d
YRUz7nNnlVFmgjoyJ7mVy1egEHDSe30azW10Ahax1uTImOjB84wYuGzlz555TeL4uShGGfKtuG8N
Loulqhc4SJtpUa8vA/+9xNFJmWETyf89fjIoBTYfxhFCg5jnfBEduomd0pjglhrkRFqwHaiWcgWi
eYZX31FOXDUYQEPHL7stsnsH3TMKLLGgmB/hvKRKxKOzookXhwBLWeaqnx1QIdF0J6ujVzK3w7md
vntFT+76jan0lVCDvNGL6c9gxefyWTb6U2QNIsGO0XLACvor42ouQFxa6B08YLcXZACr+IzJWCOa
UuAAFymoe+i8XhEOK+XfxES7yVM9SuLCz21DEfh6Azqtxcyw5S7s1zxqY0eRI6D8yy7VW9k1YJI3
fJSmQrvpQz4vieHYEP4siZa8f1lqHVDFQHW+jxIFjLi/VvvK4qGgnqloOHVSi8Y+NdCn8bwptSXx
ikTe5y7ui10rZLEWKh6nIMAGcAeZloEVBxvw2wVtKZsvXxVXU5q4uqh0k0U8r0gHQKY0hyxJT9Hl
BhRAkzmdgXOEqwn2pcRnqKGYpCQ1ud9pDl8KMRYN6gyCa6qNLHYZuK5Jz5CtV87r4pZHqTGO3c6G
CLDsXIuYkZKXYSd8hxV0fIsARoKFhBSfTaw3xmqvdGSSfJNOe9tuRzdSRprMS9E8BkUFmyZK7I6c
VpmMeUZImHqvmGPj9dgZttzCIQN7LoOBRM33fywUi9/O+j2Hd8msyOPGQDVAGmMRmS2eOqgFN29r
VjBmMLOIh4tVd6XXOF+P7hKJEjKEmADsMLKyqGjKWU0tnpsn5ot76xr5yPCDQeSfdVuNurWWvl1A
n2uM0GRU4Ge6Zzfbcoos/Y6Ve7p1iln+TEOSXww6OyqI997M0vlpgHQP6BbuChppMKlfkdcQG/5F
W/0H1rux8a6devrDAlApDLrSVT/xwPJfyew20y5DuvR9dhCKFMqgooog1Yc7JkuX5pAuzeon7HYO
unywLB6fU4twMu0YFak7fL0MJGyyhtZYSdoUWUHkeKCr29t3H7FxqkH0iZm/pzDjir48a2eTTSvI
eCS55uf7YYrQVQsqx90OAWZdfvuXoX/jTnfnmxW/bDwrBxIqC0XJSkrfKbLmvxEDrSNhRG5xnV6V
OpMUPxNft7Z/6kTYAn1ufi9I1h9zaJOGUw99gbM+0QFDz8INDs7zDBv8efY3Stua/AYBl/+tkMRI
zFp8zkBOAloeKqQUl9+Yyx4a63gU2VSIgd/hggJsHkzNmbjwfY1OfyA+NATFwHsx75uw6NtTRGM6
ARiyAfgpYhtBmqdZnb2sWCBR47l6VcFvlfuzwv/LpEs8xu0bLvh389+tHSzvLZhrD8ppC7yB3dMa
/W0s3Y/EA8rbN17sbeVZj5XLcCZSoujKfe3xCfl/glhtzxpVtzHC+cJq+nrBAMv21znWfciZ9S4V
fe6tckC8KlhWA9S/nD+r/cx8nMMbZYOi861g6ifiQY3r3gRNH1D4fPO+kw/SDxOqP/CjurUu4EFv
sIHBBd27LvMYiig67oUjdPyJgH1OCgW6OjiGpioDX4Vb+1QmF21FBP5vKLrzvpmlOGxYCjv+/Fu/
n4zbiazPttQx+SPR+b7yx3uUgf0pkSNONGwPxljJ6luIn0gN0Hxt/HG++u9+GZEWH1g8Drslo4B2
Hs8ndT+Cs9o/ZS7/qFzzN7gTn2LYjBU/FNeg/Cj2cvNoH5EP9E37iKdpAn4ENujVphViOfKM7NUw
lTrj3Das/xTXEfV9smfaDXeOQ7IcqlQl0TuZwqm3rV6zqQvawfkmwQbVRbf6uhqGKKisHR9DMFpK
8Xht2HPePHjGuu8OFJp80bCzwBNVfQ9T3bvF33PmOfU2MOFaOZPa6dxd7ZdZXoTj+luMXjKKano9
ejHU6weQI2fW4/1FKrd+NIxwe2wHw/lRFD8aZmKNKlPTFK/qY06GVF1iFRaXOiHjBfWeIoVBY/i5
NdfFKtmeD5NMDCaOWfbQ1BSq1Sc/0Y+lHqp3/fuqhWsoconIsLT8l7UQ2GmzEZXxRFGixQfMCg8L
TB+2ZB+88iwvZ3CDDTeFrs6gczgypLMfQILPOMKi2fQ8x/8V4Gz+2rh68oyGu6EBZ7kGmFocs22W
bajGc2iQfn1IjtWTykCU9sl2kZyPScp1blL6g344CRTRNHJpFDMcSfephF5olssfeOkez5FZ5FT6
4PH4hEmEiTfV2KkOOWoGweQqNd8kXkD6jVgyDnGaZ2MMZKYxYyiiTMzlI/PkiR7OZPEVPhSz7OLB
Hlr95zsdeJEhTqgs5J6UfKPUj4YoeQkIGk4AF+AAkIXMnGSCeHlDOKJ1NO2r30cEb6UjR9sFHAQw
hR3op5vR90XivHuqaRvL5rfhLFuVHP0zBxbxA9PTaQmOlcpK9rJOaDrgRgHFzsLo2KtO1uma8FVE
gbYndL3ezCva/A7/ciDbQzyZIPfhwY2fiOSnlivmRHoRAVHgVyL2EEpLzKbqqPveteQJ4GY+urRS
lWCWxigvxNbgsy2icD6PtjF93nQigJSCkGJQZMBa34gs8Rwkh19MLAj4mEWSofu+W0nEiRw2DBLy
Pj649ebPkBvwINqOPndaORoi+TcgayZfiaK/HNaILdjHcDXMTugat/yv3ME6BUpSW8eNbaCWb74H
w6o0pld443Zri0EGu6pub/cG8YO7dXuuu51iHJ8C4u3GbqOr5/KzcyIfDh0RHN9vBRvsix+7nhiR
NRg+30z8MwAajbXlzP7jYDuHFaoM8s/7cScZXx4KOWvwVtcRZxzwX2wJWdGBqIsf1u51t1f55VnQ
y2pQazVgc5fJaAoXo6fgw+/g6PjzKYkTFMF40uGfYBT1LIGNRPikBAXMhDBvVLY1Ii35JaO2eVBY
NqJOQn3Wmq9P/hBMCFebSxHNNrbYKHyUbtIUt/qLTY99hWmgCWaO+tMKb/VkQ5LWywWKPbzofOtu
WTLwcvOwcydmCScx6sn8hBTbW61/aGQAGzzKRzuV5GOAZsA5CwGyethEnAIe+Np2HsxMTMKyLMXS
SJE9SnpPxsImyBZ5R/D4Jyu2PkiFhSlOUtZ4livZW0d7wX2pM2eNJdd+2UW5QpavROTNBApPFP2t
YNhqT+LRdJievPvIkS0myysgkx6CB603ZeY2UzpZD5Oo1FHwJ0TEBzJad1UOuBW9DQKV8ms6Hkag
Ig4pER/dYJqAXLkV8bNukzpb8mSg0M+Z7b+r75adyPfj0ZjFPlgn7cpAlLGFIYx8ht6iizcVKuoW
UUhvJYkhHE+YtSIec//TVhRL2vhnxfRRE4lCA9N6CV1yusAGBGQ4nnfFVuyJMnxiUevmNJ9zgBjC
cqBU6G5rQYm8zPttQZI9TPljRLogKcgb8eczdUDi5irkHINUh8QFbBYcK1WAXYML9/E0dSB8JDRM
Ml2sJ33tjr/t1U1aoKUSt3ih1Ap/CR41KT5ukru9720HVL+7dVLw7OsXwwxrU/uywSCGyKNRTT0e
fVUP7XQ5NXsOQx1lWrF13dXrYixhiFuIWTmQBM2oNafDwO5RIfZ3UZJnAqycD9OVrodQAV/cgECn
fRs9S9geUGYSvYtQybAm53on87/3anOkoylvHDBmzdfd1cbo8QAzHP8l0pactjYx9ss13b9NuDbf
Y/+MyefxY147etP4Ltxl5ukePlRPYFLap977JH4tezmQRmmgTjQDUnXtu1TAYJLubOXFZSbiidUv
0b/vZp/13mggY3ngsrgJafc3Bp2brmSVWd1rk7GktiSOhy8VUJbDbc88Wsh1D9jLPZ+FuCsKe8Ay
L4jX0rkyzEAAqdlfvRHPZzC7yvAZnZVcKwz9fSHNDdnjWIUKXJZweL1waS+NDCJiRcgEkraMRegv
xkfu8h4vbR/A2Nkdoo8S/a7hMbgVnSqzgYnBndDHkOv5d4rOKNl9iHWlI406GKvV9994KKM8LxMZ
Ymf/tJzUl1pzRvw6WRWEd7AAx6JpydApYcMRfvYTQG4JoKUday/QtcJfGZbssd6fjh9gD9S/lyHr
qrVEzsGdhcfRb2XbrewSnCQCWQcgQ5ey/zVtZlsEHEkqCnqFBHqZDA0DtPz3sJgYcmdr0RdJ8KEQ
ihypn5OhErpVFzYTfIPhJIkTM+Co3QRUsDuiS0MBhxlF8fxEJrhBXvhlCBu1CB9buDgUWve6yfuk
x9i7VDmslUlBfh57aFjRrBF2aPz1y1S41kCaVl9N0r8RU6LtAB0vo+ihbBEaxDQvwogQo4XbpxRj
s/yr2yMsUQkpsFiGmIhCTOSHcLvkVFJSslf3nO8upqkaSWWCsYQ7jz1s2hywkTaydwhZGrinMSoS
lzG0UANbQ3Yv3SAYe0Ep2ojYtxs8LlqKA4eb5l1dkEdtN7dMlnkcm1mYYJ5EZ5imYMai0avM52VV
Ei5StFp8lir9wLzZ5wfChwRw9h9tdqiJIud4xQNfdmbaM18GfBeyepUPioCWEG+61I5q19uU+yqi
huj+4NO0OuH9oc1W2tYnNmcKoqjGRadkcttjtHHYOgskZGaJOFH0/0ei0aIFtRJv8+rynWSLcfJW
0f7HqMjWrq7XX6p5x6lj1d3tjj57JHiKWsWsBH4P/QwE6FlkcVYD7KNh/EBMF97gnpKVH3lE3J/N
nnhCe5MLWTpS3fM0W/qKDON9+IFhX15QNBN6velh2uwAr9J/rtpsG0mUt+FrDqWrlBInZrFyeBXb
/VCA92eoHqXm19Eo3h1ODsHgoeqYHPijlHWRV9j23og5juHKW4/QncjT5vX3eH15yHq13wvQLKIM
WPX7UXSzlitFGlTFgJedFZatHv8m9E6tewPwns0biBSDk8h25X6CnglksnKtVryEdZaapolI8BJ3
FFY4SA51rLpy6Kv2scrTGilg7b0TZNpLEMEFjl2idtN6MxB6i+LHeNZ3pYbPAT68jCsrDaYKijCi
rUkygG1zxmkkCcI4J1tukDZcIevIOpKRnAue04XHTHrmz/9bQL4pmKY8kJwmiEDjgN9kWkYQPIPU
NGaYqfod8gNA53xGkdPhH+04zoIfF92bgorrv6AQh2mjXc1qKS+7r70q1HrS2jzWADOvQ+gcnTKo
IxEYPhuzUP2mkUbQL7QoBsCIPFcmJIzTL+e9uC0PsocfmNonFqybr9oIjgNY3CX7t3coKe9H8kaO
6jhbz8ILs3BjBwSQKKAX7JDfVAr1Av1LVY76krCT7Wont1g+7zJI6cJPiCpxnYVLdj2osua6Cf77
7dN03qVC0sgt/RByC3UWCsPjb57R8xRFl2kHXZBdsQYYByqs0UumD0H9fhDgq91/quXv6kq0KzFb
HouETGkIbag5iRxTLihSiX09JUSn0VMje3Ki065CDRuDxOBEk3CpkyQwdpsE7BXqC4uwvhChy+ZE
WyqFZ5239SLN7yoHltSndeHpUhWF236uWMAJvW4SiExN2O/SGkMqQ0fHCwVuVru+sd+7CvVKXj+r
T7Pe6Y47TsYdx9hI94p21GFWlY/n1kiiAkd7bL/XvOn/iLFd9AlhxbxzKtLlqf+IZUItCVtAQkhz
3WrPlTM+SPyoUviMcczrP6e8PTmtJFiQWU3gYAuf2v7v0QRW0nXHjxF24/lr36V6fd1YjPcR0ia/
iU0/Ay/hGY/JDOZF98i/Gfqaymn1wKm4z6+PymzardWHhwkrPyLayjQdspAATWrN3LrZjIObREr+
twXMOWMvrGdQJqANjBqpMSL2JfkQFHMUnEOrpUr7KrTUrknyum3OJPAEem1Jyh/Fyq5JkDCtqjtr
lW0VZEpeBX59qfR5boLb7KAcjhcQadKfHm6aWavtKRmbKcLinPF4s7vDKRL5xkmqBDMy7ztxnc1W
clIN5w5H20J24qzQlYWSprLi4qUsYgBZeL66+vDCByggJ+IVHZVwS0EvgyOpHZZC0PxphXdTca1A
PbNVsP7+WK0wWh+Y4QFsgRqlIPd6I03gSwfJNV2lnDF2eihM3cIdwg0XOMRFxCxkiiobzhwi0kJy
z7gU6BL17eb/qMKjjD4lk5grTD5wLxAm6QycE8uKQlMxhXcCMkJ3dshq1LS4cV0EXv1cAm8MMymR
1R79oG4OIcwGLiydDj/bHKHGk/LbsW+vXuIFu2R9yhAVvSy9VAYndbYJAyxtGCpxO6mEhy7Xnev1
7/D29Zz/4IPA4T0k8A+wrPNiqx+oC8HtRnla4iIeVLayz/EsSjfsfc7iKnZpk7Azk04b3CXyQaJd
pagUq+cB/q5m+BRRjYWqJRciB3xIhxGIgF9iNzcnoAHJzrTlsV04mnHiXvQh2cCR5liyNExehGyQ
oDW6YrpyLIkv4BefT9ogcqRD20uO1l2EvIuWrwAglFtvRouzK3N3OzJfbbOqgWhBGWt5oBU+Hxwx
e611bBFCm/pl+7l1CpZG3SaJPaxHtdBelqEcWZQeZYKBpdMxgsCYW4WbolXPiVZhom1UfnW203Qw
OvS8/DVGPFMv96syvdEuwMBm0+LmPXGMgT55DsBBzWExzzCZv9V2C8+zCmvGRmU74SILVuMaMHsB
i1b7zW5szUCd86ZplqDonhzzvaHzVpwejzXalircvBZq8UE11X6OEDZpVs3N3+NnmUJoM4bFCV6Q
FFFJcAtcGdZbGCRyrzxtrYBg/B7IQAuBLpO6c87vbY44eE9Gof1Axe1Me1m5mAtk/kV5e72pLjfX
lcmmo26vAtp3rz9H7D8PkmwOH+YJyfTZGdgujHB7BwS8BQydEqyYfF3N8KJEr/IM2rHrCM2P0QZp
Y0OXGDixBFEHCAl4oSfqZqaxduFjiHnmB2j91bCdm78oQuDjtwH0calnPN8oHfHgVpEZljkXtpXe
Iy1sF0IGDbndjb0VHMiqabSNtq2iX/Eq/uwXziQTvnamtCubL1KQg4AcHJFxf+PEGg/pgW4eDHz/
K0D2pYUMMCn7LwQLnedLcHhVIM/g/T9cDy7xsBqEiCfosODR9Kw0DDVB+ImWrggj7qWIVBBSMchz
Nv+Qweg7DoTimoRoXX8RDLd+BTHR5naIKF+ZbzI1De8A8ZLBtm9b6G5w5p+kfn1buoG3gW2OqTSS
T4jA8wCEyExLeCva4DoV81Gs5UAx6Jp5xBbvMk12xGhF4/V+Q+9OLBY+JHN53U7Fv/eESu3LW6Qm
5m5BYCrVPRkqOuPmKdltdxWbWNeBNqeTniivRurJFFHrNe6B/FWl3Zv3T8SI4K8hljZDkSJF9Jz/
uQXGGJWD2JQyqw5qyDAuQX2Dfmsec0hbccJaUcfbtxGhCiri0NnINmF1UnPsDadzpqRx+5fCCKzG
iQ3pYeLWuSE4L8Mj/92k/42wq+gQHt4AJbfDHNu2D4Q1soQsv2gcmbLLq7SI749wtpCnjFQW2WuE
NJkL6x4+ZroXCKPmIyPt6DFH73R8Bz2T4593Dvx7PVUoq4j7QHgXVMsY62g9Mc5KEQbIX08Xb2pA
1LQjm0puJaZg0RNkQzLCS2bM5Vg/UmPreOLRr4HGklwtAlBn/3U2sk+1LCuwZclODLHqqdd5qw63
q2RBU7S+nULv85reYaQrNPoktirDfYqZ7eEUKbaPLqUfe2ns5iNQAQ//PAXMmj2Y5/LLKk97Fup7
7FkQ5dnfXDodbO3hHaCAny9vL1p4Wa91qhg5EsR8PscrHsUGjvpdnBfo9T0iH5Bc/cOiKymptJj/
0H1rO7+Wj8O6Kz3KAEW+XONSJ3yX0+7h5sksrKTBbKY+2uWFKzvBGCFpxdD2cJ3qc5QXcLrgvzsC
qgsAX8d0QjzBQ5BeKIDGgRdfT0sGBEGvmrG3tuuEm4jCQ5werfH859mPTljlSjsBSihiuOSETKII
uGAQHdyrlb3N8u/7TDQ9EDicVuE7yr9bXJw0jiMPSjRep02rnhAy4BqHsCZMtWPbxBUJ0rOkOao0
B9eurVrewWZZPkcYEp7AYzrFQFdtK5C2bs7Mm1Vug5UcNY2h6Pv6n5zRraFwSBdMyIIbttjdhCrA
tqHcq73fqP7FqTuQmsIV57CBphL/hTN8bSfjYVUfIhnrpVFO/fiUile/tdIFRBuvO9H/qdpk7DBv
skMNjS8XH47ucw6v92YAcJW+Wdz5Xki3Yrt6vHDYRTxzOqJdyJLgZzBcY2QfFqVYGrCUN41FN6Xv
Ex8oKtBrZPbrK8zeZ7G6nF6avdeJyxdEWDxpod1JdAAUOGeZI3TL2gfGOIHyzgV4wrTGpKjoOEEP
r5gaiZrppOhlzZE0JcATNKrdJ72sYIiC6kftTfZK4vEMNl7TVELkKjkMa5LZwIhh16dnl9a70wev
nIw5jLZIf6HtdQxP0mUe9FpphrVJjKZj6RiLChN0s2A5vA2SwvSN5rvwGrzrxsqEoJqKnwmt7dp+
wRY6xdVKzhVzPvNBCN4t7p3D1gUu2uGn7RrFboTcZ+o9NJGY2gYg3Ux8zUjaBZudBccsYBX4YGMF
zPdiwQcwn1LODxbU0NkI2ax6kcU0Idb/PzyfGqWH6NncC21TookIqmXZZSU+DI/yjDggJRJqeLV/
18Kxa9nuYAL4ahgKyFHVdz2zdDpAKeJ9bE+0CS7/Ta/KV/pBKTCvl/wXBgVBFOHNTjr/rxJ7LrCi
E5gZyjiPOJwM643tmOSSk4x5ZM3OqjQiwwLsHetjv4ddgkUzrYtpwsYL/Ls98Rx/Hy4MZPJa/DBL
laedpoooQek/8vEerWnsYsg9i2IZQN+XTqESCf4EGPz0ympUCQnxEkl5mkU4zvVzxTyNBj0258OO
TFy10tBB80PO8Q/dQgWtcEkIy2RIZdcs56LomLkhbpMXYs3bfbTy6m/W7uZPuomwyBDNu+qHxQXM
kDj8i09davBEoThDdxFuc/s9P/3GC9sK5KFzD7cwXtOAn9X+GgqR9YVKoEwt+DMDpYihkjwYVG7p
vxyEU+156+p7agrtdeFclafPxkzvMCVb1mpEXMAbqJmse+GGLG/Ja94pOfwCM/LT5sOauIDJSJ5F
h9056D86LThn085XhJHDmN1zAUskBhS6rK9NIByLGzlXGY9euJcs4+4T9zndrmX8MK8VF4JKDzlf
9NaoE0xC5GJORnC76CVYPVbteoKE7/qleLmMzvyzbwemXL1WEzNO0UZt4nud9Qso11CRadl2WhTC
sTd/pEzan+NNYnkGbeOF4bEASLszbjncB5gtgInWZ3JDHfO78cPAqY+KListB9H8yqByuGa1vHJg
yPSYeuhCGGgjdWd7Yw8NT5SRVIpmfhRvjVJj9YShcqX8p0VK5diLQdjVpsvowL+tymKykY7OgDIQ
/iaiSQqCzb9OJkJxhW1mUWknqxiz5aj2T/MpjyPeD/VNd8dk7KsLAyCUyOQxK/nCq8HiPZ4dqlVf
22GZ4MKjdoQMfXyVAXbzUBCyB69Ehc16S85G6kkg75bRL9PW+ve+HwoppbnLkJSeIknRW0aKA4yq
Kzde73bHZaXrdUi9qMRseOMObPTpB1rjh99M9r0bjWGNPvmfckJUW8WGT4wm/eBQ1U1jclhTj4aC
TvHLtdVy89YQUrJixohwOY7QrF3xZODJv3wFSZal2vx37fVRb2YxaYR3+9o0JrPTfR2pb8DUfKUD
0+Z64WO3Q+CSM6uI3MxjKMM/+sZDXR13F/V8bn8naKzeVbBled7Nl7uAde8s/+NF6LirAi2Or3al
gmiM++/3e1Y7r9LLGySxHVXjgsJUzxvVuQacjFUUuZo4EWc9bWN46l+IuBvjffDVHCeRK5BUEaq+
1AqaqSeUsTZYM9+CS1JAvizLJkTTxbtucGjD1mj5QOhu0omKaU1yrhmgyFG2elf0Y6fFbGigtAGm
WNz2l68CZjLitmKPg9pjJ2no3BiRqRjxaqW3JRxerWtXobH9/tYRnoXyJy3zUSco88Uss0j2/rd3
U9VNCFzY2LREqmj3Z7HkMhbULJ8Z5cEwMyE00+plO63yi7If23/RXVPTt4NSMl4Vga5Nt9B+IQ3p
2TJhvRtG44NlZqiyFw8eLTvOjVthsrF8+btrnx+R5sUSJSkdwNrrK5CWpbsgb/SXX+CuQKGpy/o4
d6XEM4CJVrSgoXYNRBDMpSSGEpwe1W4kS3cAzuNCUOWtKNX/S+5bAtsUQ1tzaeBMzS/MsvmNUnJx
Np3HfCQaKX+zOFPvorIEetKsRAQURFDEiTBG11kMuSrUsi7z0kJ+/eBaqvGGBIR2RO2WLW5yfjvC
tfAnEuf3/3w7jmRz44Wb7Oq+s99ILCc++pWAwb19MtWyOEvlqgJJKUSVZMean85G8mdXAVYJ8QMC
F6Yt4Ar6DojHCzhoQwt4aSTBWIOA1IOA3qjHlF+UI0YJ50QdHhbUcCPGlgF/0yJGA4zCrncMHVqG
DDN58yoiYx6icrlmnIOHwQKbKIQjbfzFlkI/OBaAzq02vj8IE3uAXFQtrVtYcjHE38JF5ZL/wwqu
/u7+/czDHHPBoHKDZfIfrbgDuMJzTfdz3mpeXGVAR8YGBjMYL9GPy14G9p00qnD2Qhzl34g0vNXU
dPDDMva6H5GNhyPNudXyODp25fdSsihXXZYo7webJ0ojAau1l1ov4lIL9Hdf84HeyD20kJwZiX/A
Wuqhowj4BRO9+iRHjm+dCKPE3KlIJDkk8+oLByuBXwRu17z4TVHpqwGFCk+uBOBigwSIw7NRTJpx
ozwzrgd1e1lKFK7Hwahv3nGD2ioMfK1FWE2faSJxfOW0qLuNllgcEj5xWMnd43lTBnCpTPLTl9mC
wGTioAn4MkZNi3BqBPlg9lCA/g3LJizr/ke0+UL4Jq8Y5eU6TMmKvS9aJMv4DoNe9WLnWNkP3Qoq
sxooIYjokeVm8D+WKBEBhajMJuRWI8YSCmZbbp7V8Tbfs6Hqtf09EyI68OLxMvQ2SCuLRFj7C7Qk
nSB0+po4Mc8tRdwP+aDsH3xuaowcHHMK2rCeYBAOa2seOe3OIeypiFeuYvNqDY2EmlQCftOO4kRm
a1OH8Hwn/7Ox9wNSEQcqkXPRRoXej4WEp/DKH7H8nBOC377SmfgGDCVxfrcuBkxWvoY5jWzVc3Rs
X/K4SHYEgE6t7zmT8WFlu3KKr3Qpm4fmvhS1HDSZuGzPIuDHK7m3dSlXIQqW+HpQek1+xQm5CLSA
HuTNpwlloX0SgRQPJba+Ho3gSHSDcgEMbIYtCtB31Tsi43zQ9gSHpTxhVG3j8GPRGzHGFi9Mo5Fr
LJUuzzvPEcIEVCEfLXziPg/QzaPAi+rsyopx+x86PmOIyGB3DeSMo2tXfuBe1i/WKNL8BHNZPOK+
fuREuKx8uPvwVX9Hl/h8CT6oLGQnmNrssgtZJKyl/aF9Y6gGL6nRa8Hn0AY7j0oQ875PbXtcAERd
uhinmfxWMgZ1/dDmnI9MMOp8UBtf9u/IMY83W9nwzH+UXsEhXDceJnh7nr/hsn7Q1T8xKu4OA+Ly
4MVAOvkjSHJpf3fMPRuhKVMrzYFJM6qJpVJ4WTXsnK6YWa/i8J3Y39NRdVE0R93MAft7aWrcUV9Y
HsjvrBnPfgA6+4+FMFIDZ20npFVkiuBvx48StRH+f8nx93yAHBP67J+HyErnq1IkohiNl9xQYBbm
OauhXqtY6Kc0jo+PaF9bpZydEMVFx8Tlui/7CTQ5cPoCYokxVe+vJ51f+ihcoy2nTOHcVatJa+sv
+yp0xpTsjRkUBO6aZ2QxLOlfa5sm60F2pqluyUtGzCH7726G2YaG3zFDsZxl6sd0EOYjrcFlx9jR
ld9RNCl/4MQe7xdA1kjXEgvIREM3l5AoBFs+81K5EUY64EU9N+Fkbrx9yzqoE464ddpSLbz3GiAW
PkDhEZoXr6EkgjX+JVU2dZgHJTbLEnAm4l4S6v9dJ74FLie+96lvNoOdUQ7No/dBikY89zGgKyDk
biJq3uFLc4RTcQATK6gv7oq7xN9LZMGrBJJ4VzJlcO5JXmZq1o32yIXJ3SXEDZ+rU+cJP+bUMemh
hELnaMI8ZJagaW99H6ZT41zRUTA4z/ckKIfukYQmabIDlEAOHjVJV6+ygcqhFAQeDaWy7+Et7pEr
NystokE81VJGjYDcRg/rYSV5EUr7AHrVLvZgLZBqFQ9mgvCbKJf0SmzMzhyskoEI6mQGmK6pqyLY
W4D/+Gy5hFnx54NAF7oOduyER3EM1X1F/QAmIffPSYuz1HxO1WiCs/aEfDCLby0eiJLkZcfNDE2b
MsVPn711wDkLmwCAxv3GiMc7n7uSA94B3mDAxvGTxXnnXPYbYNzXYTXhHymDB2UuoB52XjQ2/LM5
/AGCrMBf8wJaIGfYQDE+zkB0OqYD0CJwJLdTP21n1rmz0zZwEBSS0756OueRAE31rBcVyjuk0/T+
0k1oXxcUKpegSTkuwymFd0wHvKYXRoG+nBDDgD9lNun+troQY7QINEP0crwq+3PYy4DFNZ17Lhz9
jcbR+cDpxtcSkZMQT+7hnkqMzOYz0tOMC2G3e4+n7cSxpthIZ9g4CQUkG66rNn4Kbjae5UYaJIBc
CV14eVpfh3WdtaZoqOYbWk2GXFm+L6qsxhKb7tZ/stzyQ1NOsMLoXArfn2Na375W7aBtiKRWw5Ge
GWCOsbMhNPovb2uD6A+AisGsevE+IlvL3DHuq0bPaX+yTUwucryMkzprYI0puPxN1+BRNI/XQu4h
fzNG/fqE3QN+9tCRvMz/tWkXHEPtH6dMfYUhfpoH80l7wb6TvvTxgzZAHTDVgB9/QBldRHzy9vYb
L6jHJtv4fyE4wB/dyplwe1VBFtaZQzt9ii4g6sis/CA9R4lDYjopnCwFP/4kWHmYp8dYQ1zSaJuk
jySd00aehJxpMqX3X5XcWywYpIT2QfPkIExvd59H4P1/ty/hKTbOwKjws1aWgtXU+TzPKYmjtYjg
3NZTw1jdXBjKxgBQFNuaGrt7lFo33/PWPiYJl0TDh12ORVYYVrtKQih4c+eTJCfFuUqaFjI3ELh3
6jkwgwZiRAuz5WGtCTJ1lvEqZaWU7WNuuW/6kwVGsXN5oO3dqmZIeAid8wsBh1Y1m/+U81OKzsEW
UaB3Vj1ojXwyC5Rd7hvb/kBSXMX1dCD2juAozgfXGloh5z4h5DUvvkRH6GWtm+fW750YBe69uLSz
pWOSG6fPYAaNB9uTw40Y3CoshOOoHaWpvxqlhs9WfSRyVjF52OWQ3ouQUccLrJ6xipuUAkmkkPKD
27gxwOXGbdO6EiEtpLKHKhCLxoQEEEKesILzmAOATLp6siRfUUhNKVhfuVJYBVNTXt31pCH6tu5G
/c2M7wNM2reUCVXCUXu8bUCxH5kL3ZnntKJbUzICvmpprhRqm0ZIDFSbe2yus9SVVZCed6HJV52P
4+wpyb25crATe0EIZu9/IIS4jSne3yvkgbkc22wxi6Zt0S+6YQh8Db6B86fsGBJi8KirICLCzutE
py0wBqez49mWNwgxCKQfEKkM4OU1XU4bAu+XVsXeg/DAcZUD6U0op3jwtL6o25PRcTWDsPXdj/t/
W2XGBgaybvqHRp3Zzya2TDVNgEyFbGIbk7r3hDYVA0vF4KabdSVqYgdrj/rKq139ObhaziFjEPhf
IA0c2XJntnDOkBEZt2WPf6N6DYAsi3yBuUFzG8NJdHC9GZZ4TX5r9Nt7e6zEteRNf6raAKz6m6oM
s4MBms1sshLzgW+d59LJii1tGjoSWAKv/0+3hMwito7ry/5TdNWtYhlbQPae9IySIrXqRA4rgu6u
RPPoGymSnFcoFpzdP/0I0io8VMuf2R6MiJzDtq8jDcDrMrrjYBJNd1F+1yr8/N9P8rcfZD9V+xgs
hK0OhdMOXURzBUL1V07HU/MprJzgRhVUC+vOTWMGBVTg1TqBMTvfMS60WJbkX2bJruET9T18+sNj
TrCtqOkLX/H8KHhSCz3A7JJKxJDeP5tfg8b8/5ctqA7tt+9umlwvUgwdZEMXJbwnAlLdCTv25qfS
3Gu1PTfRABwC7ZAKzw5Ps+HVRtPkSLukWT8Zz8JZPWAYn+fLYBTFRT5SZ9rmlPzHQLi5Sd52k4rN
1wPvlANPXYz5VZbpgi++BbXcu8LKgmMlb1UZXQcz95heJ95cOJRkyEMZnnNBGakcqzHxlbzL49sJ
fmnKDMqzEkLjgZPv5SV0bxAdnliw7ivkKxmKwjbvmMAL6iSx1dQsIaWxn4+abpFIF+ItF23vDsQF
yA9I2orFCivV4d4CPQI5QsinmSnODEw3GzRx+cFksAn3GSDosD5cbFWbILRZAJmwYuBg5/A13ek3
6w8CbkWExAIFI2NEAjdNJ0sAdT7+vPFG1/s+MBqpbLYxw3LuyaT2YMUP3xBqTy/RBMpp0kwrOJds
1qBhdCqStvog4r0gH2s7nQxQ4RW8a0sSeYgqUQ81lD2wS4ZDcYUwYgHagjn/MtWxwqffS6OysUi3
wrC0GuCl1qLU/j3hLmd+PGzRDJ+Cs8CJZW8QceXmUV5kt014tytD7kzZIkikF0hQL3E0V3UGGuUT
Vrc059zuXbZh3ZXWudhOyjsKIEtuXLv5S00jx6U99xroSoXp+1572dT/MJ3rmHic9UTzIi7hvMZ5
i7fnKhBtku9GzTJZHwzbLH9AVgced6rnaZ3A4W7FvFoNeWgCTK5e7hTP453/6rFMhQ/HxVhZhXfq
JlJFv79ikTL5bIGcYy0ybe7vzu+0xNmXMy84TnR+Au8kFc53NL82frdf9S4EtaOANSMmOHS76ub1
BAN0IYOpJnddXmf0vwl97zf+WAcd7ev2ffEjS9KMZVf8evjn6Ih+SUfQCvwI5ai8fUfNXDIXgwP/
l8KdAaFucMlkKa/AP93ZmZsE2bN4VEmK0sk3XuX1jARHm8QcoP50XjHvqdXukJSBVA0wt0eicJWx
PwgE5iKlWSA09J7kz6TKXVsY1/iLkED0VOMj4M/YCOsG/pTaRB2vSJsIPrxpvS5un2P5Y7DeYR0C
LX0FSbhkDFJmhfKXLH6sFlV0aEWR8fUXcPGct7A5NEHZaD3zXI3n+skbUxvFhCPkka3peKJ6KKyJ
6or3h1hocyM1ZxzVy5f37L2RHILFHzsEaByfjYuw1C5k2zQzCTW0DZxDYgHw4lmsyOmPP/lPqYkl
U++ijdYfwO6RuQ120G1+aqruHZW00clCCIhabagk/l8z3IxhfW8xbANIRx0X8+kmiyhcimi6lBPU
u5VfKqRU0PxHVkGq++QEpfL3T6Yz9qz5Y/HkBjabn2QzwUoL//c4SvSBpi5bKnGJKmhGVJ9X7rQ5
eOGjWzXrelw7AqGBUU+wEh92P33y9SybLdszt3Zl9GVT37F6MRkVIqjbnX3BInevGYjUwh5U8A5f
N5MExxtWZYxrssv0nANVOxirtO5Jxb3Cfcfa53Ap0DCotwPKLrKBA8Bj77V2FMzvWewU8QURX0fx
eWGwTsK4f+4cPTKMfP6gW8WWX5RUFHZRquLI/mgZ7NGqNZQF2rtf225kxNcGfaUHgpApoForMxAs
1Hhe2A2RrHgCkeekPgst1Bdt/1ZWxUa7Q1XkjlJI4BqkTO1e295efOapbtaKWpNFSyQjUWkwJPe2
zgJE1JuJ/S/inFnm01ajKiYRCXq924nSxD/okArr2rzxe0vSIdIJ+7keH/oBnt/dHO4X6OdxDYpx
SlrFFAnVfInlNNMplK67VyOewzt92vr9FkeKSBiR5Pg/jWyxsG0uvskf4kil5KLcU2paqNcHKVXQ
xfrQEallneT/pKIVI/WojH+YDG0Amne82Ao3z32r7EKRS/DwHGI7R+KDMc0ugHLY2miYyNTXRVyl
EQU2fW0H8R48kQ7yDO7vuoUfAJvCCC0FYMMBgxSzoRcyZ2zpYwGTeveKeo3JzQg52W9cN3LFRA7J
kVXozxc5BREMtgUfdr9jAKycbpHSxqNpxqAKDyEhAZ0gf6+oAHrTVuvAN/o6PNYdet5gkUL6+/qs
Xrjy9pZuiqWzT9EOiP7gPwMds/dSOk5+IhTBUdwOQP9hLUGiXf6XnkFSHsoC+hSOBnnYsdJlXoQ3
MSCrAGCn994nYzVIDBqcdbZPwBZcJIt3DE1kDOUg7tGKF7puqDT4F7D7gubM/8GoGPZ4zBHTsJzm
BZ6B1WVTn3GBwrVujl+UJrFq4vwfAMHmWwSn41SyFhnpHvXP07YfOkHL4kYHPVRQFh3BfJ83ZfKv
NFXSnOYgriya7LOXxncEopmYooNvk8jH5KQQciDFfl4RsrFihTqXSqIArhSbIVJjVLBC9SlBSCPA
FvzYLcUvmPoiPm0BFejLg8mOzLJIcHIMXtGtUeFDCeWCPAh3pGGN3/mz6mDEweaOeNUe37mJUN1X
bvHU8LUXoTCW1FLtQqmwSmVhnVOuxa+Xb7RZpVmzdSShlMa2Gb1wGUo5cmH7dUK51T8Rf7LEkq3f
SgrDyakFKxsv+p4gNYkqJIEuc6QXs/6/1yShbv7z8kB8oIOKl30D6rs4MePhauZxtDxXtfM10DTe
85r0q0e63+GF6DIOfgvqbR3HOLYEtV3wQ1tjWcdRP7oNBK1HWnLq4YoovpFvCx2AEkpUL9lk/Dmq
Hvmna4QgIytjw3d3Kx69UiI1Ekt0V6u787ZoTN4llHra9mOP/uT1j6HSdcEixMdLIfrZGmuqZgNT
2loUlakq/VK7auxFQHeEIdYDLUaIGtsra9B/5oUrCACH5+LkfiyobR7i5/kWgF+tdL/zHV5w2V6Q
r7hCheiZr1DC7TLZdZFXP9ZnSIFEL0uH60ulfJ4bccg0HrdWSj5zGA61LFPquziyCyNKeyrVIGQz
N7SF96/keq7JeYBeoHzUofzZPeW5gnsBPEBNKUzHW49jBFOfCKMPSGNzR07uvxyRcvYTsbERBsrl
M/q1wcHHEZrD/S4Z1n4EgklLG2KVfn8BjIaHOHBEFOXGeaqNxgcfShsOj4UNSxIzz4W3yBAChveh
GlAzXIK2IhUXdxzJr5yVita6xv6L9XFy9jRns08N4gDTzNHRQ9yMJoo00mbC0kXYYCcskISF/6OP
9Fohob7yD6MkL7PRMihBYtQ4d4CVhpS187hslReZPbslUyfH1cg4Bp7+b6lPcMO6f68+RduehNle
y8eE44tf4CChur3WCUGbOp8KjTJ0QKnpGIegJq0L2WCo+m0PNgKzZoNPnjwDWVWOUcNN6V694eby
vVkqAbZM3018PXRuU1SPpjbMRAT73kZgXGFH1wQWx6uUC6ns8YCVtVlYIoQnZeEcr3LJ+AIRtnGY
0BF2jikF0y05YQ3xVv2TB0a/HzbCc+XCTyXZ2uW1uf3dkDem07bn1eCMzu2OF4ka77xP3GNPykkS
V5j1vpqibp3VGnmMNpn6XHnVRtSk//fDvqW5pYWhFfRClwNMXKX55n5lepTI4jysM/j03474aaRe
OLU5HWZ7BlMJUNajpmy3uWcj06Sxn2j5W+o7JTd1JnKH7Hk6/PtLuvF5MTWSiLOxgQUR+4J5J60w
viUOwJVb7+1LD5FwVLveSu3IHobDtcEnpw9KiSevoAaFqCZXw9f/Jns5C5iJEn6TbFoH4KfMtu67
Wz5tq93d85b8yzV0/R+7J9GeVsYaPw/RjVyPBYqwD3xNTvaOWDJUY7LcTIq924/vJHGzyVtpWUP2
v7bWy8g+JeAdJ4cuKmp4/geDxTpOaOjS1ltR71qXxKw0qag97rvzXpLo8pRJBZbu1QLeQEmJlMgC
sF+hKYnGmH2Pt0HRldTj/14EP433d0FafzJ1PLDSLbZJvksrFdiMj9HVzRPoqWsymSqXzB0gFa60
MllMxR3FfTICN7vdDxY5NQ/0pQmd0OrKZAG+WUqUXFShZIc9K5CIEa0G3Wq4OFM5nlxtOjubN25l
bZDn5Wkw3osvne2GZuFqCOpRHOvqFpfGN7B+NznAZ0zSfGn4NZhr4dyOGZFeqkq1PnrKPbwivMU/
OHnhfxkt5ddBLLmiyfYHn8Ye/rJBKZmLxlAMyQwXVVHM2OH2aRwJ/4OKeO1wud7bzF1H0a5R3vA4
czSAU9jNNoPOSGRLsiRTB8S5FhzXgIOLi818MDs2Ql7PcQ2ejWlhrYusDllOW88hedTbJTLyXnzl
gXmcnlePGAg19UQhmGD6x5AFABG0eybilf1lTer/ENVl5iaGm7MQurnZju/MdBHHf0BVYjmyZuCU
lhXCXa3VxUhdDYs3vEqlpTy1Z3WlgS1YbxKWRdYUOC4NVsvjwpXct9tqzhq8dxqjntrA2F9MMIw0
LLxWRcb01XYSVfTzdBxux95vW/+djc95zdi3B2qkl55qO4WIEubrTkhloYU2BdEkX5KhgRGfic3M
wGuXK4vimzVsbjrv2rzXsSFAXizx1rHvUL9RGwt1bAoi7CAw250D3J0GglYPisGQbRMoiSmDNYp9
AMHh1bYiM3airwIGV2baG5C/oqqxasF+98uYvwEx80QVxQMfMsxyJ5gUIWP2O2w9CXxk8jRdMnX4
EVRmbSCL4xuTEQspxydoX3G2Z70HlUfqDqzd32O+ldV4x2cJSep8xs0kRVLs5aQO5DtsNtqVLn+n
Q2Uik92/p3R3hQl5eHLfB/kjScGZFSFxUIOzDV4KK8WDCHsMI1M643lptPDpLYfl6SeY80a+E57w
RR5j6diSdUKbQvvKvVbANfMKam7NZY8TWuRRRHsyx32+opyRs9nlLrgwxYYbEYJtDG+136+pbDja
Zt7RZqUSh/MdA4FWqRALF8ikdgNKL+XZpTExLBm9Qd7orSV9t+jDt5ZYdKWNXang4AVdSkz20DaN
3e0Gw61UXb16x0MrS6C56zYx+D0ZiTFOuxrJxUbf46CwbvNPfhpKMyQoai/Vu5LIXoXdjlufiUUy
HkgZicJFAPDOPdZmJ5NpnJcs3itr/YwpuTRJZIX17EnuWyyrZpY4r8R7oKobmv5+MN8MEIBZuN+J
DVudGpjoyyG+qGZCMQ9PVZOswwVYq95nPQ1zSDohacpovAo5MQjicsk1ajSJ4rI5+ouKL8OZB8j6
9gPxNM6HCiukjq4oTJEbyJB+hl3cYZEDMP8/TggWNByBBJf+8BRg38mz6HirTZUqUFeBo0fG1OOP
XiCEJQUujMUgmoo1aDGCEYwjoqwPVGTsxFeFVBXVBBFcpY1dW5//PLLh9hhM3ETL0rJVAmKzCgNr
L/Pe0z5CtwRFpR79IFR9mdqKLPOJF0Wab40LYDaDx8rZSsTGsaFKPejnXNvrAyFHwnUmsM0hBz2a
gWGjykxjVN4nDPJDcp1x0qRjw/DwTUEghaW2r/IeRseQIo715tY8+iJHPQYkgRuEbNpqYSovF12N
Ujt7L/n+ivX/I2uQrPxTXsDr4UMPWtGuuBrsCA37r06lk5xexLMtX8ol43tnKia80+fqKwWGQYuD
4O//jikCZUMUVIlsghZsnE/lTDoCoG7wIvZatKSdD3W+G0jdI5tWy+/GVLBKngkC50zo/riTkrmI
Hgy8fa9jbBIsIcwFLQhtPpxslvSnCmZGoK8B+o5OyrjkR7Uom13L4/0wq5UOgHopn0LtdhNipK0/
OansaWLRrBUEb7izCqfU+hRFRRoZIxssND+Si+cJreUKANLxM/ID/bLAzu2rzjMNhddvABY5rRJt
X3gjS9Xdd8ZbKYBiMPjZqxsyoTJPnbcFPNbhai0m8hZZYwitdmruh9uRwISrmZqEndEidbGMYytl
BaUL/aVhuEUTvKu9Sq5/10MGy14SpGD47hulfpaqkQbRKYzK+UNOJC5Ae1X2a6vsTADKQf5IiZGa
epnQR9KhWFIp3oUOKNuNauiPySastTXuelJCkP3cyAEK/53kUTSjdeCNNkoBI1C2j84Re+XOH96L
FWMsmbnfalnpPfMQy3A2GgdZu4TEbxX+0yaI3SMH/n/Gbvr6SN5Bb7am5aQ0U/Uy09AlX7aD7nQ+
v7lwv55g/8vduHg/F8qDdO49JwA7tqBKlA7lZexhzAY+8VAvA0I8gqpJMZ/ynZ0gxksv2S+lCGbW
IhqgJQCv2eBEdFo4ONEs39bWRT1b1j5Xg4CbYyW3f5ETUVLc+hYML+gvMonY4sLxOZO+rofoTFW9
DcgQgrpUy9MwcQLXzF12y/FokVEdDd6LbnCXTYK6cV2MReyMue01Mo0pzibsE7NPncO68jpz0Be3
NQzTE8kKWdohawfsdk2LeBI3/PR+ocEKSqowjgcgO0Gd6ybbqkr7KDH0QAgJXlrxOEVTiRejtuqD
hRBUWFi8jBvp8WbrRofJ8Pg781AtWtis+OVzE1r96vOkQd4nDnDHh3yfIcfMbcn0iDhHFAAa8t8f
J72aIIb2iGoPotj0vw9fJgv6I3J7uIGi7uwZq6xSt+4NnXbaKSfH/ot19UMoUOsQb9Ps4gdM8Bmb
yFcZSFoT1xIROC1t2SMwXc4hqn5OpJW57Qmn4vSsh+MVli76FY7JuKPWwZR//pY82CKrvRV0W+9v
hg1sJoA9Tn2k6MFd33Rw5G1ix1F1ZOzrJZE0BHKbysb+Reew9B29ezydHUx3HZevWI2FTzwwNR1n
k+zz8lv3JK2jXo7nsam+yoPJqEJVrS5TZoTdCpGqnUCVuvZlt/LIrm4hYvsaDG22DvO4p7/fYkBq
ZiIcCFggg0SqYAOuoTo9zQqNFgN8oY+6aKl5eUsM8yUEQ6NYSULnmDTxcqu7YNuaEc8x8tfmPAWb
eiUQq8ne5XHcd/Vid0jGBSYvQypghXQBKetSPrBCcO+pPy2tiOSZ0d67SA2A6kJ2amzdL/rjGb8B
ruoJBNkfQGF0D0xARU0iKzzT4FT8sV+Smm3y1bNN3PbDvIxzGQm03C04I7l0ibvc2kHTpK0T9Mp/
HlZy1AGwDZC0FEuGbif1Nxw0xO8i/G7YlCR/9+6MhVYfGkUCI1m5hBj1LSVJL482UfvgJMoHTe3d
TkV2M7Rd3hZx4a0TBu7tZKsABSTBq+3pU6rz2wtgTDpLJoqkJdxgXWmlY3U1HqQ1Sg0Iq627WG2T
FKh6enn8lwwphVZEGE2tiHf+9OunGveZMECIiiBB5O9BkjNKt/rTIURSHBCoi5qfWpCe8DK0P2FP
B631BHQmZIFG217xC4llBJenmFZKU6AAXVg2KdAUwybSHV17N88a/G5cK4xABmDO4Gk/zPmmJxcQ
f+pWrHiiIvQDeNjhpHbpuLaGNSnOVFsXfN29SB+4QVzf13N77pIsYdflDp++PXxeNRFeWfdu7DY3
kCoqWM/3xJ1am69UgG/xhxAHhPODA02qGwtkRjNuGSEV4vbSQjow5ApGVlQVpFHQ1p/bJsmdELKR
FylaAXE6ph4lh0rECNukRYmbbtJdp9tsr56WKtveEF5SGxEeFF2HHWC+w6B84CC9XpXQXEvKY4R3
w8ONsaePNuldkthxM44KjVhB4710VGzHrGk1qZGargJ+2Fe0iwH5SeMIGbaZxnmeGIYpKEWLQR7N
zxWQTONfdRqmoGo5eNyPJTSGnJHzsVcrnCHbAL2KrgUKSJrLZeJkNnNWt4vo7hrDR/kIaSXgzX2D
BnKhYi4UFni13Q4vCtzr87CoGAKfimr0mDtvB32mDvT9I4Ofg+SB7Furcu63oeSy9jCQtKvDJqv2
Es88T48cf5Qojfw4SDootGTGwODCa2IFxvanUsrMSCG5LkVzZxHHV+RjlncCBwzSTMPWfJWcy6OM
NcD/YrX80h6/t/NiwVTCAHi6O7ILR6cT05L5hseOxGF78Y+Fej/LAeNOWqoCjRopdkgJshi+r5S+
BVmt0rAJle3Pxj0sgaaXSOlNz1e1wtQrjxtm9PYaOpQ9CIFBmT499/UwzBtPF3xvLQjhom5l/iCW
znJxX33lGSgqm4QHCaCZPZ04Y489xatEzanQOKs+rdD4Q8vCLYgQmPBLiGemxG70YIGzDl+HDhZz
PpQe2YZ6W4+zaXmxY2mgWZWrecpioi5+1a66Y2CuHnfd9Ia11Z1Ifl5KIR4frc275lyOMM6fi6DW
5v9MKbCqbSoiAn/Ml4UYJE4zQiQZ4TnRKXYEUXvWGgFLjUCncsthIUsSmXYAP5PALoUV99rCdwat
p+gbOGBbOXJxuSMMV6CPiDWzbtxYxTDEJjeF43yV2rXut0tn5f+lcfS8bxnBR9dmDphm3g4P0RE7
JWiugI1FuS6kSANnzmAVbLNRjxodEjkAaf30xUXyIHxjw8KbPJw78Xo7+vPV6567GyDwC8LUa+64
JS3AnmC7GVdwJLmFmj7qmJ48HjCdhwphvfvUmPAo2Rg4kv6EV9IM1IDrEiIZ/CAJsbnW6sGa/Uqf
tfe4wff/W5FudRydx5l9xgRYosPnDCrEIpRRIUNMDZKkPphavD4RH3IOzI+0d+fkptswuBbbz43v
YPh9g0opabEF/rLOKSnOJi1vv1SIRhcIt7Z5xaxLV0IyxmcU1iLPubdub0cWBM/vRBd0x7jB4LKO
/5RhJ28tIxW6dV9mwe46qz2hTb+adO2Uwj/zpcCLJjMISdcLZK2g1Qn1crX4CdGN/L/UUZND+615
oXP7x/1NkR64heu7mmN+EGBzAuMz7gaKZwv4r7ip4XL5IvHbkrvfS93uGoVkGu7bC8hNADH9odWX
7hb7DdH9e7gR+j+255zAtvxWPjLI8RsteQidlHIgXUnL2DudDm7Y09xrcI2r3PyizN9Hc9q64YcA
xVqcu6ScpSiKjTXFyqZj1rhh/U1ihWi8dKh/MaYd+fVN5lW3He2ca7pGRMFyfw5An3u8hrt/cQLt
hQJklhYNOvpXArvx8eYZFxqhbLXwWxXhHR4MbAuKyCemWpM57N7/Pm9XChcffjpxu166aKiUvOpD
K35m9+DMj/nyNtxkBPTbgLwUVH3NYV55IAatl27NbhrMvvv0pSUlIXzLhEvTFxcd00Fy9+FYH+fv
aUYSKJhAaata2q0A6GwwfTkKoV9DsVqKPchzd0LoZMgybamqyd0wGKCQGlA12pnPkbFZy2RAzU0s
b6IosUUhM6nfisfN3vy4OzXZ1ir3XraN09IX1UIesxgEswswXnyxuMKwq0ZbC+an+RKrTHCDHCre
xkaGM2uBiCn2frt/AHQRI0m/kWgMl4HHN7+AYM3FDFiig7+MA1uyb+AY1Ik1IYVB76mk1gYIgjel
7N3wEBC97ip729HBvZ1080Soj4ZeRB+oO1lJyQNCmXdSQjQlMd/s9dRwOglod11mhv/atz6wRQd5
/YP2xjWAQUOlQBwYtczfzUNxWW0B0SKI7Fl5sSMitH8/d0R7FD2kTkENBNMiibY2ZRR4mipb5nWS
cvhCqLMYeLM6APr+7rU+jkmdP0JMb5e9WrFCFrjW2DEKv+jZfSvin0WI1y+UE6XpcrotgJ4DFC2c
/DRpcXD4UR2+On+WlqydpfgNBdjlAfmdUE6zACNL/hygOJCmII5j23b3C1Igb06kwFMBb9Usy7ul
SB2JWXZxcUMdSuO+p53l5l98aFHCLJJ8Q4vsfWWYvzNhSQVK1uy2SdCc0tD37Vi/GH7//gXO2ZYu
M3f44Rzjx70RywZghP9IAY+1f1xGWWBU+/4ZaqB+QcIdIXjL5es9EWuKJ/WWpyeDUqSNvzgXMOv1
QrBchztFCAndymFhJEdL3EA3BmrY1EiNUNOz0I+R7azF/M4v85UPqjrglfL8RHk4ObAkZJrS7C30
AG70MdogbOP6bn39KucpmmDzB9E3MpZWf2QDzW+qfByBDpGnyXyFGw5yGA51+PFvPUy2l4W6AaLb
dDF5qpOu6sMqz2YHE0JIdzMw6Ne73VGr5cW6OsZqaCdKtTDir98ZeCk+7hKdqHj5VsCRsY7aI7lD
eZVlknhpfWxpSpM41SOJ5fR+vnQwJ/G2k5vh4kwX6U/N3QyvpjGmmfkM2DETdz1NIh+8dkoQ9ocO
CuH9kavrRbbQcLVy4sHgMiAPCW4PIud05dCVFy9Lorg/c//7zYFFC8IJAKAWBgFSb8na6DIb0A+A
ypWkQlIZUQbFDwEfnAu0k/WmxMpM2lPQCd9RZfay84Lz1ZXqv8V5gpMjwnN1i9M98ek4lUSAW3dp
5CH85YuEF2xWBwLjdd+PRbVbc9RQl0DFUp3cykzO6r8ZUEcT9ZnsSI2u6DveYuyVO9mdtm5Q527+
/egANwmp1IH1O52oI10JeAhWrO1RyeZakUuuNQC+47VxvnD/ryCSOcH9znrlCaFdGvlcwrP8QCnt
NNlbkbTI8GQ7LBbW7SsGcArgE6oJDI0pYBzbUUZqAlzWh515mYZ/n2Bgv7rbH3lwTL+ZJK1ocnO2
parmjPAWJBQWDQ3ylkjw1xRPgLzsywPV5h5LNiBnMl1KRYDwdz0iMhCktJMuSamzoubjoNnf2fxT
tmHlRqGHKg6EZVmtHfhyYV8pJ1KgWxp4YQT54vvjUTx/IuY05txoA7cp7UWPtIbkN/1xRvvaSev8
m5D0j3MqhAlRxxEha5+TY9rKxDxWQ8zktz6DN24pepOAWKxCBp/G6l1CvaOnUNHex5qN/QoQv5cT
l2zNBjEDZZsNe7utElGtHTMOTURq3s79kyTQzet5jxfNScK+B1wxaI80eCTiUqklPMb6y54Gp+s7
WX9WRgqZ8YQYhwxMUWsoRTzod+DqfSUvErItCdv1hyywQ4Jpv0XqBF/I9w/Nvo9qc+3eEd7xXRSb
wHYhoH+j+CPk5aAMlDt2qAgckrSnc2gy4Z6hOB2iT99tPAYf7lr0yKNcA9e+f/deGJY7liK0B3oK
AciGpaPZKJTP+yk73wUY9KNJPoQW/iIc8cMCRiGyt2lpeP3DIph5fZhoVsARrHPfrlgX3k/QcAd7
4BgDW8IpkX/FINiwixo7vqDMWHDhldm/9NtBdvSQcWtjWaFY7kVGghIdWMeVGg9vCT/8CqB0vbTs
iAtusVHsQksdo86Iv59dcba3RFeu9UEocl4t4Gl3uSUDYpKnu7wc0tIleOIkIZBKSxhusbxufT/+
zokQBMiUkNH4AD8EBAXCTVlvg80iMC/5HYeic0XdKz16GauawQVqg/Q7lSaWn5FFnjCTAYykOcLv
/vLwSJsoSa2rvmYI9rF4ib2GSBXCtLjs/6B68kaVTxMWonw4yb/I3RgPQFm8x7H6dDQfvSJ5WnHW
zgiiERkGnmAuyuaSPDMLE04ayTzvNZu6sZjunxtuC0fXn+6TDXumjwH40Q5NmZbm/OEidfsD8WUK
jtTxshlqVWJlvia5qPuic/MO9L56Umc+hmp0IpKFs7evxG2Q5jtnrSbAwStmeFtv6iVz/82oh2tH
uiqRSnSJmAbx5nKV5O7SDCmQ0GNB0p6D/3b69pM+SgEbKg8JOwytKzdRuC0UK88SfsyhsMCzcKop
m6sL3cHZPyVVRyHC3B9Xk5y5DgceSJZIRPkF1oDVTX9vUasvYxidpduHiWWHtt5KcBjbuwp1IDnC
lre8d2Hb+IB1988nRtHDUOGpSIrDAcjm2lqnsa7aWZm9uUn0s1kskLfJmInurcCV1/+6WxLBCzOC
el4t/xr8XVShaFtMHnCNFvhiyLFJwNeYTl4H2KCtOzmi3zYd8+k2Lclpg7szqExRCyzyKYjnaa2h
EZcs9KugcGWEfHt8lFpTOCXU1nE86W2r5Iu0A7r/he/5iuzKbx1SWD09kw+ygIILvg10MF7QhGxo
UPsNgluqJ2sVp/1E6/4v//ASCRjU++ZfJjiukzLT6MxzcCxvkPaXH/c7arcZ0ErAx44AI7a0WHeC
uw9aciHqx3HzZF7vRAOBHl/mCN6pIZjIDLIpALTMSEsO2rU32xnWKZEkuzMkyJMvq7ggjCDOtJWb
Ikemx3/CINVzihlLIwF28HctPmI1X+Qm+PLIlrpNiGtnZTBcq35aATNfbJqcamBpV/ygAJ/p4vZ5
OGbCeU7E29f4khjcMLB1JWF7BDsnPmMffGwMVW/eyHXSDh+lqtux3zVb5uWWJ9pt6XmB4FjCQeZM
W+P9qW/bCAIoVnW3GvkgyiKNZOkoa9NR6IqgH6h4zLmz2YgAStzyKVi8E+JKp8VHdKrgGxKR8PYZ
3hz2uEKOTr3KKAAiYlegtRhX4ddutHLnSAkTdLjnyUgk8Q2YPrWkJ5gTjIny1XD/qhxWWFcyyyeR
DJVIQqPJWSPPd3y1JUCMURk6HrMGQ5RIV5cIcWp51Z/2TYEUCb9duxwNYvOmUxNAu+TNTVxqiJ/K
VwSvPotCcOJN6h3h/X7QRta1B4VPE/sz+Lyn6zKM2KQJjqyukoXxod8EvhLgAFm8u3y6PxBcHWO1
9LRce6FHkCtWPbPQw7PMpc71jxV7o5OJ0A6TnEIZmB4FphNL3liDO9vlThj5LSO2Tj9WJ6D639Im
NEBnu9bOwsOo2yTp5ID1+73sjwx1QN/ao265DlbE/ukqzg2DtyJtWy0B3XRM1oLbaXLGVWShhfQa
6nHjNY1W2iSPb8S0DaI+gF7VW4lItIxzu8ARywOQL/C7P26m6Qq07hNnoGcjp+aP6C0WDmrC0KCp
yD2/+vBBQBOc4ACpYHE4vmpq4OIZhOoNmX8k/fFrEc+3BC0kvlcptGrISkhpqE/87JLOfYBEsea1
3JfPDIds2k7A+zGme1FV/4hJR3Rgh7WCwFw4IPj86pC9yGZREpxPwcjbZyf5lBXErFMevPFwv+v+
yKXU2slKahHtXXSBsc6582o2OgBYSRdH1QjSQcTf9iCkwUohrcE5v3bdw1s+F4mzmIBMcvBxf/mn
1dNb26j2N1IqZE9JTjeiveFD+w4eRpy7I+x1IN81ndNabZUMgCFcZ4DXJIZS4e57AXoegXrk6fca
5Ii1DFzN3BsujSlF/QrkuwZijEgK7lDnG2VWDbogz0f5kRxPS+5/LgAATKF2PKdie2nrj66K8IE0
LS1KSnyV9HPKcO5ztRfQnz6BRDkZfU0bD+6usNxCPwCQKEc+tLESuyYmbGiy7TeuIRA8Ko8XVrRF
eL4f+dECXcv79DDEuqZL5hl399+bYC3qSPcYk0pwF7kyMbaTKjD4kjv+LkyDGrBvrtRl8S0QlL5j
9HXalzbnr2toPsLBmnwiAQVVW5Mxpw6eKtg0S2FGeLLg47V+fpheIbUpQ8n++4d8Ghea202Mq/Ns
wFGlaW/zdtb6y+qXD87stJ2yOa4e41b0NnovPiJqrp5liU3oIA5i+cuxe/I0Y+IiOa+dQug+TsBI
NpqoEJU6VfU1Y5VrAVDrc5UUfmKwilAgw/Or/zV2eelR1eKMW2TXE13nNTFkx/iIT/kg1UZhHFJw
c4bc7l8/gtvCRaApPVCMC6Gg3jK1uLOcyRe1ZZfYBQoMvfQgVGvReHZbw3wlpoo7ck1TG6cus1LS
7pJTDWUkOydkQRr5Qjk3hCGe4tU8HiZCcEYhhx4QGL8ON6aIEGisMgihUXksEgTcuX+nlv8OZkui
i+mCT9lgjp5eVxenBH84NpnPWwcWXA40dO2psNp82DDdW43aQLR0sVAEMy8IITpd0ZJNUjKBVBBv
P7lq610j/DpShbyCX7V4ovgSo49tZgKUsGpmd4a1MJDqG2tjTGaZIBc3ZqBfMi2M3mbLXrpUJXC7
SioxRiCVLqxOhOT7PxEaU9QgR7v2I6GkhKWu4Vy9Lzmd7ttkV0wZIQZxdiWKrRdWTXgZcdGtIFcy
Ew0JVw3M5/tBkWxRP+6DFhLVW6RF1kLech18uKK+Gf1Xcdwq8sqVs4ShOztLYi2Qf7Y26Cs9GYmF
xzC+6W2qHipWx3KzrOh3yC9IeGFFyLByIZPZaXz7bzB3Y8xcAlGrHaGUWAFvoPYouqduM2hJtAjo
IKy6LkjMQIgrVyemMnFMdDKDzTp9iQ3WaCxy9lb5tvtLhysihHkZPbq9sFex2QxF5NnQrA3cb0JW
tDVaj7Fk/k5wN/KRYQ5ExVonlMC6p365PmRDYmgvUUSTF0g9HppDAj3EVCL2jVO6cL2xgUfooL9U
qVXA8+u4r8KMpAIOxSpQCtoQW40GI3Ry9XZRMX8vIvvHG2/E3ua+Rjxj6AoyfGc2EfRWb73MYinR
csqzB/rcgR7pWuo7zmbBD2D0g1/ILs8E5wkugWbWpXlprlLoul/4aeFGw7Netm+ukc/n1wEQkA4M
Ux0t4FMPCwMaBgxjXfVLzGnDbp/l/NWMRIu6MQNJ0N7NAICizCceaxh6E27FStcYMyHjJ6lHNHPC
AYbuNIXetY/8Pzs9jLmUlK7SAptFY9y8EdunJGSLm+DuYCIa4Jhfvn4VQAKf/CLNssAW1EZBUhcV
AW/hFHBYRBj3WZ+DM08oi8j2FP3NzCg81lHJJS2blC40wJKaQzJ3+a1xvUDGfg3eEAwoyg/lPLgJ
MNmil6QMzrRZFDgJUXu+4dj8brtMF5VKL/TK2IvlJoJ7ZZDdqejunt8eaVx5NBKo2eKCOkXXdMwU
yLwMlaXcBm10lI3hVDPhOYPoUIp6ScyFFQZg+LCarRZvfAAAnLTM491Y97JuJKCVyZ5OmniWR3oP
ex2xg6ol4QvumOFYIYiIprLC70DtzDIZLXKEOlpilnKKV+dph965u0yicpv86pF1Ic7RV/zQUrPW
QPmknEn8ZFd4iPzLjd5L2dHHPUB4vT8GZwekscFbTR0t9wFar3Rz7gViFEHiFNMVR9iBCC+FEfON
EQ1Dzsj0LfWgbtVpS/TnaoiWcjz0dQqJCIB12JdlY7FdLpu2R81uIZPeRdMeZMH8gEivg1fpqG1e
TRFvcRE0eGVwmZ3MQenaTveWJrgo2yW1JynXfxpumr8csxLu0bkKyTiis/vfN6lpOlPamqcQGSNx
htlu9RmqwI3lG1eCqcUNvTbTzIrum8BZVhu5VnK5hrfG9Ow9Pl4d6/PSRsFyHmCLxvYh2IwWoRAR
ab8lx4tbuIFV6T2L/8Nn4W0QzzSzr33UfAO7Cm8Puh3aiwh/O0msEaKgupaGNQC2ynBHNa2+3vD5
qwLPdlONNqS7+Iv/0NImRE8Z3aADxBMI28M9fz4si2guCdG/CzDk81ThGj3CVR8jXOrN4G2DDK27
Im52eo6X2gjmHFNAKTc5bT6s6sQkfswwWMa7ltacyDKrfx3Q+I12WWSTWmpt8VNCmQHGsRTM5Njv
xCShpZw6F+W+N25evHiADUTFw/iXcQB3SbbL/6u7e4HDcb8oZ7KxGrGJt+yG+eoQMZMW6fb5sp2b
xdQqcagikK899vKhNCj6Anqqe3cpXCgqR8PH9FfKIsGzBs4Czev27wpBzqJnt7l6Nu9+rNcdu3ZU
V/uFgcs9BFcqG0jCq9ip+OHedEBfm6qh5SDLzJUNL0qLJB0MrjvKDhs/XyNHpTJ1DOg2kerxOls8
s76WRKuYNMMH6ZiACPv93KByZilMV1kbUXRPUdx6KfZXtiVNcAvmUmy89IuE+uCIhJyJSKYrv2s2
xBtc7I4jj7THY9TqH5W8r1baDqMfOWlHjJ5oGbNg2Rexn3mOBXsQdHhuUHLdo8jTKHJwtAMb0uq1
N9dPYAHXxFCRzYzwAyDImFHTq/k4rXtoTOcVepLAGBH0FqfGLku25yBKVK+tDYGykYFF5vUgI6kr
yrVjnOekmZ860gIyNTSghlRED8TvJ6n3G9u6d+88YRYqeXcU6zR2lkmDShdIgPEU0An7crCn9w/+
G2pcG5wpBU/q7YiIidSg1fqjz5G9hn3FyHKd9QEidyAVIfcN/Uwo0rw7+PYUxAIICB74umdJzZQ4
hz9j18XTCLHsyLpd5Al9eJQU8kdmVR6/mF/oewhuuo5EBmpau7tibef00leTJ8KYlEp+UUg6l+5E
crizTilLUJhG5NuuP7dpUtBukl9LkVvJsMSHTwyHKh4rm0Nvh9/fJL/HpyWHA7ROYLKsnwBih13u
qQeUIjz2ew5JIXwfEZlktaRfZ8Jo/IFoHQijcZOfEQ96X1+u8g4OOV76FG8kMMWMEe0A2IYTgoA0
cZNCZujSRsHyPIaulx2Tlf2zFvCth6T/tfZM2ISwr03js4GHeHEmDyufCOx4JuoIHceu/dKddvBE
YwFdFXanYdbYhPYX+MeqGZhRwGPm5boTqFLo+eNj8Ty1HdeFGyLOE/yJEbHMV9M5kpB4gjDJZZhW
zxGPXBVxuyUTih87SXCO3XvPytD+G8g8gG+L8FMMEEDBz+MT6mMb3LVHXkEMPS7Y5qgj+86NOKYW
H2tK+z5Kt5LmkRNq7PbsTCdmCArCdceiJU/PChbHH8beDZG0uHTd0mryCQtMUi3zA17MUUtkrmd0
ESwrMKqYqNZesZrShLUBiESqOKwMp8OcNbo7ktlWc/kw3KXD1b29IcX+kYdAu6mqXJSH75g644QA
GiUI2Lw3CS5ewqhZi6vBqSQzHuu3QyVe66FU5zf2P+DgDE+qQzZcsvlq4aF5/aw+GsmYc7apmSmC
Fwo+fHZrk9yOdoSi3l72K0ZWTbhXJZSJ9xmJfDFPF5gYFhlMyodZg9mXcLXI9Z7nuTkPJSb/N02N
434/kVqRuTSKGYU3bCRINt0f7H7jQoqUB0EtHUGQEKjajvxBqC7eBl4h3iM9FQsg3rF1UXS1nhWo
iaObtTL0UyxYhgDi15VckXEXSuCnCO/AqaifMXlKhSQQ/7kl4S8G+Ejk5jnEpqNSPBVjkuDULgMt
DzYZc2WM4TEG53YrgGHx77+I64jkS9x0icHfljqqaIuJdRQElFEgWYjjk3xNt4fg0w0DdkEED8Rv
PX3uHgd7P78GuY0ACKK32YqzLHhUIPPbiTu+NUQ0xB7yA9C1Ibw6E4NVEMtzNxwCqDnRjO93AEr/
Iw7hHgr7AEyoMdK57PQAhZbYFdNJtmNX15OMGGZPqp3cYRpAn0nS9iMI9VrcuuAuctQDq8GH7wew
QIqzEa55PWcGnnmeU7dQLKdDqdr8prynKh9QHV6tB3T94PGPbbdST9iTWmoOixT4Wj5rq5naDU/i
YYDsMSxb/vPByoasaU/pkZk8FHOUipwuV8IyO1Q46u1wXhniuqTaQUqnMzXAnH/tUx2OffEAWkdN
XZsRZWcggPpK/A5QWVXDxtN54YyLBshFFcP0AZaljPor2HmC96wr8/j5w9mQdMxRJ2gC3NHFRzmN
cPaxbHOGMmPzuGkgCm/46sWRopnnjbPZYhnN2BtDEXPAFgfEPY6uRBlMNVdPnVjrHjEljWsIq9Uh
Qagof7qhHib8fr9CM9c7whFTHkNubQV9D7W7M0eRLkB9UwZW9rCkAO6bafu1vcgLO2/AQ7Vmp3Nh
i3f8VVwC4YPc9HRGn2GRNGoAR+hBHURVrqp85q4BMgZHziik2l4+u8LHYsCBuReEZ+SeEsVAnL+T
HEii3jBzUq+9HLJMpagD5hX0vcGBejPEVS/7ciDMabpoPH4VFyEDTRgHKw+5ZlHPzPQijkABhiWS
zQeDTqbHnoVMNVXtGgjkXlbB9nVA6oqtTVT4NUt+lP7tbdITweuXpkCVOlQoE/MV29Q29qA3ktNN
O+bPWVB/Ikf8hanRs0kVc629Twa8iRODFV5HcUWKC3kYwHExPEvRZHXnpC5s5GehFoqHDw9xoPcY
IlMkeGMcB66ohcyNZb6QT15RUi2gWqy9PO3/0nRjCXhNtkT7aCooos1cbv25BhcDtf7fimH9+Clh
nXQbVjr3kY3/2hZWwaeWVOAi3CE1LBWeRHBNmN+7/cBzfGDdGIhR6xHM6ezZXZa0vOPWgO+qLLcP
Cqe/uJXwaViSn9NcPNk+QJrN/UqIT2lhc4gZhStCaeLeQtB70T3PLeYP8BpTN0rlbKUcaIT/e/+z
X6tuRlVFFwyHrqH9V3Dh93u0muuWBuKLpXnOUjDexHMY1nlb2X0TyamgM/caCYwGTn5cF0SweR7y
/uhJ6ebCiVMniYetvizCijin/xjBhiAAA9GZzZ5/zYVddJwqLJGR+QOLR8zDFHI5VUmX52z/BPgo
veuy0ccq/Z84jbGOyUCu/K3ugajJtOnBT5DARC6CRvOJ8O6EcSK3iI8MJkdE2Pm09sD5ahxe9JWS
qKm/r61UQx6o6eudd4x5m6B4Kg5jDv8hfrYoHb8PfqQlr7YzZMJYIuNDdbNr6goZZhxpwPZbf36K
pa9dYlBB/MAwy58TMjqrUbq+hbQ9VYKZxq77GVDvtwu5Z42+rNuqLMTngtq6RVfpOjK9qTXIrgQM
8hVl+8WKdKoGaiv9px4zZbrj94tiyUtZqlL854p3gBYNpuS6MZ97K0qROfoooYgSRB1FuqAtHIpG
a9bb/ncXqkMOHHGii4Y1Rn0xYCOE/1k/dm/L4IvxucrYumIBAO+/JbolTQMPDGgxR9L13+SXILnU
Mp9MyGsO+nxbJiQgwtpa/UTD2eaPSKkyev85MAumK4tNwGDt+Kb5YgA42YIfzblVCYZ0GsX/FlKC
DSdxuPliV4KGJS1LtdzOv/mkhDUPCQdnzc6xh1gz31LsjLvoFeOFKDlb08d7MD+PM5Atg1jpZKAc
P3O1L12bgqpvzSPmCnlumdGlYNXRQHAELinCUTZsR7W4IaZTe9vjSV6mLxrJmehzWRVoEGnvE0/S
NgILXcu/6iqK1Jn1lqztmniCDKN9zd2TlcJgZfWHmXr1wiM9Eckn5zXylgWWf/orKYJNpA6r5A7/
8c4GRocqT/Mmzf/vRah4RYWRF+fUg8JuxOxA/IPxTu+10PvrGPL6drquVYDZl/fGaRL3sbxTeTQS
KXp5de6S11boGGPNppAjKPF+rp1H4c6mf+5NGxGBQdRObJux3katxJJcfras8O6v3RTEjrZSow/A
eD+IgJG7jSqt3gQ3cNt2QDL90cb2vp7WV3T1jPiKQypirFNFhy5+Uxkg4ZkliM4lUsk4NmIe4eJn
1Tw/JxwbcLTmP7YdRpaTRIjb/uSPHkA5YTEqvYyy40JpufcTzJqqkKebDlcO/VtyDXmxk+pHWpmR
xxOlk6qqIjYrqI+7436WhCR9pUsU1djydPjbuXCyi85WbzzttuX3cKD1rpTq0v7WomZz+lK7lcyw
p5KA9Net7lEnjQYLOAwtO++nlHZVXy2nmpCNJetQ6Gsz6HcPb78yHluEH72Uc1oGXlDvvc6NMaI2
vyjvUMlsrpchDf/43v16ZlAFK3MngkuVWyCQRwHVSj5cMiR1cVT7EGAyKjN0NnDR++yEy1iJWqbs
AyfagwVT982ewLgGvEKF2XyW+jaP1/n9BEZ77bTBA/6ZCGEub0F9fjH9gGcvsB6mA9ZPHuUldYX/
aYsE6A/jGy5f2GVAWaHE2OE6oOXjLO/Si8p/dqUpYZ1T3m2b/lbvasXn1mTDz79OP1qsRCihJbLo
NkcldmjNxyPbclbnD579erAdkG4S1d1CF3thCqkVvjqkR+wpSvbRJEq4KNcR3tsyceOgBnj22AEE
FM+iXypVFA/NTdfP2lyjgfwSou8+f/yT8VVT99nEMvjclx+aW6gPDP/T4PMe8EpcSt6RpltSEGWm
hJh2mqYj//F07YYBAG2BjV4kQ9jW2sPLzGf+CFEChXbWs8d62Tr7w7Pq0+aEclPhLCfIenBQo4U8
Uwqa1Y4SDNmFnipAzoHeCjHwSlZ4wFmveudpzFlRo1ROlhNRHHgjlz/ImnLkKoJoup7kQwFP5qvN
/jDpAFg8Y0vyoKj3WsFnkrEKauY8azc9dUucIo3YOeKcAm4z0+a57I09kPsk1pJt/WZo1624Jr7B
bkTPXbElOjEzD/+Wgt0Z8D4AtJlbuUVA090CE92lowwS9PAZkaKhWxV1kNDQ2MsnRfWCNnGNgpou
4R/Wb4Y2Dor7W0H8W5JR5mYKDT0FfdY6pDWPlQW6Y1UURrmiWcRbPtjnhiNPFuZQc4RkQ4C9sNua
hmgjM3d9FpLi9XpCdWPvU1yUKC0N2R6nogv9OJ4hiCpA9W8PplG3TlLG4IvJMolZLSpIyYpsxu1E
E0WNtP8EchZdXj3uMuqkezTkK8wsQtrzdY6pJlFi4dTKdT0QVKlVSVubhE6V/BP5rdPkEgSS8ZiW
K8RnGbzWoL9FvsjLMnhlzJB8ZWlUS8ej7/fDjL7zF+L/33K6KnFgKVrKR+iii3wdyH6VEIx6M96+
5IAcCzeRKpeK2D6nPy1SV7XayKeVdecI1gcnmPfi0EktgVME7ub7GZGeFOHaFtYY40JQh+2+7Q7R
jsk4pNi+dyt8QAy5MYA7AnC9q4VbtxYhYxnD7+qIjMZLoKr60I8ZUGeNBTenAVZv7Wb6NaVESDiH
vhRorrWilqwmHbGwLQ7JCB7uoq+Hkz4qZ2yA6Hf1QLPYq3kqbL/L57EDqslZBz7jvdpYj6suIMTJ
6G7TbACAcDv++rQTB4U8Fxu/cELEPQj35yXVpQ3GDUKL/H1J++e5ZzyNYXq7LaGOWd1PSSvRvszi
ApariWD94Q3oM0wsfg3ZvGp6btcG1FowrhyeWUcf9YNfcCNiIF4NwoM5ywE3DEoUxK3YZMSIhT/+
2r6boXHr6Gd7dU/FqMkw4zdKGSNbMdLq0UApCYiNu10BWxjjNNgemKLQ11z+Nyh341ssxCP61LGs
4UwqRgi4hI9G3OCBsdfXIxg9rSvysdLgE+Fnlgdm2EvYHGSuuFF3m2AIHOBaDaO1B2Mp4dzJv29B
mdd3YoXS2IbzOvVhulgOOfc3UKDk3sEs1LCTI5uiGtP9GjGkwznQRtw3CCxsn4pIp79e+YcjuAUF
jcgdjOl27qKfQH18PMf/G5YPJWjG1zO06rG4AlScL0igYtD4bFJ9K5ruE+34QEyW9Qhd/QV6fGLr
OIuCk1aqsNx2jAilF7XYnkImamZuG/xFSlkypqPkky0eyr/dTUaGn9jWobyLaQ+j9+ef3+wIBSNV
crpbylOBw7eGRVRdIkAGQdXuE5ahsbDp6iiZ0Kqpf8ELJBp2U5vRbqWxUwdvv3g3iqdAxoHuL/Xn
xOdKpiggG7WK8ZcYBrZ2XCzF0hIq4nK5v5moKAEqr4S9+RPsDzcnGm6JlUjtgn5eFirWDRxxe1cc
zvbDQsinIne9gC+4J0iJDvHo07hyvMTwt6Q1KlyQRqY4zbqmEIDLNdpcQBW8xXzZMRNBG+xlxb4R
Or93Z9j7Y5nw6XtfAJu8AgSKP/WdKOhfxw8QHTGOhu75XWZVXwnDlpCdRS1YTiD/yo8D6kWHSXok
PVw2n0qpOfRTcAIGVUvbcsdfoBS/fYZ7Nw4BjkHQkxGN1JR1QZtCwIuevkXY/KnsBPyX/jP8KN7c
dCFVkN7dMyPlV+RMxgseo1Cj4+kF4jjJsJ3x8zoOWaOfd5qbcKT9vgHZmkUgbGLcHTpFm5DbJtQ1
E2m5kcDrRHbdhacr+xyZW7Nz2mcsGzxAs6ZuRx9XPjKc/0YNDtftWzvnPfk3D2MdYu8YlhVJlIhj
g1Pp8Quru3PfQVLUE9FaDhtYBGaPEtZVphRfpupCJTkpVJX6g//MUR/N/3geg39omNROsL1FXzDH
f49he35hidC0SIUogyatzKgg3IduvICOmlekZXh2DgCyYppb2473b4Ruoq6KlYhloJt5N7ArRH99
7/IKagH7xE7a7nIPScJw5SHns2H8pwgzNFluqFxtCok+90IAZNNzQVIs85FqkAImxLAA1dwqAbiN
rox9iF4gkS99Dz8Axy2lwj3c5qdPLa8wVzixyMnHE8dgxxPMZxVMGMZILfKJ0P0q9cagUrcJKGsJ
lIBYL/qoSQoOunmDXGjZtLqAxX438AFDE9G/I4uN70pvVp8On5ErR2eLTDZ8gMrzmmyQY/hjIn8O
4y1ks3AW0JodSJOmDYTfPKGijv5eAqpgvOztp15Jr/z0j7uJxFL9NQYttfqiZwz6Xd4qHL4KDsP7
+JZF3I5dEZPV90hbCQZCxzmfdMyV4YQmwQFz/0kqSr6h4FRV3kTKTP1rvNMKIn8HN3SWmG63LAD1
zYETr+eVcwgXprSZH0E7HxCoIIyYgY1wvQSMPJNw0uefDUSRmel3yLmal1Dg1atgFZBqpfKCGAjn
7sFeRR20An8B51IJRAs2S9YmTO+W/IksezG4LS2Anwz5dIgv/mdv9VIRAnEBNfOTYL9uO2jKaIsh
OZVDItxI6WPHAngEoUmaPoDXhbmdpSuTfbmbxlbhgUQYodTx//Ku+c/SdBbPYH9iJTwuSQ6PRBoY
NDcGnyaY8jVNWptbW9W0ACTAfBWeQhw2Sie7YrVf7y6+4+r+EECmKLG5qbDgcLGI7m3bQ9OrNjhG
jq0IEdPy282C8eXwvnXBBor63aTcaSkCUpra8eRpXkQOZPZh+N3z/l/SG4dGgwaFqKZqqxEP7n+j
1U+Xy/8vZQczAYico7byi6024uv4AM25j+l0TQvZZqb3RwrLXcUGoId1MH8w5UY5AI5CU6VYorvI
h5mBRF1cuYJVbdLriHO4DkppSmzZDSrF/XORF/40DBFAXPBZfJL3czLcxy+h19jxjObkrkCQTGfM
quxjlvfVEsKU/aJ2UdJhGNjGZkE78yPxGSSPvXoWvkQ/cYq9xJOffDofXNkOMFZBnZlLco0U60V4
fIVU7MyG7rTNiSuCg3veqeTAZT1z69cg80pouY+NH41VuPf7ESd6zAAH9ML3TubKXUIamD+jKG7c
P6NRVppHzBw8l7cwFO9FrJWOpSTWTcI1M/3U9wZbrNvYszT/NFaJ5AISuXHAD42oOPVSIT3GT2Hg
dlPN2cx+mY3SGsN1pnV3CZPQyp4fU+EkZdQUuAlA4KCxywTIst+h1ZHzLOQhVtXiX4cGGvp/vKtC
XuGaoCaawbj4Kgp4HwmVv2kXU1UiBXkdsRDQJLzgyAI9oBjuC/t8nCCvHE29ngqXqn0eU8ujs7PT
4q6Z+wJJC1n60aMaL2ORIPSyQ7g7gRtp2U4S8h94m5+3p60kocjvvKQb4oh2k8Rjkorw2m0Wt4TX
FJWYUZMQ+xwH03Yqdw6+hserCoEUOv2gT+XSguWjVij/C9AfAbu34zDcLJwX4x/+kDjo83LokyqJ
Ns5y8D7YKzNqNyvLGuDWCwRsH2VJ5gB2rWOlCxt3QViq+l62F7AsAjq+JdnqTIchZOD0nt6EEhJc
/Ld3I3Sk7mjowLEx1bDbEfPPkfbI0T0ExWtGf445znGVdQ8WWeu0Xgl3enksFqWx95MV2SLUl6gr
s7qiTe7E7nBs30HYOKlpUaKABGN8TZ3S/uCjYzcJPE2OfzJBWNk//UVC57p4jab06f/OSQ0zE+V1
4JtyzG7F3xhL0TzZUSb723i4ZsYlZpQgD1/LbTZvDavrVTmhJZfwyiN+QCbXvwf4AHPdfZppSIJd
TQwkOxSqJcrLxFhD3ctADh585Gfoy2z61e5KXI+MyEiTBPHdXcHMsWKaRuZ+ELug29GzKMK0KdaJ
7O9q7CWpOY6MogdFIA4LeBZaIeyEPAbXLRQjQmIn4yTyLMFNQ7//SBxvaXp5bgSX79Q/LbPgShrr
00jMiUoj0aFfg2YGwri4WG35rA5OOF4VcFsvwEQdzWDi2IfWdlao7AlTQpdsBANJaNXu0xwDxiYp
ZpXw2Hsbp3nQRJiSJw4rk4z1yUqPfqrYejnXU0KLmsMTeO7Lgjyrn+pHB4bGcT1W+qxER1Y4rKFn
eyS2esA8Zs/qK2l2H/uLevLIpMQhxKcE3YOGLtG4aT6QkmSMtOISDkXNLucrs4CqzWPY5i7lhgD1
TSh9e0D9/nVzSSUr24EWsTHfYCU7WbJvron1JSRQKWkBuUhDP0W8WwitHWNaEH95zdluBnVwTQvb
cowyHYwsbHXuHtY0PAeb+pljWMO5uzGxEoucSJZMxCsOOLUf//rVRzMUYMvrmf9h40ntG29F+AqJ
RBpuofMTtFO+GKktwoFyfo8Ss/AcdYFKFntrkCDbXio3v73+Dr/WanW9DUnBLzH2lE7mNdinPvOR
jCh4PalwFlQUbb0z2tcmQeL2P/R2VEmMoznjE3Buu0lncmOajBJHeRk3ZxA/ixd9zm00inS8JySy
nNNEjvGfyNTV5gyKBFLeatehZHgt1ZeOHcYZEz4Jl2q66oCq7s6hcJWVk8UMLvS4ImV55pyAShaz
YjLr8Bj+PhF1nqXil++H9/raxLuDy8hHe9vfSdFRy+V1R4Xysi4tOS6QdmsrnL687/GyoDd/ciEX
wzXKWTiK5qZnaqNER1CblPQfVDAcaxwoYJSUABAkcqxD6g3lSABJVePJl4S/Ja5DtHDjs+ahZTxM
e+77cbGzcTKNx1cdnomCosLMwD7bkgFn4NtRcQPofXK4ZPCpzebjiGqDBrbBiXJZlV2rrr+Ol/JG
S93w9DtufW4Q+kGpaxm+i5djke785JCQyRFqK6cqAvDAqDg6hE0mHGIECuELdvyUkMG17ahr8ZZF
Ywi+oK9XkfdqA3PTJA+SXhy9dC/RYUHUKj0OQmhlpeRL2PxaNYTq8YFY5xGBiPAcxcqye+JTj2+m
Li6TeWWFgnI8okXwZt6V+wCIpY7vSC0mAmHg5BrxdKYw2kfPTO0T3o2Cb16jyZ1FGyC8bfuu6FMS
UhTPFkcgVSvKAfW1aMWmSMQ//qJqJMVO5pNK2j7jVhoBGGOGIV5H/Hez9izfkj+pNLM36U34zclZ
UVi9upVDIkwBm6kxghPIWg7NgAMZLYldc5dEAlvqC0Qytw7tgehIu6+rSnbw+k0reJYY/X2pSckn
2umPb9jKUn52RBIa5g/1qcGxDBSqxSwScG80c2sUPShHIP3eabMN4MZYTj7ug2evBJ9i2u5NN2kH
B07sPRhrIDu43k8FJ8L3O7X0nXZVobO9V61NxFiNkdnsz35c3fAypLeEs1cUHTFD+u/+sAinKh7W
iVGEnTLZi9ICW5kDuZuIs+kL7ZhSBOwVl1Ws7D72H0HtEWItaIqRcDa8VgTLt7CEZACF9xhxe3F7
F1Dh8c+Tz50GUAyovEJfC6VyWOu0+Nl76LGSEWit3tUJhTlSfOsFXiTbqe+80sD0T90QMH9H85ht
WTVeq9QzOlqCln9nepGDFbbWlbucFXVwcOpQAX5hXqmmLwoKCW2cIniNrmbKeHZWngZaNiHjb+CA
ij5FVx1JmEXpHOdeGrK9qzxPATs22Vvhp5wd8LGtcU8YCUCqaUw0fMYJhHDBAnVJ3y5P+jFzneb0
eII6+zh+9mwadvQdCUYUn6St0Wf9hHcZqr8ea3krUAxA9f4MuUHR6eP1VZzDXDx+lkzNVZ62B/KP
P1VGb6BzIU5UgMUpsQ3pns320ttE3OXTyeGlycICTeDyHxmv6w315N7FSpgsP9kTYzWwKhg50Nug
J2dSe7c2N0aGFfOq06QK/Uz7oZXvXPPj91EC5LXZzRo8XgsHdLIvXSAM9qAXM1ls0827I7NZH8fX
mKFcfHfc2znqKUvkjZiJK0L10NjKxivM9TFOOdw6h9QLRfXYZFLxOnRm5CmmWX8hCMSYdhpKWNer
uKVSAMUfYBc+NHshMbsgDReyxUvdb/G7dCG/7uNNvN06L88+L0r6IKOG3TER6QiG6U05jhZUcfaz
7TX2Fcgg+m0I0tvcgv084P7UtJiecjB7q0VQu6siSwtwHF8qD80iwew0IahYV0LdFu2hF498ozCH
D86Eb7MOrtqL7kdUD1EbX4tbvLGS2aLX3X6zsAvCa7O2xGNFaq6ysBWgbK19XLFW8PQF7Js2OsSn
YATe9nq+fZAH20EjK9m9xt10xWotYuPP8V7lEDJ17G430/kYnklGuexW5YsTW0NBzAal7Q/XkWQp
EXuRGkI8dBG4JFZiCZIyq1GbfRNqtdDUttvyKnViiyyi1FPVUm5kT/221VMtcLaXzgqUVcPjHPsH
s/9DfvOTNeWur6Q5IuULdcgjTdFRv5LAZ2VE3+PBe9PW4E6y0Oyq32tnE/TDrl7MOgf6TC23V2nJ
JOyfDxrOCVO9oZO8Gd5g/lwdJ7LvQdoNYg7KlkzwqaOj0GF6JJW8y0Jt4ifXLtxu+9+Np1LRje2p
VHm4gHBgcI2H6wbvPRku/G77k+/CacK5YmuI5kIFPIeU0pMfpuW+INBLfqxESka25jPycsKsiMMC
SOaSCy8sBT4hAWYxqjh5CR3CCOJOLP5StkAV+JuFCsKJKK5hRZM1AxaPulBeDbIZxYXJN6dOZUYB
4W7xd6eo0jj9BioUxJ8wuCcC+ABdCHo693cMqIVL+5p5vSMcCQfket0lJ2PQpdH9Is8yTiuEE+5h
0kSuX9+D+WLcmpVVvsN+cGV9ESgQrhx2vCYZJOMRIzxxZqd7UkDMQ7t2H8LkwrrKAQKvbIQJ2eQQ
gaOUWKsb0f9OGRKxSeH0dj3CSvocmYW35XrX/HCwFhLhGkXjD1EDEhD71MHNi22M95ekXdRVDfom
FfDeweZS06Pfaac+BD5JzRXP7L2DQXaN+ZYHmeZut+758gqm4lc2vYubeIKtG5YgIw4w2Qe6pWVO
hO8N8CiugjFYg/BURZmBcKaGFgNVqKKeLt6Pr0YjUipXcSCqhOHYqvQTSncHkqeoQWEx7Yj0GDhg
Y7AsIdmoKWUIVELw52PPx8jfc9dVLF+jYkKyF7oWIQDYvwpCdanu208xc7/jMK5TicEGQW9LHzzR
n6Lu0ibjrNCHwlgW5p7Jkz5YBIzNB6Uo3vJAnaBs9UyyV97/dQucjjsWvZOPYBWXDnfzPgL/kfvd
K3+EK34oWzBH2CBj1dotNbwMqLs8YdEdCnsy7Qt3eD1OcbH4setH6yJjMEOXO8eb56KhkD9FJtoU
z9/zbTW0i3ig2vQZdIB/CVNGTCmKvP4xxfUaKJHzfU2Us3Y9dTBgYmjZowy+cQg+vWIHMDOxqDRX
qlCAhwlBsaYUzxuUvMpYyw8HfdtGfz50eF02BbZURpo23N71GIFih0XTCCAYwlvdviBSrXpaGBOL
vq9BIAXkAr24hzJizxbooW2Ro1wu5exxFBxxGR7D2tmnW7+tz0P2WxgxpRMJ7SPxBkVVYoHqYPmM
FN/iLj6OzU0OQV69R5d/XDm7jG9XlZKsGo+8uTdo5pUWZGGjoDYweMkJiAbxQlquTdiNZ+xRaG7F
8k7rYjsAG7bPWasokWiBQx3B/e066xqlsPBVDzscfMrHT3JmRTKEEc/EYOggwaVsncsSSs+tl5d7
Ij34IdiBA7pziJ5iuR5D6Wt1WnpLQp30+YvjwO1EcULlCNF9ToKATubCETeYoKaHmGwJZsuPedya
Tj/MFxCXOvYEWBCcuE+LjhvQKpSEyRy3RfAUxh7TxE2m3AZ/nkPEA3Yhd29CQmICprWE/dOBYmKm
m9s2WjpBiEYIWy7V0jZ6qBon1aO7W6XQ0wJPwfWAkIvx6kNPKVDWcqRJ36TXWERZlepdQ5sSjoDA
9adwZb/v5xB/5/JEVKQcWxinSaRcRF480VCNhY6XGdykyuUwExi45LGRU+CPpk/sNVSH3w0FmPdg
/Nv8hKNlJ8HpIo+lHGh4Q2Cpsw6yJtdcw/1ml8LFm7pCUjD/i5uzBugTbETMf6ovokn7Ms2ObesY
bskCqto0/F/FHSbV0ZAULHpirNG8Lp4hbIj/0nJo+DLSroG9abWmYrrG6Fm/k6pPPF0jMq4tIUMm
rkAo+Hy32sm7SeXrHokcMDqTl5TgGSQHxg1nw90axf2jg3ZrtOAzIkQNGFQiR6OWx0xV0rHDOE9x
uB4I4Fg1rMHe/Q28Is2ml1qemUP+6Cf7Yz0VU9ocbOafuD88UNbESth4DHNSr337bmC59W72jI6z
KvDapWyO3Z/U3RwfjqLZV05FTuov7f8U9OD4yk1IF8FKUrnpTeZ+SGuIa6RweeQDD289vE27AvMa
UN2xBRCEuz/yrEYxQSOYHDqqg/svlk6JNNOgnuAELHFDdmgzQiGtV6O+DIiNyM/uO53AMJuwRd4k
VeFpBXkhgDu7E9lICpmrgmNXePY+G/lL8ueypuHxNwlM5CuQ+mEd7uxxheRkCK1WB+0cJ/739vjr
UyLKDYlk5P1AAJLZRgVWShXJgjtfK1uz30YqAqLGpE8zVnzh75JTWrYtzBmgltqQ3KicjbPaOP5R
0GVN/kpt0GpqNcA7iS96T84nuubX7PHdj3VceeVTPOxk1EOQjHWrhW3KvteLryR6MGFiR1h24upk
/1mxI59psqoOaWQxnuFS1Z5oXw5CnqIQv/jSsSh3HpNTuSiXoNgKG5tItnITeWeZfWmrKtZ8UXmg
Dva6DQuJarAQ6pegtCHWHhoLGSKnWIN/qMxucDg4auOa6YgZwvWthmSur7e6QpNnxXZzt5zJB1P6
+P5fWqUTcOZVvzSy+9qZYlpTJpXh2mYXHK4GlBIgNmK73Ul6+kiTljabNj1jzGXnPm+atSr/GGT4
udW/x3ntZv73sI25sYzStd/KERw84Tre/ALleKsfuaBGnIkT4790C3iELuZ1si+TNKvafnx/FdyQ
iXwi4JCkXZwZsF28q4svx7sMuCAcorvqtU+ezP80pL3fwhxR1/HWfmydeWNzu/wECbSfBkBQoMLH
RAnFlIEb+en21yYfBJn29sldBCdgSOwE9Ct/2Fqi4i/4CgVBLsg7w36LSecSf8ilRXNvs+vkhZiv
l5DTRPA9kZf8O01viNilQvGKawyMKqcnTiq6hvtVdPK1b0Dq7jKFuhXSMQxgl6aXbScn9zzrMgOZ
mn+StI3S026Va1hm8G/nFmzNitHQzzTnntlVJ5nKi4iFG2oTspd4tsD7qp0G5N/qwfjSLRAxojoD
lGpuD4LW1pVAktwS33XdnxByBaaq00M+da2i0DnfEvcTsHYzOo8MA624nZLVfuhQWNvxTjxOmnGs
XWxmf8UCq7AQHtXJUZzsDq5uP7gZ0QDW/vxvXp6I7ElrmS+LxwoS6WSfzCZULW2nUQhoY1R+5lb4
3WjguVISP9EnwT2eYfa0vzB8Vj+PBaZsZgi9T838Q4OP3fYGn1AI9vtxX4E+k4AxLC+LMPDT+H+6
3LELQERJC+cb1DecSM1zE7f+DiKgj/Ukb7460rYHZZ5EVmOtGGW1N8VZTjhHDCGoV/eWhCln0yP3
/Mro8glihnXlr4wUfTZpMhR9tKD92D5+puNlyVAQ4gLs3uflzDPso1VWsI+Mh09Dp6TOKdjX45h+
hkCMScZGlgCzDh1JxPlGrcVGDaRW5GojCzo8m3VuTtl+LQg/oLErSwoWnVLA/Lqv9LeWfciKu74Y
XFT5cKzNH+s2PXgmmJle80MJ8euknm2LgSAa6IhmIDCh45ssywMv6CeAbO38OgQ8oeq7F6UDvQn2
qV2XnLfKbnNvKFB1rDw9dCNAwHfyIXL4TfO2Dmp1ZqfqWAYTF+JTxPm48u0JBHNgC4OJNdaBish/
/jjjGg0wh4dXqHeYdSiJnm3CkpGfxAv+pnIYRq5VrKU1LqTNKvk4XBJj06xSb92a8dsoXUofDTgl
Bwpybf7aVSYohoD5zcVNC9vPupVOuIM6zwJkCYsFKxtuKNXYNA8w5bUjyK+Vy05rCD/Wztm9k4lJ
MDdlsaDkj6pqDBP/MLKoF0wilNhUG3QLQqju46CYtQdh3loz1byr3tCmKgFNLQXv6E+l446jzTgP
frnA8JihmQwU+CyD6H6V3KX38ar+q3B12Qvf7FqoxZI7vaI6krJOoCMUjV1zHYt837jEuPlYMPiq
rdm5N5nKfQWbWn0qveNVHWBuUViLMdAyTpWvvyIMz9Yi6YjG0U5wAJWSxy1TW9RPAEH6198/hQ5h
Gy1/FW+H1yyN6mxMlZ6Kn6izRlNGrR/FqJITxAXpQSgxXbrlFAE/lKoeG2jWLuPvrYJByonganrq
AkN7rdHxofeU0wszshhoCXjAoYGLJZzOmpxHSD8Gteq+XUZY/XgjxH5lWPy8sD4zN97SfYLMkkhF
sx5Zw96nN7Lf/Ji547c4duOBj5D8588VAYQY7o1zMnFoXvp/CBAfLY3S6m5GchJ7/fV5Fzhnn4Rx
Esl7fRkmN+SdaVZP2M2MAk8xlxJn73EL6PuP913hQ+2qI143fG+bv4X33Ar+NRPDlu4FXih96tr2
f+Ju9xvRjUv+1koIvEYtNT2icTDA2ukuo9OX6RF3aaj5cT97VnVTIAKbG5/OPjnHVnjyr0GcTY/u
8xSW9HibVSZ4wUeTk8x7zQDQOyFUKEYalp9fS20GjZF3u9419mUOc6XZskc/gaJKk+k1MmnedR3I
hPnyCxRPTjs5Hl6SmzCZl1kBQS69m+B+ZZWdbVbu69wV56kLOC1Vf4qFE0/9p7UZaP1992typslY
uuy1TJHm/8QmrdnYKHsxtrvUwvueOFa0rul5cjlhFZJ2z0GCEsYKpAjz2watTwcCl2wUm2rOTZnY
uVCl3hRAskdeDO5I9gyv+fut6FYeoELgMe0Pu3JqRMmS5FocAcDTti5pkU+dfsFu4dBuJaLGdXZn
l81pM+sVaVGdrtDtdGXPOO8hY2SPGEgRewzI293xTvqhZ/t17bEx2Fcbyq2CLhQOxnNXm8Fg5A+5
l49qB5X3+qmaZJ2NFSKTFP6sWm2f8TxZSz0S0DNVezuc7OlowHclMgZQ9NR2GBKpJuQ9TFu5Cjzl
DpqIrJocrtA6t89LuYdHNswIy8h8NOuH40s0MWWOgd1lsg24cKiumT2HESvZgdfyaT5+VqQ9fCPw
uIFIMppBFIYsBYNuh/tRSmqZIyGyoXXLWmt/dcPlXH2XZ8rR9QrzwKe4SXFaKWaayQaijkkrentl
jMiaEudlpiWz83tQqxmcGcxAw1deI4pfYdLEa1CpVd9jKUcPfgyDmp79Bf9iwl7TyCGbUchETPef
PffBVcIhN4oOyhKIymUopOcMPg24+/0lOB1Zhz0mzd7l7/x4YD1lqJPh2CmbyzJJpMhHcHowAAVn
h/Os2Sgspv+Kfx8MWcSZ1lZctYPADDs/RSPT5eJVfn+XWWmxODO+wiRjRbC1ZHh++hTSofJ4whUY
MPUJo2ay4QgrkieFZua5TEu+dmU2kmyitQaiadPksxr++8p6apHuBUt+bU9LF3rDfSEm6hgyxzB+
9VVH0RF2DWFU2FIpJ5gurrwjk/9ujQueydw5Gn2Nz3m17/F66IThAZDWQbX2TPoEigP6IU1azc7b
tx3WVHtdKEDWFMG3KqtcjXUEKO7YuB46KPtrDR3Oqgq0pKv3V4d4bbFNCmWRJ6FSXCjlfUitsbHQ
7YEUHQ0QHDlfECj/9b7t9wRWvd5+qPw+vTHIF2flq855wI5pgDR6deIZtrI/+dvCN4lwX9J43sL5
kCd23VoA17PrMUEFmNWBj6wes/1+1ekrCg7VjfRyAHnxCfDyUF6sr1d91Rur8VUlPYu8NHU+Cole
Fizsv8H4nIxTxeSM92FE3eSaZPcWTIl8hvFyHMKMKRaXwsG7MD/Cvxw+E5XPCFy7iMRdydeJD2W9
1YM8ria+KXpDaga1sFiuH7kQCoeMIkjjmcl3O8EEnMFb+BxC0umLomcsAdlgsaJV8gjyG4ZB/MXA
cCSavPH411uLby4ZxKzdn+FOlgFtk6ohXPqwMvPocR/CW9Htxyk8ooviJnF9Cbw5Swex0tyuUlMk
ykL7Mf3DMTA6uvgzvtnHttmsBKLUjkbh0iUBLLVRhaww0cAFeDgTqFzTFjC+ycJj2Gg/7spo05/z
dPMd3WcGyDKtyjw4tdssUxUtI8/PixwrYqloudDy9yCyndhvGA2yct8zcrB+gGT8ow3fHEBDDjtj
xibMIwzVzUXotI9e4AeoJyH+TQbZolvQ+TZCQf/e6YJNNobVOIAHP5Bmwy8SG31uJLsOIZoGYLaf
64n+O7lSv557PXW/24kvxjY45VzpizTodltKyQAWNZ9Bu7cPc5f/wjZXnSAHTrIO5TPDUvqLPu51
O+WJnxE9C5LkON64MDkOocs9BkElcJU+S/RdGrKwspIL4tXolaVkWJzPf8rTcN3wJQwybHpt/2Me
951rVRdVz5k3SB81Vp5mWl8aqhdvPxgKpUjAX12wcY8+lWVtzr65YyhZglunBGJ42PDT9laTU4OH
BeEqQPbOhNVYtTLUiyXTXmLotasigEPvB7wvZKN2FCOhbXnUoJvK4QhzRJwltBELa0s++zi1Sgp4
egzdvgcOfnpvtxNqgcAbImb5qfsGfVs2EpgF+64n0Zmlf/M7kCHx+qwk8B3sZh7ook1kGZQRtHrn
aLadz25xwZxuCdnqUeXsQJgIZaspGh9Drg8GJlzID6h5hi0cWhhK+uwwSxNJDBo+0O2bs+sWRa5t
5jKZR0xkCM92Z+zQrE9s4UFB4fkyXdwNwZ2/h4Vsx8ygSrrjbFpSCdX6MmTadrCuIlumPOZinOlm
o9hsI3fLYw0GWDDLa7VXr9h692/lo+p5/9oW6K1ZOcPRD3KJCpTnfE/dRwbivvQrH4mBp6O/HjIE
mDxfGWZtlncLv5PWcYLgeLyzKMpQLCp76Thj7HTsfQi3FHRh6kg732MHfqqdzRJQnGLty34VOue0
y4XcwQOr7utY3NFHS2UJoIz5ovQTmAslIMdVHNWJ6YP9kLWG72Q0olpWMV2nc/WO6ILcQIxNQ3e4
0UuNuw6wYvgxRPEBNbzAvETtoaa9aot5vCfLs0WZ6Zsk40n3Ooov5zLoEcihwb35b+/y3w/2TD7N
w2uo9vG551Hd90tM6e48gVbjDT3PZfec03vCocR6WDRkk0UW1byGuvO+SBRYq65XlzTOUWtbEw/h
TJeq62T6fkJddDFLIlkAPlA6Fuu97Yr9Tz7lYrsD8FX4SvnnaMBJ6YGRp0s6QF8TOxpHsOZ7mQMX
9GPPz0VjkpHl/lIANVfRDA/+JH4XcOCBwPV0PvHKNh5QR+rRwvN2zwEC1OrG0ASYRjQX081YgBWp
ev+qIZSJ7M4Eh4/dWhVp646ZjTntXTCMOn3qgF79pAa1M821LIwp3KxO1mvPjo/iQtAXnOOUfIM7
lXZPIJ3gte/Z4z3I6FSBNkdlxJ5zrj+t0qso5QpsZWhtg9K/sMbQBKiQgbM+LEsgST/G06+mQwUI
MJCJ69nj/HADHkKonSsVupZSH8MHucOVbC7MRVrVGbExDLblGQX+cKZBkC7yFkNwTzkG8+wFdJZp
7ASxAz15eUdDJTouVJy6rLFyqLWDW29xGxlGOt7qJZ5d7DRxjKcBqNKT4IXJLg7LSgg04l3Gt6Wr
c4mc1bAbq2+uneuicO94ycEBkLM5wdqec2Ibl+49AZelSAF41IV2lEkWXY0MbzfMSLSD6M3UfvlG
oSLyL2cre1acB6MeISfu+hkjqef0pafUOdlkKc1R6Z2bhv9/LfERIqq1+hbHfvpRCBV4yNOOaMvB
q0MrD91KuTVcCEPj6uLUj9A1WPTEmunv5roFY0raCM7JkLKqUF0cwpEeGXfJ5lSeElDdleV5Y52H
GgMY3F4n1y98Iv7pyKtu2VR4Dj1FxJ1V0/gM4Q0Ce/ldzjbh4GZfCxdItw91teWUr5fLdofe1V0v
iFe/NKCy39Ue0daSj0n3R/CZ1+bKqyDpBZnHr+XEx6m+Pnn4+PRQkH22SUm9Azd+X5UushKx7NhP
ozDwULhKIFIHUY8JEHdECQIJl1qnpeTSKW32DBJ6b/1l/FgehpbJSidnAU3NRxj304/sS4DTxJr5
IVtyl/+XyV6boxCpKzy/AvEM0rv7ZklTMYxanVrcf47nerWd3AEeCMXkfPSvPp440z+Z027hv0S9
ghMxN0GmnQfzdPoPJk+SikxWjC24+f+B9uBB8brskDymyLrDgTcAXJ+xaUeN1prNrAEs3+D4oVcx
JSyMKxbMFJPsbMyP3UOqih3Dd2db6ARptPIOxE+JOcU2eYE5Eh0WFYgZFrowLJ8CBLoj9O2wo/WA
NmzYdtARPry5CzrbYySyj2jqzEMe2/EcSBrhN+zPbLxgEAuLVM25PBvvEGHq2qWYPhVOiauYRQrr
S/CYhk1Xoc8/o1s1d8pw30KhhmtAH8leOkS4UsFq1Abu5CePzS8kHQQiOmwAvRoXrPCi8VhId6TX
3klqhn0nOh8nBbmLLprRSmcXjLVQHIJEj2r79Z1NLJpgog/kYcyTSP+MpF83HKvfH8ysB8RpTXZ+
Pd2fEJM/S7lJ/ojJB9gmsylzdsrd88gCI6E71Kn/++H9JufPLGo+tV+H7e7n2CMGa/nqOiqZR2QA
qxuLSxwiDMi+HVlMxYmuxu2FX2zjuP8gqi6QPSfae4cqM3fGplXTU0IpDsq9kBxXi8u1gxfGfG9+
l66bf1/EOukkauBinmc57SHZpToUjMJHuQa+k5G8dq1O56x/DvDlSfbUIKWFzuyop1MzO0bEvjj3
tAv72FoGEXUMziqKQC1SOPLo5jlAWuwvpPvnvTatDK+NTP37vuKhfhuw4gNVz7FlYMvfKK/zhruU
FfcB7HrF+d77NYQEpAcGL1aIZBBFlzTAzUvHfW3/RTiQd2C0227ixDZrbCM1V4zBEw/haCFkPkrG
yJzloQQXKQIJWu7UfQYGf7d8WkMbd1yMSsBdGVrh66Q48eD2KLNBA6CfJynBmUl4w2Zx8oWKPigo
/XJTTHFBfQYeNeiWWYaq6JJJVjtOb2e5tyKkG5NDSRLhwmbB7TD4vgef9MgrZN1K8vZ+fQGhzAdP
b4uaAktLH7chOx0SEXNdr3HiI9xZNK3ysLZjSB8ZSXZ5u03YT+oBgOSIxESt0iT7VRixtkfC4LE/
H9xV7O2NcFdBu1Xp8b12xFuWTOyOIn/F0Gz1GcGZRZ7BhQJ6Q0DwEvnWY+cTouBYx8Marha65LDZ
MVz/ZF08jeW/c0xMBZjHkwrkK/OqLimLn2Pz5E/y9MXoOXSHyWt3trPJ2DvpRtY13/gQtsx/v6uZ
cZQWkYLmAWtojGKB1WhJIJEZV60h6K2GXsF/ilBZcxNIIOOR6Vd2vIzsxtLLny9gKKzg8aHWOYt1
cHmvUlRNOOwi9YYVDlL6zXu0xCvlv8WzwakyvfOt41nPDNH6TeSgnTCT3irhnoyEDdQ5CrGIVEtW
Es4q/HmLWVjUufEbMVpBLtJISI7Z0EXiE3WgWGGBScOv3iq132Z3LsCHVDFppxssBQ9hGhVB6ZgH
Fpi/BAUiT5EMrVnTJvasGXiTtB9ImH2hUQFQhaXOLl/E559a3kM6+BDRnePSGPVlPEqZitpKCK10
//YeXBqXCzSr0fL/wSKSUd+jKSFw4bIAzwLTXpzNAblJ5ui2dwZ9p6TyEVeqrJQXJCdfEmbBY6BR
We9JWs3wi0FbInUYEuup51ZnlUmKGeQRUqOVxzRtuPMUtiu7U4t1jpq7jTGgIMFjHsYVnIw7Ks/1
UKY+cB7P5aFz6aVR7+jWld+WDsZmTqqeITC1iBY/7T1WcvGj2H5xJy3sFgVHbA3gIfKDdUG9Rf0U
3eY3JUmGSJGCGAY0BPhdc5ikZV06PoOErUGKrkHOjj4kBWxf2tIgHySc7WH9jlQao9owmRWOOHfc
3RHZlXMfXdCTl2aq9Qqfbu/updNW/S3FQcMy/EZpMPUvJ6kPi763T+wetZEnC5ht9Vv25WKdt1Zo
OBM8KvIRybg7cWCMw7lUI1ANAzvuh9FNm8vTd6EOc16hNK6z44YjFgPyjKJxQilrko1HGsgk7HrT
D1bdMoxAvgau0WViHWO2k+GFuxO5GMTg8H3o7EAqEKkDSpqA34EFZ2RSmf8c9soR1CVnohOGI2My
LfXBP6yRIbkpJWURPX+rZVs0QtTGSWy7z4gcm+LR6FGkW4hje2fUf6x8Fa7T166+ZSZgzivsCiT5
1A0gLw/1k+WJchHozWBqAcJPSQWOxw0tJs1Qer09XJpQxZaB3ERMpndnLjclFw7wBciJSoZDTC4r
ErJW0BzO7J8HBy0JJSupJn9+Hys228Grsd1M/jLErjVpjTS160jQp00RNosqxYGjmSYOVZeLR1XB
lF+t6wLMrbnW+rqHNtx0yZISSuNYjYe6qoUG+up21EPBImooTysmeeeBBK39xL7h5+Fnhp/q22Qy
spFjsDV5ouZ0Np/2hSQhWV3dsWPtac+FCBM38l5EYRLqCg6bNZDJxqdgqbxiIwaL9XWv/LQRZ/lK
3pJRQSISOfR9LSep+hd4dVP2MYCPJiYaOtWHmXqjGXrnF2hFpNgmTSddfnxSUH2mZUTbiLsPf65y
4yNS+Aq4vVWPF6+8DRzeL1D82/pp5/UPscHhWcn90C6dI22LwY4qFbTWevfrrraTu6/GAmIZ+XYa
TIxzsu7B6p3/c3QpBz4VDOiryXpsTO1vhEO3KlqdU478tn7FlidhFoHAInheA8+yBuxaJNOCmng/
xPxCDm1oDVs08W+/J8ghj22oB6izLcw0/W+zWAsf2lGuLB4RXp12p9tFx0AXcCkJ8Y4CbVQJA6xx
yEOlrZ+8mNJLvhI1mfAHt/gWwKiB0K/DpuoTttuUWLyO8dn67TkYNpNAtYIMrc2eGpk9JqcJlrxP
CrJss98/zrrRJJdQxO831hxr6uWSevSPza4xo4XeKuByrANklllJxp7C0evJHk/tK61kBdQicYE2
WSFIvGyjZnKn0A9Vtk/jc21OJpnj9OhZYJ/g/YjIiAIxMkRkfH19KfLNZkv/oHbUEUdAW9bXmVhH
w9lBML8gd61QcQsJ8F5VPjCMqnSVriOmYI4D2r6hzKl67casZaG82iK1kPNrk+A+27KEFNrIic90
UzHM4t9nUBnV/P9d2bAgVX8KSDFbtyaSwd0gkcP8FzKlYq5JUwZGKrGLNuwUbRle7FYfP/LXDEyJ
7hP6bfrhq3UB15Xq0d00BNJME8FxeFnjFgNmgROAu5SG6TkcPZQmvWe+vy59FKwDp8UE26r4wF7a
HJxEdReCuuBv13HUOsswT/5/kUu/AH8tCYdwLBO99RH1JnoddUTT64BuebkxIS+2UnwkS+g8n1am
bn5kfoT/JN0yUCoHeJ9UwlYhRQ1yVFqHaR47984GD5zVuMuAky0tiCsbLTPIych6aTfOA+2ezrex
X4W3R03kXV2r9lY13NWS/Yex5Yuc1lbdFaan7kbU3rZREyvsSStblKJb7uFieG7vMdXomWyK4kSv
IuBlgtoQVsw0vtdp+6KLdIvqcrTsFCwQdpH2jvVDgktFB61vR/OmF1dp9Yne5tENKyNgNQkR0/hF
/WLn1X+owtBRUUJfX4F/xE343sYgU2aAvtDxuu7COxf82+0hPoZkpc+gE0urgqEXdDbufwV2fdpB
aaV/gFSjYJ19wRS3wHre3Yq6+DWqp0naY2lmUFT98othL3/xAJpU51Ox+iM+bngakae7ofGor8GA
hjCPJJQZH1ZIJo4BxcAbnbZP0+PGv+lPn2qp0dQzpXdRxPoqIsCTHcZbPKVJ/y2KZBRa+wwSSEJ+
FYTvI27bTanSyj483IG7fqo4dbQVyy92McfnF0syORjrltIb4GrT8eUXHCUo78oOqO5v3Be7ezAr
j8XRTagh4Qz5FyLkY6X9aHl5SSbT62o+HcsgEggwmt1/EvRDcBUq9uw10EPT+3RAeHeYFxCZjuyL
Sm8pqaPb7//GV///9X5fq6nVba/VytEdkMcnHN84LAZN1IqqbhskVx2ONYKiElEVbH263VhLUaMX
hSc6xC++E+ujxUIMNSoKeNm+CePhRffhYapWOSq7ooeKjx5EIjpB2vCIOI+YbUBGla4sDqYPziqp
3iREcRbPBGBOvG7imvNFrO8ux2wfROi5mUaTuWyIjXFEuryBDEABYvEfQVFDT6vXDUQcl2hqBf45
CZEmZFPuzDoSc76RSni2gP80oBpD40AK2HUlOHUfKrQ3b1+2VC9b6XXGJ2keurluNk2xLgLMEbuN
zn1vGglJFs7ibBia2wbYLw/+12FUtOBoyLi3yAcY+rMEktLCkmo9PrzjYi0U2ycefSlodCUIjwR2
AGkA/YAHaG/DQVQkJ30MV545AyhB8roDx8PusjXMMN022HxUm1KN2Kn5KuzsA/sZ5T/Mf1BS9Gux
c6bzG0zDntKQXO/B9KF2OyCAjaevNZZLgE9d0nFrbO5t2G2aImKpzk85b9Bf3FBG8nT5etwij1nf
2704+Kr1b0ZKjj8SKaV1CBo0Zd0zosMAc23AO43H9SvrJ+ETniyN7HzNVf8eovE5Gbbo3zAVlsq/
Oc2+GQXI8VjE9CaXj9UdI2CR+akB6+6AzUhmmHiM5hADZwhDIAlYKx3m2/Oihz8P4N6iITSPU5sW
mPKshSvESeppW44au9Ng0azugpsBWrjZsy2DDiut1jzPrJAvFQ0IW7aLrCDI/5yeQfcc4txYJoMC
9X1A3nDYob6ZHUgNoVkih6C+TKpqyXZg3bGjZpGXvkaDKTuLraGGwpQzLfSyJykmwEZkG2FtwMl0
KpMXmWqSwii/+ObJUCLx4wNWhUHm+8RZe+BLR8ndKf7xNggmR8v2zj2QgggYFrvmN5vc3Bmm3JPx
NF4ViQ5gIERb+Fy6W3JC+YWVNbLH+Uuyn06wID+4gPnkNF5ytWIlqII4H6kB8RcU/12wl0XNG7OG
NDs6PVAVZZlisC6fRkDgtamK/xKtuGp7aAcwEE98bqg4L6wF3YtwBPRYqGJyEL2zYu4M7rfDIpcr
AascDTJP4sdi1c2ZQzZBu+g8xllkvpX6IibVwob9lhalet08zTHe1ca43SZpuottyD3r99hjIayv
ZqTxHkNh6PjyAD5yCPJ6XS/74LG2cJavGfaHaCvZYcVoY6vQwlgrhTaaF+a883J6WWWm4wmEpxsl
+buawN9/LcODzari01M5EjVVLv3Ll+wjtKMf8l3J4CBn9RT0Th/yEkzMosvtKY1AugRhPW66BmWR
JvGfDV5/528riN8zjFsqsBasE7GDQgumD3ONIkKZGOday6OhfFX2XIhLAy3f29Qsay3Pf3XJIQBu
qvmDwEoYFKgNwyHRpY6XSm2NUJFrpr0243W1iEJ1AXUmVLl7Ao2NhBe/zHnCj5FZjEmMmWme9zc6
4NhtrNHq4XN5cXyK9P33xGxMQ1fAm8V8Pd0g9Y+yiDSZgTNDMI1tmpMlomddp1KjGepLCxjtCPTA
4nhML0fjQhFoavPkzKI78MJZn8feKFsCiAOzyoQHikM0RIi909JsJ8vvPaJYr9LbIa9/U+pMxxXX
cKZpxiSOv554Vuw9THd+La9yyqwiYqn894y30AtnkWzD96/k8NV9X73w/LWPxM7OGWrogTo0xT8W
bVJhLcDbvNhj9ZYNJTYBlm1OFROPPCSSPuN+8A2kfor7xQYvFrqPwZB4ZZGXG8JRUU7dV7rvMwf+
X1NdRg/g5uhV81YbB9ys0XXA2TMPr8I3vf8cxzf6qNnuV1NybuMUyg3ltlH4thNlTIS8eKlVeH5O
VTvqOqJtnZFISrZEd8lW22i4MiYcwny16aIpTPKY3X0lE+fQTrPxKvtwmWjlQO2RG+VqHDWkhaZ7
NIRutGro0WzIcSVP0OdMwsHOdMfrMXCzMywDGErTM6+12FI8t18Dz1InTGDqW5dxS/rXtnFoScJN
peaHI1sUsNzqtIxQBhhAMJifC9rzqjUce1FgASlwjQ/wy+uSVpNKz6h3moEALyuGDQcGxcQx61gs
mnh2Fsxdluj0DoIpyaOQJcGI608vcis1YVP1Va4iS16DhLBsgTMM96ev/7eR4wAxgDW/K9zUR25z
4kxzEI5VMUfWAytGNCvG3gxKV9fNVzVsn9ZRoQMGoi16jhMlqqX5lI3XS59Z/i9r2lYMC1yh4C7V
v0VIRMzRsdcLUL5PP0nNQbpBSKp2QT9MRvRLd2daPyhxz6RBLCWsnpmWtie8PgtPFki7f3I3cD6E
GQgLnsWRd8CAFRRXBGwGnQ+o8GqJFGgh2Ip4xCrUMA0PdBO0fhPqQmmFuvnWHDisNQMO/f2Tk3cz
kTC7SjR4uqju/0cERqtKeT0N3yu2nHV7bstjF+xBuOYoOf9QEbRGaVJk4c4VUqVJUQTdQs7Hcn40
a5swfUC91M2ZeK96n48X/z36Ifei85TmT2TiYUuvWVr1btKpxx192sZag8FOfT07mMf2yGM8Dldi
eKVzAlk5kULLRn1cXJ0+PPm2w76AIBHv65f1RAFOiu101lanMIPbsbR5j2unrWzZxwJddG4NSLj9
i8FqoCxjRfwZF18F1w1+zQNi7v5w9jxSufYavo2iDp8zU9KDkF70SNmZRlwUOwifGjO/xfa0ZoTJ
i8I4mGKUiBQMei2Rlx14gaTyiEPeh3kqA+5B3JG8TyqTdWRtPhFKmal37O7tdji9PdHB6mIm1V7n
+H9J6IuGZ9Ir58Aw+ImVyVQEhrhS4bkCVW3sCfwdUAT809dM4q+J+OlXJ/bx1J6DxSfYdo5nSkZO
06KBoc0yn6t6s+D4peAr8YsIxjoNyVEYprAUoTt9odYCMq8l1raG6HOJG/i6vzs6kRqXwx+OeIQp
t9IcUF2eJLY2bUBYaoKHCnTYSJuXCEJlqeoabed6SU5D+b9d5C9iu+UJ5TD5JmywUrQlRRiQbbyB
DqcV6/Ph+NZKNfd9NU7PGFZjZv7QbgxigmVsNeCPzFRFnnRvxJLacvRRirt0sVzN4UO78e6yBkdj
Y3kUj2r5p2ce1LXuWxnzfkMY4JS/ymQuG5WnHWemFk3pjAievHzEkDuri23itN09ZH89Iu2uZbd0
AnHjddf0XCDjcdBwgD+Lk+lHM7vYp6h/AXIlp7gPkaAjz2dWahVu08UzTG3eh8u08pKtjlYyHMEM
HzuRkWxZq+OBicoxc1a2HW/s/g5cXI3r5Bz1fmXDbOrQHmuICxLdkpTAtd/xEUGz5is6Up9xC9Qv
YOkrfOXhE7FRCA/sFgguqAMB14D3BThAChk9+U70myJ9GSvpLycUASfFnsrYdyABfVdutfzhDD2q
dDo1/54A45ZSqkvMqKRM7rGv1Pt7fW5K/JalgiUkjBt9cSV42AsbQjI9CBMVAAouqB8tNisPIWG/
CPz9d3Z7p/X6muRtVC7BzwuUDw26ozHujyrRK/Eufnhouc6F7ukFwnwVpsSRyVXa4CSZKQ2KDnmP
X2fHsh+DXERs/DCllVGdt2MCFapOikgHOqn1kTctgmXx3PnMhbeVvFDq1pN6PixDErRawGuwV/vO
xDbdlLxQX7Ng1OY9Tw3R8VXnviMleR9AwIvMHKzNlcMpykDitrGjwbiaApJkSanVXuaMAwLgUsVs
yX8JWKXHEzc5IgBNe31Fh0AHsmBXMEtS7mSVHWWYYLxshmJzqFPtoec1rjLkKZKrIAEbfg96Qt6S
1yjJOSxJpd/qfl9qyIDnaI206sqDvJJ4w16KzQTqeSSjQdpDw73VIK2tpr08faKUimJEnJh/d1/e
m42sDflKGX3SCnqRYkudwUfZEHUlZ8r/vgaPNGCPS4/Rd3tQ15K5oLxVTnOIH6AY1Y7vcZuri0+T
YUIEsQr7Slf4zjrZmI1EFKCmPqXb8rfd+eWT/kFg2oojlicatmZiPqXtlenI67wXcMPt1q7bBktn
32c4RgfkUmXGzXoP8igMeaJDPUznrfSqPyGmGYAzF/M5uUYtqW+Qa2q6LniHPnIIrtaGIwkxD8kS
dQvzxLimt9eFcK3F3TUqG0YIJr2+MB1d6/0+yWtSw6nUOCaBiE/WQn/bwMsXEklVeZnnDh8iTSRC
MVdnLSwuA77MYZE7F3IuhHWKprIDnHKi7xFFwCtgy+UUqdsuYbPjARDMR54qQeR7N++4WR7+ZjUz
TCUA+6Gv0KWaNZiyrS5tD429DqddGC4IwePWSBdBXfAcAiSSGUqphk4AVb1ccAnXaJKkYKZuxe8i
Om+bmnK10GeSwHeUqXWKvfpOsDrM+Dytw8XrFKcPhm1JZC1QR/RNIzRgggyfJcxM79OmLXE0a6Nt
XJ1NMI2BMYI2lzx4TjYK6JwsCrNM3A6gG6rwpSkIbBsHlJgZelLnIZGwl9muHgo4K8DfcsoOnV0V
nKc4NcH0wUug3l4fBUWXAUzN/omCrN808+pcEH/fHDWpI4vOvJwgvtloeOBqpTKj32D+RJC+X7ID
uPjHdTZMC8wokPh0YU70Pb2v6JBM3YskjUH0vVZqLZvfgNfZq8fd5uHrjoV2eQMP8GHAbZ1EFMtL
6TxjOvJweF3lAbnO7njLVBgNXcWI5jbyTZe0jg292byS0bPNAJmW4vN/Je8B6RGnIbYCLhXXSj9F
UkVsmi4ziIet9p8yiLTDjk2j8Hh67VIurAc5Jmkf3ngyX/1vRRVIz/RiUmxomBcLDZ/FUu7j6HdL
vtIA5/DGVAFJm/zRYTEFElkp+Z1YIN/sXZJFe8GSnHb/dghOYwq2SFULJ7hoV3xHYHO2BsQNrxOs
+Z6wsmlZ5LPlPlJo8v6yWQOHmQGu97NZLBC+VYvVQftBR85QBEzuqSJ2qnSiijpFb0fLQr4Xcoav
j5sKy2L9yv6UyAXRSKvr0wcShuU07JFVb0SMq6ItgJxfN5FrWy4u/U/nB/7UZe3rI70zC0u4fWdn
G8DmoP2kWRQByjrwXc3VpDanJWCfjSUx7N6oXzVXvc0oJvexIPxjQ2RdSmVu3zvhFmRqLt5W1aQO
JBxzzqvMvW6PnRzCMpZGT7fAswRPbFjEfTm67NweMfZW1IJNgaPsaYNFkGFNTWPrSrNZg9Sy+Oa7
I+7uVI6B/HdRbb2x4AknqqNAUCkBhFx+wsbOZTLjDbImsVBQf5oz8IEH9kxJS9JiMaj1bJXrhc5L
ypFuwgywcTPP+qSr7oYKVmAy0uBUu0cLVjVeowPwSBo+9IfpH9eOfIb4kvwJUOc7bxMQfSv6Zzkg
ot/pZaB6G0gIKlgDfA+pRqy/d5MU91tY3er8x/D27ajTdXXp7CXi5Ep/GjzDxUOwYw9ONurTiLam
qkTe3nUyLitUyzEilF/FzrcbgroFjJuPBYT/jhwBrYHcgWNDUbahMLn/4sZVWT6vx99lKNqq8LtN
QerFWxDK8TrFAWJIcTwH7K5RA4f2cy+ccaeN6ZrVKVgHdWlkN+JhM+tgndGxoSwfFkVXGtswgyXj
pdwrbNyteQ/thUf45Cl0qN2KFX4PK9fabBByJ9GsHZnyPvxHa3Fr2sUSEAlUcMBfrv8Qs+FjvZf0
5U2T6ZJla97ZSbkpWpnJ0x81LQ3JkVaLQalBfoqu/F3ljGW9pXtggizZX8EfVWDaTo9ELVZy/7iN
2CxHvCvYf0OTs29ZXyo57pGoK78edZZZhbh0JNfBznDiYOPgLnwrfWZq9i1CjHe/QzPq8GP1w6Yn
eTmjHnpmSxYktd2y6cre4GBR+aAILjnUVO5FbvbN696wOiEueWQ+1MRnzXf0lrCDHJ8IVJa66CMa
7SCRlZ0PdQdBqRvJEcDSauI8ZXh4u9VYUgzQAKrzYe+zaV4AmZTUhB5PF8+cOwDnlQxdUck1G7JH
DpXhk9wcZmz6icZfQdxUYlS2E4TdA7or4DYffSj1T/lMqfCHU2HTpS3wqVe/KQCgmWmBXANHV5XF
eN7wMMUQ1QUBDGzKXDKjPXKmZhnMkP/Cv2yhtZ0xce5FjiYlsMkFwC9Wv995NoFMozGwFMnyKU/J
M2Q1QAlyXwT64kc0RV208tl2PuJhylN67AC2q/1KJWPakmg4Hnr61tCiE6LCt8ioOBM9UyvSx61v
kDRXAAm6jCan0t03ldlmjGYc0guaS58EQmvJDxdE9XVI8FalMOXeJ6e7nLyjOHiWGgVjxDnwt3cB
yfFXSu1kqHBecN8jRDrMGKhiEBH3TUelSJE+APtNEPWwta4m9DjEqzRpCD/3ARdECCk+DSef380o
rtGDDis1fdYZO8LGS7g2HQ+Figgan5mqVSBITQveKEkoyb7+n4tyX7NZcT3iZV2z/5xMfv66qvq2
WQbVzvLT5BZxcsVKY0FDwGw0fvprg8hNk2WcjCwfO0vcUj6f0F6ZCis3BLYqMopCoHjf3zAfDtRV
6ERdCnVMpGX/RXQwH/mApKSyY0z+40A5VP+jioMcOde/jlzd7TVvSKwzNrBWiKPAju7R0VcVcxS+
QpeLwTAcFxpGySf0o7ad8sXkCO/JcIE++1dj1hjS0/BGjNKsQ3bXt1j7e0C3CzyLorKgVKTre7Mu
4A3Xm5Cgd5FlSd54iAdumms80JLo1SEff/fsDyj58SQvRJTurhJZ1H8DQeyVWnz79T+78lLepfLe
C9gEtOsPUKnxIJ2h94Au/4XxOleL3EbzpI2LL59THAeIt/R5jxFBT/OSEM72riS8c6wCWvOMydHQ
4/9Tuzv1di3aosTAT5iwEM/jiBT784LqWSux7dGVhGXsnzsqPQO+CvnWHOD9x8HOLlR8YYeKGopk
UAPBl7xhsWbBV2qN8R9g82nvSuOQ5tGWUx/G7q/HBUxqx//juruJs5E3XJEVT6ZfFG6YwSHvFqR4
eHGitENAJor51oHDq8tTPiIuOalhV7zIcORWe+edmtFvZ1urLEqI/uPbEQmwqnmoolksRBTXuTux
I1vnaAylTjv7nmM7tHZCJTCbvlql+twrNK37pkwUaD2CMW8mbVQyvflca0jM5liNjFOwN3IH+nVW
Oourqvhx4bFAhkO+yGyZa58IePPuaO5tL3srIQHSHt/9hFedT+8yeju5r1HzRgaJCa0ybC8nWt8a
ylnN+EEnFL2EXA8NnW2b3g1HHsPkREOq6q3c3lDxh6P1gC7L4A9SQ/3sCbHJNs/MILhUsK02DDij
LtFzrJmG7reOCHuVgdxYOP8Qv42OjS8K91ZlptYea62HFrXS5/qi5lqot2Vzu7kbXFEpgePxwnkK
SuBgddEJRtHo6Ux14sawqIKGGch87gE2VyPLIjWoYVrJ7v/BC5xjHA5YpgexH6FqZ+Wxdcr6vlGO
6Q7Cvp5QeB69vXrX0xRxdW9H4q6lSmjXKgH8aTj2k1ZbI3y+IRmP54PdIxO+8BrFq0HbAuRTTnEk
EhAu57zJcn2A1UwAyZ1D01Me3hQl7BMC5qr1tuo+5/0gjLiXddsdGiLcTunOsbhWuEkKI1YA69eE
HxKXAYniKfOtKEa6p+3oOQNn0R+0e9UanhinceWjYy2ishjxBVIfxk6459M1mh9xA8NZG7dRoftH
L1rRh5isOYp7r2zrQ6GMpLMM3wQktQeOuRO6UrwV378JuKPVxDyWqZNA/zvtzr8YMzzbzs/+08ny
Lt+jm2hwqlRooHv2cSk6l3H6rZtAn5qsyl0D6uQsZaTvxry4f9nWvUT30rvA3a9cCScvdJ0Pdxk0
XWQkb5hMBkoz+foBDzZ66P2xMjm6P8Djv+ES5g+b4BtHVeKAt2wPzQm0VdCOi5zHGcTOxDiksf7W
K5HUV3U15paSdNLr9O6dqAxKGPIHGzz6Fs9sHJkf2WPdvVTAaO/sQ9ii5n9MATzELPvoV4KoMpzB
GK2WXJO+rXvOI6KOUSp0DLv+8dr/V4efrFXZ+NnG2ypF1ftlSBOAHSJYKxK7KuRq8JMvf6E+UkSp
uqSz76Simqqb5xZKpGFZNhxWmGfWa4bkPzkYtLCNjZo/siMwb/HCg9BVtA87SIK9PWFolOjOAGFL
fSX4R2KNgnLUyNiP0B80TLW+VEOyPLc40A/jOTrau8gmaiAatcAOzbMqD7CZQSx3pC9sex9Fhiwq
HMbxAzFgBgAzg2QI6h1lIwbusyKNoZVi8vHPZ6EDt2vdzPKNsjEfM6jCONSUh5dM+esxTKBWTEed
E4nxlEhKC63YrJYV2f7LUfKwlSe+WSwcYNUpRAvZfzKO2vHkc5p7hDQb1/IYDrXUODSXsD0cnjpv
qk3OeI5ay/ZSgVSkBCbTafkNS8Q9kf7qnWZSI7IfpbebEG3z4sPltIKB7ijgy8wq8UsC3ouDlIhd
YCEOmGycETs7UNoeof8YmNlWI7HcIIGfTDApQdVIahNMbT5wTOjgYvALBW580/FB/gtIrup9Zsak
BMAddC07wISME3QnsoAVtDUjwAcsd+iY/WFWWSG9L7SZff5BaGe4f0mp8r/lq9ck9ZlhD2xogSnl
if3ouwYWXl+sBKaMRwyXDSXPqoA9WWQIq9xi4j9aqsHmI9qmf321pYVdnYEqyiSZVXxxUpXtOJ/w
rlRcU/5or2RY8N0iI/f1AAE4P/AZ4sJYBeWCfCONWH+G8wjQpal+bKrOD916yU7SEx9lwM8lX81Y
n0i8mzzOrCyptckZIuxwCi8cbkOAZ+vwNSG1Wm84YS/EmyCfr6BPKmZivtPTMy2ueIRRnc+HD+5M
RFf16X3WZ0rz6MemOp8RtAjWHv9x7SBoMrJEe6ZwE5KibJR8Nqa0CoQFJtg5NlwvA5/owyuFFrHE
8lWEsgxf/B9qnEGNPC1DxJCcf7L2YlWg80hzLDi/bknIj+1e1kxQ4pDUjY3BCVYjkrWRHqcfaPUI
HyaKhdwTup1EHefOwpgIVhSIDfyLZGpo57IOvdXZlGAcCauKz9LTwWhgg5ZUKalNqA1HKdLGFjRk
ZvNz0Wi+WMOAiisW0BTOi1OUc8HI2BXZhy0cToPjEVqL3cm9+Gde4qISFDHh19CS1ASqSDzoHgHg
rVbSnxNGGzoUGXA2rfkWqu9+IPymjRzlH9GctjFdhQz5PLTCAhvEg8KDDyE8+OHjL5fJ5thmf6zG
AA4wpsn/FkAtgx1Z2kOw9rUh3Pr34C41R4M4bjtpas1zN5zUMtkdCwhMnNXzwWG+1QwbqF8Dlzi9
X3MvMJXhAkZ+WfCqrUwgezy/EH7UO6RWUkOq73gbhZcAiQ/y4hGvrLd+GqJncbVkvVxEwAdhhQHy
PMmXCiWfZ1v6stoHB0HQ5GpnJc1ExfuW/rlGTG33Mo44nZAQ067wkxlRpQIcyPXVQwqHn+8edyJv
JMn/T4KUpiaWiPE6pXgKkZVtwEkXkI4GqosBQ1oEBZCQsL0MWeimkeToW130AjTLypUgagKSFiia
BNacUXqqLsLh5eZl5aqK2ZRBpWJSi/pwW5lelz4aXCuo0XD1NPTSavO7BS7jRgiDNoHeUw7wA1oL
D6Jwr0/DrnhxBwtsfXHrk5bHX5IX/iHo+3p/GC2nyPpCEiwwSKtRkOYCP12dV96vRnUqrbBTMu76
j5q8Vg/vyXrFiH/m8LRAM4ZciXhop68aBw16VFrU0P9FujnhslGVZ/cstjID/h82A4CUbsjeMazk
9r5le/ZOJEEBcRLX4cbmY8HtEaUhB9IzILlg4XUDckXNqfU4GGqXNvAHVNrzM+y86UVWLKVrfaSi
fFiOn9lBiBPompMAuWQPWaQRYVJf72En041sCbgoD2X1SIyTvKcoMsbWnLcXq1Dwq6tS/k5eHP5D
wWy8sQ0a+grKdJaVVyyP54/1XU29TINvIbB6bDfWediDKFDIE/st6V4t23qV3WwDaGXMLYC0zs1U
Nn7JNidbDFIiPi3t4dukgGGvDzT/n9tWiSY2dttDOKngWYxOAZVHoMB+9+Mj/j+YrULbyJ1KQNvh
WKn3++FEBEoiP1SP9rscyw/a9ZkpBWXCurPyJma5oItD1Jb7iUX8MPTPDmNmiE1/PmmoTC46imhu
gI5CYxdJkKCArOpDJX8m4MH+m4iijNdOTxJkI+q5jGYiyMB8VKAtTRK3ikEBWQLSao6Tcp+KPa4p
mGgD/v+D+7NnM3HpaYMCAHW4+Ajv6DipyiC0qpwCVly9KGRRjbkBOEKTUHIAcnZaPfL1xEc9UW97
X0vPS+zYcKSd6uiAq5iukLqxwBONBCad8hwv94D21V1nE4xDmgaQdP8PlWYW0iAPkAbDhvr6CGEr
eUWKax/1dh9pT7M8vAI/EgNBLt/s8MBLlpc+lwDM3aPdFLDl/s4plcPMwyvvq8xJmk0jBWxqN6bZ
qQxFdJl3OrNRPwV2t6L64rj/jQsaQbRjn5+AF56O0nn7HDl3lW8ASnM1v/eLpQGXZvhVL0uM9q62
oFUYY8k3MbObtyVoCFzGRN64YQ0UPwZ7yfJVSrCaIJNimmR/8jHd26y5blWnLERcjfWR4XmdcI6q
Mok5DPw0neIwIP8hn0iF+MjikL1yb5mMy1bD5re2GOf1Hn5czskW/4M6PEaNpomF6UASGalrgWHL
ftoDjf85HSKVeLY0+QVcoWVHLj9PMXMC32EgPZ1xTUXvY83LX4HT/Azwxg9cCYJUpIiHAGyIMfK/
Fptg2kOtv44L1fCfbGqSYp/cVT9evEoON9jR1Ual30IvxmXby1cqskZBKfveEWfAUXlWxG78n2z5
JJbQY8Ap3IL3B4V3CW8/dGAawEwFB3g0ysr97sHCSWQC7WJW/QLne6KZGdd8vrMK/OHeDC+0eE9/
86YnTI2TfmggeG9Z8682UmN+avB1UUDJ06lPqMTUA9FaQlprEH0P0KLtkxsxl7lqJZIfQIpmw9r0
PgbZAB5VwCLx+el7aCptVeh3R/AQ5Cv+KifpYZJ8fYGPjwlW9UGEf+TW3vm1NKTjRMccSPO9VuK8
/ySOf1lx787Pqqoa7qixiwsSgdMK0CyrHlX482gingJqa+3dzrCC+YEPq5UFGBxuuCCqjuCSbIuN
pkSbGryOLiKoPBLgXszvnRsTX8Z6yaZX9Nu3hLS5/wo5S5uknjNEmex9IbUxp69795eeDvVQYi5r
eKeBD2qxPhgwKY7sj1RjyH/zdYDtp/tZqAhV5dy3gfVT5WqXf95zUV7ZuEYLNWOCmwh4VLqPMSgT
MOcWhxs1GGNmbJEyyjjmOBbNHWs1HOYaSX4G1tVGcoCvnL/3iVE+wDrKSNjOlZAyPdWP7vek3eIf
v7SaeNzo8vVJFUPb5sPqXz46h46UrbppSZTMSxMny1uiaPvvg8cOqc239pwfceddcX1/z9EDJync
BxiNdvl01jmsODsRhlutzbRw+/6Tn07UlelWeqju1sEyWYdrFC4OAuicWMlehit0XUruzgzN/Hng
qB/I8Auw4lww1rLxtc2PXCwGxPWF8SjXNNEnsg/bP63dSr2twg0NqMg8bKIa8n6sUxMNk3NehZ3n
nRYvIJ+sVMLIkAVUhQFyAfFW4+YKHjpoOfb4MC5DrUdDefZVz5SsdGJn6/Nd9wETZpZvuBDCv9Wz
VLxo5fGyKXhuT56QD0ELJaspK6iXZGSU1reCSB4CSwBLWoqeKj/spepZJJxRw4Xn/AbTfD1gGUxw
xbygVcm5bjrlqz/05MP/XWzytqGlu1WGk0UzN2ZuGExNdgVpvxGpl9/dKzLBdmgxH7LWlPOwFYz1
vAhd/fPRnxC5kbAtmhx5a2Vx45ZKiSN3fA4WxYdLnOE/QeM3FQ9C5kFEtOuF7NY2iiK53F6SK8x5
37R9s3VzZ2TzbBarawGerNRv2/uGvec9FGcSAEur+RNEwuf0i4d11XskINIwbMTwPHVDjJhD1bXi
VdZ6Oexib/Pzqln6ZJrFpBBa7vI10FiiPqlYSHQ+rijRaMcMv7J7iRKCc8sXimgJe327qG3Dh1xM
vGce8/SpKLFsTKKi+lFVkLmM+c0qKryc3fk8LoF2g+MWqiGSE65gRaoHhdj3gN1QkI7CZqwIpjYH
hIDzFm0dHhTgtscYApEU/F7oGho0MR1/jAvb59tz/ZZ23SJDWb5weaQZHnsAWs4esNMFDeJXzreo
u8r48oar0Ct4D/5iSDIjDqXiZ57jzsABnT32xv3hJvg1V+r3g9nyv14y6l0vnwtgShfTkQf0RoQ2
RsgwEcvBzEJpEwnUzowTZmBW2RHDrGrgG+joktUkoq2u03/Nm9AZ1Kqt0N0JwQu1Cg44XhX7g+jZ
NzB6kibMGNHL/83N1iwHt0Bj5c85OwLHLyICqCnNrg5B3ZNR7ZO21Oxw9mbKJ3iRUqx05omz1Ydw
HIvso9wGeFpduSomRDyHPWiiST7lwdq/Yd1DPFal8nPVSPXrHcxq+YpFPV0hYNQBk2EkYtPpdZle
fIuID5U9XU5KwbBz5x1Vmqw3f7AmmKKt43YNLicsfF+j7Mi0qLOuK6gnYobB0+I56s6fhA+r0HX1
kejVoEbteAwd595JEWpnLJ0P8aQ3xS69WZ8rbL1Ud3tDQeW0JRBhEnzprGze8Z/F2AJsdOrr08+O
UAI9jZJ05JKLKdwu0af3Kf5ql4BLlk3qvxp4AyOCjrnfeBn0UYqjt/TVMLS1O/jkxQeSO0LQoOkh
q36vWoPjX2/HIddtVjaZoNgUmgk4GjHxk/7IBAqZRF/dIQwyHefX5LiQoIJ7yfw4a+muqAUjIyF+
5hSiJ6CtACY3Pt1VLpXm2z8xmoSAKYMcfJF0al8cjOngBrEQYTg50F99yGaGP/kEyM3ecMo3Guqp
5W7BHawI/R3AA0awtNLUlR57ghZNcPKSXwWuiAwSGWtbjhCQxs8D3spwgi3itJB3yJGh6iaqqpQQ
UQJlzxmBJZppnmugmbepQRNr9+YOMGlX8x1OTNvI8oxWy1oh/Ulkd7CZesgJpJNH0WdW/9UhjQWo
O8BRbX/abuR7a+KNfCmC3m2UBzq1HRcNNRy+QAjWg7kPdZ+q3WB6LqF766VfbiCh9xQyYQigoDM+
oqfm597clenYpztmyMDC3Xwp5XKIRz+4mq/QVH+VKS3MYYKsvgQO7gOlQkYv0jK7lNAvfvegI6n1
dmlkujJKiLAT0fr1gUNg+WAia25249PqzIHnqlsmJGfPcNukxZxTkDhaXvKMTWOT7TlJk84lkFJL
xtc40ELDCOWICYCspTTf7TrtGT1t1Z6769D+cWKZwOuBjz05m2QxsxZ5F2FWDNBB28aaCwRz80dq
y6PbGpFy5V3YQXDtgL2UG62qNVLdd1iCa7R5FgV2+Z+kuBNNlhGkx0uAGfUEqw1135F3Aek8hVFS
rutb3H+gKJrOgxLEUif6b1Xj2UsZUD6f8pdjkFNCIQmqPn50So8GhnoTZqLERAbOkdD9RUnXSDaE
ePPxhlcj/oZOMCAgwCjqPBQ3j0HjJHppdZVfZsDmZO3jBdunETdScfdODra5oL0TbXs7nQqPQse/
1MHj1U0mcpKkuW7d/zPMJROOCNZMtVyxvga4ZZUPfOFmrZ6TdmDoByeD7knpU1GTVcxCXnMRCcQf
RUN13PmMEXaVne2vsJD8aC1lu8fsju6USRe2YwjDjZn7SHCePWi7qfohrUs6SMDhvOzqdAHOExHx
/Bv8MImGVtKZkkkmdGTc+uZrINibyWdX3EfkcDoYmLmxoI/wNLN25GiJFkI369TBaKOrr/Xy/4cM
mvwKz5MD0zaiKyJo0e1Dn29G56ZFjcobJU2KfvWoqNthrf6awZGkUbfwVl25c+Zq24WaT6hPR78L
doiSMh5/Xs20QiAcpwVdVuROZbfZ4HaASj0mB0vrYQUIZZj7S9qy+BG92U4gA47MoNgi6Lz5QXQv
WZdfKvrgYgWvpNwhZm7OJKFWlWXpgM3xbKrrRt8jWNwDMT+Uz9+daSJNl3dyr7m44ntx72VCQlGk
yRWiNvyFJ8PupquIO5LQrvGCWYd6ayYr5qeLHoTNsmsWTJH7bdofJzhphpiS6KuVRsukfxEcpHBP
hGjxJ1qTi+rbTx7bBbAba7VLuxpGet0bY9Uuj2MbRk1lHvKd2dNJlyRny60yA7kuljzstV2z3OXG
Up0oE/b5yofHxTez1IbaY5ARo8E2tg2hTgajJtLCCNXmnNfXcWajc6Yc333m1hDwmbyGZOFGxrlO
1jZYP1fOqFuipw8nC3PRLmWkJNoyqxTVUxsR5ffpF3rEr1FjsU/boop0msZyUaVFn6WXkjkpPuW3
LQ4oWMEpSPEYlYIU0IRvB8NkrhrZP8kmdQuMvnfeHx1nD8OQcRtC0/yD9J2MPS+kT5bQExqlBLGh
04hxBqYQMPtz9sJmpGs8i39H0kcZloTe18Xe5Gyj6a0FBeerxmuk/Z2l15K+8DERXEjzUzA6q93K
AdkjwUSxPQCFpZ3g90iF85Lci292VZTG1Zl2ofN3bINic2D0iRRSK6nVM97Fj1SsCvppqYKKi5Sn
B9C278esSuPWb658Qqhsoo/iN4f2yYjWTR63yhtfbi9VFEZRGuDiAGukkZtjs4e09XPnHpXf/GNj
ATyVWqNU4DhzpMeKvXFvmT5aTDXAsuUYy6W3QIkcltUqNAkouSBwJnuSD+VOtOmAXIT7Iv11XRxF
stk6FQEBVSuGPUG3GQIkMIco9wwJ3dNBujwqwODpdwy/K+jXudVO20VIElXHUBIxNhokUeglDnt6
VuiciPJP7M6Zq4leVo5+qoZsHfZ/MBUHrYSO36VOHsJHR4kG1XuA96LJP7SFfqaa0KFuyzkD2vrT
QGxbU6tmeMs5nVXNk89YE10Js7i81Uf+SDomZVycS0JUV1fTzjJX9Lm2AZzuB1v62e3VycMRz9Ab
Fwtyzdov5qlF8Qdv3Z9WTkcJxS0Y8bnlth9s8F9YU13RNPsPBzrDPXKAYaBXoy/uOe12Fn3oorj1
sz0pp+QzqPNRqV/TPaGmtafxkFv6v27L2aFEXcsxsfngqm6tLiw44HhDlr9WoIedCLp71sGWk1JU
8P6/jzwb3nO3CUOwCfeldhsIRHj5QI6SQ4/Up7HCDDr9/WXfJK3WiDwuBF3lPO2UZvAG3Vv0dbC2
QCLudkf84D7rHv1ykMtJLJJWTabPTM/00srhgY9uPG7wZ2/IuijIA99WmFHvYVV1zTAUTn6f2UNj
rzPdVYTsGotSB3Z1yOlX8Gxwah/XhvM06mdHrmtIOY1TzJBptpiHSQ1vY5DOlT5lGYvpxHgA+t4K
AZuR2vVsJoKYAiYVF7Xuwx4f1BMk9+dEqNVxogc1tN3sy24PNQcy5pkuGNqGoFk6rBc6Ko70VQ1a
tisY783S7maJ6b2/ojX8ErpZ3r6B3ucSw+OrPL3+/qycQOMjepTR+Z/MWhjA+SxjWl8mPaHXOBeQ
O5LEZERYV30J5FKC9aJ6TF0ziXycO4CWRd6YyhuFSfoc+1ssPuhgGrfyDlwvznqU2l0zZYltKDo3
y5meS763B5FUFIwdGJTE0GBwGqpBQyhiV7rzWb5f7ve9UZveYM3IHr8uBM5GVvOwHZFi6tsEsusi
q7hDBNo93HLQnZT7YkHy3xvGixEC/HWU0MJ91golzfIri5JFJr9SAVepSrWQaz5B2kk6i7FBiaC4
sZvy4kM2FynuIQeMpcOVSEbByCsJnQ615LCbbwLlEXzDm2i0jSjSm8Egq7DeqoRkzohYFSdOqOxg
9G4PeqFp12evjuulOlPVIZV9VJiP13Jz4zsGK+LmuL+F9uyJAxXDdj2nXATEoQme0Qyw2HlkNAW4
t7BMCc45aFyTmkB3Nkuj9czOUK8AFppd0R22ypLmdtGFnUVBO2uf4aAribl+Ndp8pE6hx81pLpUb
Jl4Z3MjAGcWK0z+n3aEHwoJSHI9KrfKJlKWIxL3y7R3bzn7tMwbdju4a/r9HRjpZZPvyK0+gmu3P
Yo/otYVJShjXs2h2p+Sv7aaitGfEI+nqUVBWjvzebiGVOPEpAVO6P0kv2j1TlSPtEeWzI+Jji8e5
NSpZfQK7HF6t6IhTqlJFzzLOsPxyka64/zxwJnRfcPuPHjpoiR8UnA+5z4K9L3ew7XtNMB2AYSFk
D5s+7rC9fYnhB3ZAVs+w7oOgHJlCVV+80T+zb3q33C3R9pAmHFgBxlSUldroB3sVh/MzGEkHMcJo
+immnEf4EyOVQy0PTYdmz8SI/R3/Fb5p/mdDo6jPfrSWa1pHQAKpGyAgk8uPD/xCmqyZQViXck2F
VC7Mp0NbbwhmYExZ/NBEbBgeMwm4eFmiUOt0JiNqUJb+SsAqWeDFCM1jh3qChHJpkNnesGeyyArM
vqjngbzMkbhjCMU6Fw3pMFdikXWBpiTRyKUYT+7jWl6amq7R+XRrDNE6Yj7qVPkceOmWoOx4UorJ
e+rdsKOX3RZrejtEuMPIh0dtIqkW0UFzHknxZZ1eZlufOvbLkWM8mJYax8M8uO+kIgaknIvswCDg
FGbd5ThRF55V7By3vcaP8omqAlqJ+T8FbCEjzUZTmbpzV1aHkxnWkOeBfBWfI9KM86BFB12nKhye
FgjWD9oIM6jSv0Jdo58j985uKCt/rfo6q3zmuxk541kvoZUBuXKuqGcCloF10dJ+fLOs+rT7eJOT
9YC+Ids9PHqxtaRxrxYxytRsw3iKWJYrjS275JnyetHXvlSXCzuJ/qexSrenF0ANqEitks9qfrIB
sMbG0+sd5RxTsqyeKKPfTEf8pzrYbYw/wZn4I3Tpc9tcjGDuiGPfAdbQpvpqoxbuEvWJ7YvIZ3Gm
1rOFeydef6ynBsIsD6+JyVcDIWm6c4L2zWUwFwjkOUhZpwdfef0gEXbcdMUCmIsPcfvcfSQvzs5B
XblukJrGruWGexyMdU7JCtrA2YeMhc8Qh6mEEt+7rA5qM5cYETTfB1hcwLUObItwam03CooCXkxb
1y+UJBzijTwrpmY4WhoJ7GEIiGgVMTklZT6Yw5qTdJG+1i1t5xR2NhprwkaVER4BVFUulnQbuQLV
mmbrabU9qpQqeoYRqe5FiIXUYr6uPia6/UBBmk9dwKMnNZx/sHhhQJyrarq020qEBQkf8Kcu82Io
b5yTpLVckpIPdXRgxQ3+YpkSPpKoqgHTwpww/xYBzPMXAFxuIdQSznu7Jp/hCFaL/c/l9oWwYnIB
AIJdzQciFzeYhsNrHBni0gawJkld+GmQxj0vhFY9UZK1qml+GXX0PuIFwoyEC63cAjCamvd8YhIj
a7D6EzA92iQ75uZFXp1TWZdz4WDGrghQ5ToVr2nlI3k/Sk/kYMmzhSLRfnDIE9ndiVWT47DDtxVO
NoOxW6IRc/pq4wp96zqklGAsdNm0+4glSdgq3GkVt3g474Uvd3+GFx1Bb270IRYqLlwgkSk8vqUY
XtMz4DLiXtVTGXp0FaODkSDnKsDizD3esYnJ66CmMNrZQl4CdL7l1bKl2WAyhVKy/5T3rd279t+g
AcBrBrjMnua7mt4kBjgDkNVkjiIxzh0rVQ6ktP/xLJm7z37i9oKGiZz5yV9APUe72JwSId6AWtpu
BWrQFUv6tMS+Y5gqzAq5DPzSk1Wz8mBFX/G++kIoIxBbxPu14GjI/i3XzJh7ZHqMsOT8l3rBLADn
NqaeGUxAgFHGR6KUcsTZvJF1eEYcSgzGTEv9LE6FIi8TwsvsO01qhQmrb85UR38brm9EAY7naAJY
14Xman8H863VT78VMqK+FDu3xHfrZZ39y7dpRS2LNzx+LXmJjsZbRYxxTn1zoUfCyCPJWVhFSKkq
2RFltq/7l6z5tl8uf80MT5F9KN5KA6heJmJo4Pi0KkIJZf0QhffPyIttOyuxcJ5MLeypGx+LVTFb
pNyTKCncWMDrdP5PpolPx4RAfAU2RBOXi4iL/f4zGw6TrafCTUCRqCI3q4Vj6GKLkotOlAcQguvd
hpezqu6FE1TAXhCYJwx0p+Z/NmsDiH+Z4nQyI8/slZrILZza86zyPfO9Yw1gvW24RlyDnS1N6rhW
uUUlEFsMnDDiICNE2Ca+R8njYoMsTiTt0VpY9q09KLj4Zl+GI++C/QGZozCk9hm4hiNGsnDRHG+S
N9aVSIZJMPltuUkTDO7B3+dLgaUNT602wfj+PBB6c+AXMO2qB/0i4OzxJCBFaZAaotkNp5naD6ay
ghfRquxzUO8Z2KDLqLtwrcTR7LZ0cszvQ0SKrq8le2RBRE0UIWdYrNbYa8M/yy2g/PfqTV3DZMs7
rVUUKI+UEugsCr5bTymwhLoQ9vHL5llpLtM+yT5jwYvEr8dsLm4H+rokzQm//jzQQ1AFyqNRUBwz
wN8PumVxMMdxaR742XDcoq2cUBdFmGN28inP3CXBZ/PrmwyiqO1kamHZ8VLD8cMwW65Ad0aQk4Ef
UBnSDrVE7VrKO7B6CgBB3ADBDnDkEWpj4oVns0B5AC6gOJKl0AV7irjs8YP8wR45hqAk6NnMYmbZ
ksJ7+UH+Dla8v4Z72nSoGBwJqs3WlT3ZUMeaTjwMfKYueRqf4uOphK3iP9lWfxxABDEj3te9f0T8
EjhwvayNxsWcvfnjCwBgfw2CS+Zo2T8KnbdEtGl1P14wDTZbQWNs0A20P/PhI4hWNfwhVe0eodTl
joeadEtoxQVSH9MrdXzmLtbUsbkADhZN0eneFD5W5titokplos5epRhB66jRCO654bxXZaQbawFE
MGXLek3+ZqWhqyaRNUOW5qPxJ+gwiOfD6TJhu590SL5faqOMA0QwCDYnWj1wWO2lTyA8+9m/9jt7
Bz94W/UtI3eL423JouDZC2ZXafOsL88Fw30OxI74qEcUbQ8kUjxO+B9QxGrFDAE9AZI9FJeSGobD
FRYAIQIcTP+WmaDAwcDP4h9L7RG8mYB79N/HYOJXbg7Nx2PZJLejqoaj/EgoCk5quYfEgr9ROfCx
EmCIktHdt4ssRoRDlVb4XZ4D91sdwKzQpYfO43Nvo0IJvKslavA5RXeRyuI4jaBn+rzThUQ1Y/Kx
s7uw2qEnRGtL2UhJyMx/FqjTu5QlvWR7iUHIvsHIC6T5rObpksNYiGLs4R8Hb44U8/mi2EUoLwvZ
5NSuSX+Hgn3bG9BG8Bd19kCQwTsUw70u5dL00Akprkyt8TLg720h4VIAVk4njihrhP/QvmUjJNgc
huBrfV0CafMawlj7WFrRXPeFP4cNGgqWTgSMZKA9Oq9YHz5roCyX5wwUqwV/dt6Hj2Q7fOR49Eqs
J2pEekJg++c2m0ncuwQgERKE4BJXQgbb+j+VpKsKneJO/4ENYxqqPNdlo5em8FaXp2vE7ND+fDcZ
+gIf7fMm7AK/mZNQ88/n9y0tSD1gH3NQGXZrcwYayWLFji6Wka27QGnlJXxBWhDsjy+myxlf/lbt
TJeQbS5jk38es3Zv20458TUno3VcE5GWN3ilrq1gkGmJtZWQPgOkfniRf4/+3KhwS3axB6Y2QVtl
OLmYaC+meRGY5jv0QgXf+jqA7ZLVozpEB3ZRk1k54LTrPekbrgK0qVUVTyKltNfCAKdtdw1vwMFD
lr/iAzCZlzLidY4Y6N0y/ujA2Op9sYS4mnq66EC+sR63x6BTQRmMgzmS8MnZ47+sYO/ORrCFvpLF
BbKZVoSrz28mk62B6Is9ZeD0JeL4cGTf4ryiGGInJRa4Ji1oyPctOW7noBUSmFiiqzHaWqL1IZG6
43Q5qwgcztVl2dlQoI46CUDzx2JZrOCHb+YHn9bkMspRiaduSU2xgfCMV/KjESgdiMnVOMVffva/
ieuYgjrUQP7sfqH1biWhUt+Zrc8YSvDnoV7NdSz1N7ZJk2NtH+b9ZxIU6EfTFfOzEP2NR1aMsUke
GdxFRxAVKa9w3c6+1eQvGzyhad+wqRB7rEz+4uB40mCHj115SFTi4jelEPcZm/l3N65i4RlH7JuS
yr6k37ALRMuSpEnO7vYo+RkKq6qgnh9grgG323Tjz+VPl02k9Sa0w4xtvNJx/lGgLD3QOC3uokEF
5qkhVfS/kklTCR5JzHSXtWYEbzxRBwYxAp7jT+GLHID/pl0o3bcHH8aqkA70gWN7WwV/cb/f1Wq+
0zutfH3V+yGXNiY/Tx47K4oqphyLFSTEABQ/oEp/cWDFxksCJHEAocxExGAd7DNdMOSTu+8Iuslv
sYBnhswe4TAMByB/+26jrrbnrtdo4AxHQh+4X5To6bmMmji2c6I0d6U37ICnuj7swh0quhP6oH0w
RCu8gNsrqnzE+Ez4a5gVBmtjmDCidzz8qhhFLlg12fBQFcJ/uBzDVZr8fJyRdBxbw3R6vXg2x2dd
FYuWJpujoEe0xF4rESsxXnHGzGVAYGCBUM1kXMvTOPEPWcHsU6U5pc+I62sAJ4IvaD/wvBWeDEnA
9Yzd8z4+rJxnROtwutXcYjfFsKKkklEhpQvjazW1T/vq4Tb4NUT9VMobGMpOI5u5Ubq+YhtDir6L
JNK47j+8dZQpPpJ4FNCvOd+zQx1HYcDiJBA6d/17MqFfW2OIEJbXTUiXdiIId9J8hwhiLQYvYMis
cWMLK9w3IkRcQlW2EK7b3N6zsheg2IOMp79KTD1dBMHG8YoKUB77SmssDJJUaxvlL+7Fuz9DdcC4
sg9pasWeGhBEp20Tcc+Z0wfBiH5PG95u7Tlt5lgzDpt3ResWyo+Bd1nAm2jBK5vILwYuKHnFYyQo
u8vvOST3WSQPjaXNk5P9S426oMFlyQmWivPd1Idcw/day7YVWgvWrr2fJfHl9KAgFJ06BLhVBgDV
lXMgIS1eB6q/F/8V1dg4PN5bDi5ECzmgseajvBeWHajEtfJq400Zy9eGOfE8TPDakhQeNN/Mm3go
ubVe1TeLzoQFc/z3q1pjQ5kXpRksWKUISTfiFpLTe3z0dFFJ/tU5pkbtkhaPjmn4iHHVvExPKxD8
JiMBaHypgvyqhYejBaR18IQtKgiQ3QhvkYRaDY9SxFC3PEXQ16BjHL1ktpH44o++E+g4muUpl81J
1eQpoBaNl/jY3x/Rk2GNzpIGK/t8TTi9eKKjNRxasyYQY+WTXZDExtsva2O/js/slPDD2WLcFLQ/
geg6p8Lb1hzzRvunb5w2uc0DQ87shp5TS6IlU+lQsaeJbCeY1J7qEH4recoHJlVH3Uvpy53o3OKE
CO7azesUgN5SfPsbugk+X93ykBUovW8a6W60uv0/FoyJw+H5DfCMUBEIp0gEcvvw1BkbZHS4p9GN
abwbZALOwI3zHecXxnqLB/SJLdHRQz7VWddy6fEoNQWTkdbl2oEUFK6j+2U0t1GRyCy9qVVhSAsT
9QgfCk/e4Vkfwr30inyElsllUYGv9HeEtU2Yyytfrl/kuVXz7OSbPcfNz8qz7/IL27pN46KtwUus
Z94sbTEZjjlozkyFP/WW4vakXFNBfWoFbyVgUDD7ezEpQwPK7Jz0kkCrCjMUvicA/RRUpm2QQ62i
t7bAETDVeF9oTAHoIdo0D74pyfMNbGYJga5FJlNNpx8SDWiRkOQMMNtIyPvuWy567elQQo7FggsV
aUxQVMWR2fKIGVZJG3Sc1kzBLeClSpB1NnC7XXatfeOV66hoEJ+wsbzFtnu1QTSikRj0otGuA6A3
dQEzKStqAaEl8JzKVYpblMRJMxdbB5o6eBE5xdaPXp7A/8niArDmVahpG7sCSVoUdvYz5axEo6m1
jYvXnRbipHu7TaLBXy1qjfNwUhI54pbYybShQmLAXosbsdILg15bm1C/3tzKIWgpPnuac3zMxAWT
x0ZxinXeJW0Q6BqAEqpiLskmPjUu1DLXi5SyGpaJb0KVyeQWZ0hJuZGYCVDreoJnAKxvY5wAYFhp
HOGsmTtS7qd/DUItQQFqNdkhQYh361hjYac5p9s11B9HMJD/P3iOlFOeENN/utxFoR6xTP4nuXxG
xEiMMk2MQYUePyhohc1xAPGI0U7kP17I7LYeMVfgEubHvdeAbDKyKvPuGQGfn4MYbIKiN0HVwQR4
DYN9fNaF1hT3T0KL1oF2rStjIN7aMEWfXP+fWzgcoNJR9gvHBFg9IVTAxV7xwytRFk9E15YYiqCh
4vqlqo70wQ7y4lu8SjAmuxKIkbljRq0FEfId7SvShfjFQb2AdfPExM/kVTNEoAbeuJM6foq9pRqB
wQv9LZ+W6wGTiEtK7JzVvnGaUij2ZXMk+kOUcj2ukvHfWS3Fc1Sr+4YVuLI4A3hllrWQIep6lSQQ
INoKu6KhA+GLF+3HWCY63SF5Hb8BS4WqYLjp+rTP8dubgzHPsm3KoUVbGqqYnXMTdTakJsyd5HEd
qhDHawJ4UoMQStXvimkZsuHqVQ+C+lXpl0Jce6tHgeFiZiR9iFTe/y6n1r8k5XUX7AY9fbovCfzA
cgWf4ALwfmXcRD9uHmEwe2gl0Yx/lMYoHjRiEHI66VuWuoYd9HpuFi7N34nCvf3GqeUEq5oUXWa6
WgWzp9eMaP3WauGvWxO/rUe5FHyEegshxLEUrx+TiQJY5QfeB5xzbNrcdOy/tuEFj6spDJCmYFf3
U4tGrx8/eNTmi3GQeOsZO2iV/ZTBH1ydj30sOkmVMtFzQydg8rPYzS+VH+j1o+i6wWe4DmADdn7E
RmGrbvjbq+fyMb2qeqTouvJV6E99je2bAfGezi4qKeXy+/yVjl4Rz+Ni1r4ZcWaJRXwFhJTFg6TV
9DNkXtFUFX4WK80v/0w7yvg9K9UXcD4iQAh+OLc9o4dO0Sd8ol7TuBTeQgNHDtE7unxc39NRfvNk
w0kZjK1YbUr+Wryb3y9JzrAwPSC1WlaH2BnjHQ1YdzmMcWk8bv7ZKO/DqD8WVm2uzsJCZzbi6IRj
5D1bNcq5GSCkMnnsYshMFiJ84AA31Cq7bFxrFWTHPtB9f3KQ0kiWuF0oQhJIS6T8Z3tiR2AdILpT
c227KDBDf+QhLxFSf1uPdkSsJYhZw4i8BkoL/DX/JZPqj2jEmqEDNx53gmigrdJ0kcqC83FfD8Iw
pN+k8GyMkoOqhreyjoEaqcQoIOBOVGZgIUZUjat+atgsLK84OxZulqNh82wyZtk0yjuvOX6MWrL1
BWwATR1+Fja5AbDJsbR7BR+TLhE0gQ1iuMkXHsgN+PnO6h4XBDyXyHGXCYoxamK0eZOqaVdWSE1u
ufp5yrX8nBBSQ0k4PzxrSjXGC4Cc1X3HFlayHXYeigz9RQsjKaulY4tu+fjpbXyJW4eGBbcp+Dgn
k7/gWEmrG0CVuhY2jYcyWSixaNPkv8gW6rq35mcjTk1C0XmWOBbYO7vgMHYIyX5iygy7OX0knddL
c+/fLn0LZUFciJ7rk4vy79XiLoGTCp+zSjOMEJN6+Vl13Qd+EBXW9Ls8WUG9PadddugN1Pynw+kb
6hQpv5/q+N3xcud7Mf7qyvNc8bzUniVYYt+B3u+Fr5En/qoUA29Hz1EXfQ6Fr4ZJekaRqWegRJGy
DbZfSSrmGM6CtczpiyEwlmxNXa4F9Swx3d5MQiLvDWF8QSrKDXg8s8Pdbv2vvYsV6rDVPR3nQJEq
rFkhRl70imF+ckDtFFsuaqklXrK02DzDiYp+Xy5e1ce5evb34HXIG7/z/rURWRTLSHKB5oWtCCZ4
EeObDtF0u5TNY3TYZUFlX2iZs1vFFsPZYePF9xcysruxNnmsYQETCEg9ooxWK4RkW+UREVODDHh6
2G74y6/YJxkk7JRkEDG28vbDtSAGCnz1iRVRNhlEQOqIHSqYpL93lsCr5ICPDisPiDSkFOMsuPRE
MnXF7d8YxnpiNbujG9zCiJV4/FC0BD0dMkXWPa2mCDOhU/1jek3/pN7mL6xAE/aoXqtuH3srQSQx
p8lbVigws8KBheRzpt1xjN4cje5wJHWwmTSEF0osXcQQgFVufYEUBJ488Pkg4NnFP0E+W7iEHOt/
8go64C53SbyXt/uxUrCjuLb/+6m9jMzN+HeCqSt7qo9vBb8xqkbtqPXOeWdccCV9yYMLxf7/TxVO
AYPkUcr2/Pvs+HsIy+APtf0CElpUqm2NMRN1AQEgXc9ceFSZxNFgQSI/0mI2Kv8ZA0C6CFCpQfPm
gzcDuO4w+JCefGjlnhaMOwmZC90NYaDn4zd0evKCGynFZt1y7HtHUc2afXNSo9DTwvOfCW1da0f7
Ih1aa0ygvk/6g9IYkuIiEeh7CBXJwZf613SZ9ZEGodPc6eXAQSP8XD9YAFmNxM17eN44H0hpFIub
uu6D7wcdE+2vt5ThpII9zO2ubaDrivGPos9iabLmleMYGw8HxBNKz4/ZQYj0kwXM9v/b7uEb00ue
FrP04L8LpXdp0ZI/UK6E3+kuWn7pt0pRVDs6lomvtmF4yYWJvVNWDz8mK49KlhYG6Ix+1dxnM4r5
B1GbG5OXmUlAyo2FRRvspV7si2Sbc+5ltxgvR1L3lhXXJ1hSNuFVb4QYI/J7zYRgeydJvmtRar55
6E1jbTl51xiV92aNnpu3MjkIdXBpcqpPtIGd0dIj/+TskQG35IqhW2qYj1sdhN5MEPrxAFGsu8dv
jIhhkmHFKUu7R5KW0643aCfk3jAoDRaGgsS8CHC5ydfluWfgnwZVjtLBR02uvG8o2qEbwElJ/l/h
X/3RYb950L/WoI7gyaaqNeIaMU2CWi1GwJ5B/biFcQRD/JO5bZxIt8RjeMBC/hB74kP4RzRri6Gp
AmvPn3ozK1Uk9EOOpt4PLrkpA41XAVgLpm7ydCzvSTDQUR08epEoJMoPR++I29LcPfil07h3162A
fE5eaWijB/WSWZLFI9uegxpbLhIqs3vLrAwEy1yMYBEVzFh9vDHY8n8rPsemBL5dL93dsOKA4Z3H
Fpctd31ATq6vbDKpzzbRjoflF9gbG73SrfG4lxwcj4Kxl6D8X3otZOlZG4vPUvJ3kIPWTPuS6tXD
AhtrrKNjQ287KOZkMiQKrvG9fM7917/wQDGZ2q4QHlPu1fnbPVC/kQVbvPGb9NlXu7uExg3kw7ve
Zm0nH4LRRELVtYRVNNvMICTlgfbr5h/dlAI00htx8JKaXrh6mbefM95yiYXHZajhr3UB8q6nGOwB
F7pzPuxQVRj9MXISo6Zd6gavinlEcFTGVY2tNF39/OOtyIIyQCW8r+McnygKUCKe6CX4VIptU2Hj
aUZemXcu+ITJu4K7hcC6XO6ZA90JwfgGHQHAAk9R/EpRsPJuJnMf5gknUAFlXUJ7IAYM4WYV7Mnp
gAqp82euqyGy1hwS98tSqZ1Kk4zQ5JgeWdSkZmmbK17ogHlZlpSdM/us2OgPzDSop7Z+JVnBR+32
L+uqF9eaIyCI/96bZQZg6iusIGHnX6wAjXmBGe2lFUiCf8Qq4dXEBOIP4G6SaR6KYn+wHMIo5CLi
ukExroMc7QHePEKrEhu60ctezcqN3qxRQBM+4UtlMsaIaqN9KS/1QE57Uee2ZotB5Vfi0ANfZZwk
PfUCtCLR6MwgOeMUYlxSfO04DwQYsU9O5MXTYVIUj2+03vMSKG5GhAnZjC6N1r7jpEQSCy27RnqT
3ii6EnPqWg2ztgVUvZCx/Qe6K4szFa0hC1cjpFTPHdOWhKGwBOuvq5DsO6O6QCf1xFqOCQIgTCeD
2FJ+t8K+YXd9nEIzAGkLz9wZyMJhBXT0g3UKjhxn4o9PuIH47iRtci0zKLeeT2Doexrmoltxrl0h
nWIL5+crC0ov9cr4oxh/5OnJriAEoSvUED2/jx/NqZyXOhGl86KzyVJ8rBeHCTCJkyE8LpqXKrGR
vwjAKzkK4Jg5noVh4qZI3dn29fjaFCLS5NcyBk5cBLAhBs94Cjv4tsv07Y17cfKeeYH9AYO0QaQi
JJ9sVodksU765d+Qw3U9Cu+rT4/xBLIkBAeBSodwP9qyl/Eydm1yeCf/eD+HQEcqKKBsJLd3XqKD
mXKLlG8l2ISyl4SWMNXBq5CChRxF6fncRBqSmTkuso/1J6798hvAXMI46Jw/7VfE/FXxsfUKCy0S
Jcw4DPbpF+M3IT04U3u9aWbQnT9kjxpEpta1MqgXN925DQOYswM1ialHe3JTThCBeIVznhZMzo01
S+om461d0/jFBar6g5+9lJ5iAlLjrJh1+jU5sYItQ2miLFR+buXD5HQX1L//dQYY+6e4Yt2M6E2T
TNyEDmeEy/uRtL3wAW0rLmrEabs+wK7rXAjWsUcFjnsO5SxxPcc7EtdK7IZHYnad2Oh1ZILHGXr8
vp5k6QA5ZDrP8FLqOjAUKjk7qM+Pg6lGydB5q7geAJOwoA9NXLrUSbfhW0vYyfpqEN3eMbEGsAsI
y8fMwtpcbyszJtaHeeKc3r0ED+d2YKITl0qbNaks5vbQgaNVA5vXHsp2cL7NlfELNUWFI6a1xWD7
Q5fA3EG0kZsmPJVW98J52SYV0ba611cJie6ADxW4cwNSZYguC1xx26gmUpj+DVEIuNwjO2nLfsRW
dTI7p+ccuVslr9+gluyTpKJ9Wv/wgWRFSbCWvE4wkxKm845O2zkIEjMZ9LfYfp7NFjCJmfjdVIYJ
t4Kp9vPTbxghS3XKelQgrqBt8WRyyBgq8JAWsdwp6qMxEnVfZSLyftMIPWotE4xDwb2qAV+yIvV4
7hA4yzLUZhFkt6LkNJZtB+iaWUIPbpI5XIHZiZL0s08qUBIGRSI4yGx0ht1KsLmZR5P48JnvGcmS
N5E7uFPT0grkiyvQ9p4pRaJ2ENlLK1e9rewQ/lnce8paqy66WnoWfCtp0BXnoW3qLaY2SMJ8OXRL
jx91odW9jpCHten4umIrB29JET0EmdKjIKHVN+lOBuoaeXOIdVIogAAsclpOb/9flHjBLkEGoD5n
6gphgMqNLG2CCfbAwxKQrBK/keyzLJXIljDT5hySxflVwwjVUXczCHw/ZlaYiTLEuRt3VN58JrgR
9jrlTb6FL+Dna93ZBNQ0GCcFrXX+By3I8sPcES1bb5HEPBU4A3AIekOaohow9NdUXX3bdO/JK/bj
non+kWFzeuYBeD4pP1C5XzUkGOMnH48Bf8vNo5pyTVHCPqeBnaQJ4ip32+N427hcEpew2AGGXcmK
VxHh7YMj4JlEsPhDLY3aWHQvIfEUO8cQKoNbtyTDc7Uzl3Jlo/S4vMlyt1sBXgLrr66gQD8uG9or
Us8JvdMxuffrKn+Vt5PkVAohLny7p1p9aiKjQt9luhUc/lcVEZ4lfa5YWfOGDpTYPyoOaX+AkGbS
3vGfnUwvTlGg60h5nz36VwwSkjvcAZrLC3VHG/joqHBVNKH8MV68aHayFAkFWTTN2SEY0sRXXX3b
fs+pLarCYX8RzatVEvv7WdkrxUwPac1CWuvAKqcLqB8sR5BwyOUnQ365uca31P7RJdquWx4v3EUJ
qKuXHkScKekKqJ1Y/1SXhZdICLiboqGQ5dl6hh66/Y6AYa/hIDTO7ultO9YvD2Gy25k4d+Ka62YH
DMJ6P0P2zz4mIz5dP0rmA5wPIBgUXnX4Zka7nsMlk+7loxzUyT9h6IzvMhZenMBYvAfQRqEFUVTR
EbRTxySW56L0TZD8wwZms3izgfm0MQ1JG0ZBomyoVWbZF0lokWEKK7GEQcHPCIhxcNUwF9df8cFM
dy/ZZOOlVTgPqMMbO5AVKkxA5EdgMKokNq+7Jpfp7EosqXgjDhihh1qbY5XEbcizP9B7NdJakiqt
icoA6sshVdLULYW7lM0T9TF7M68xZbPNip9Uc37yMwE1L8oElASbTt/wvEgy4+TD/102ZWlMmbLV
y427fEH8Pnt+RjUWHPKZ+C+HI984Yp62wo3+RuG+xbwoi+8Msgx75jIOI3VVtbTOy+hLmo6G3s4/
a/XrU3Vgqr6fPYFQnMTyLfleJ0RAUcTJ/77kFJl8/rZRt3K2BwNgpr+j6TPZ6m/sTyeMC7QdAms2
H9wXndaogzcvDya8jD8tV5MCLPvjrnej1XZ3nR08YKKKfdan4gSO1yo67lS9NviprcHgBHZ/OfyB
jesIRUu+SdUesZ4Q29wWDVOy7DlCIux37AhRwo/V6kLulVeEkjOkyTYgi/GuwHlIVxkbRHysLeYO
kon0mJTjlc1ZxWEo9qlNFmAoc8H79og2MX+twne6xOPYzO9SwPKGau3k8rlV9s0CeYAIAYZiGRsI
J1BrRS76zcMyx5K74o7SikPedr1m6DJp06vbkdsfciqrRaWsgvaw9NenJqnZcPcf8jKefEAZ+76e
VR858ZuP70Xkwnuw5rjiPPnT4733BfgURHbPWWoBR2ucXNEgrG/uG5BaOuHnWxvgKCjhZOJSRlhr
ku6oBUzNJZYh/y+1n1Rk6Kk/srJ3BCO/EsOOfgi6vGyxR9+S2iD5BINM0ogMUOQ0u8t8MLH1TxrI
4LMSKEw4RIjrmSaWFiJOR63yraicbiBFvo6vmlD3RXgW6mlnVNDm1TeCmeTKXNxslPUlXzV2BXRz
Gr5K8pkCtL6IKjN4HMdzFc+UI//1uAtKEZweAJlpriwy1Cx5p1NymoYhF8N0j5vD7hunOW14Br6s
C+HxlrjRZAM9OKNJDlAvbGI4MA7/OggrMJ4WDdEcsYr1OEd5ZTO5RoXVNvF0SowteUjdY1aES4ft
yF6mtNDjWFlS0B2Lc60CcAgTwLSoauL849lNRFyf/VK5kJPhynrtECty75/Hl0TQz0V+albp2uZK
gfP3qsXJyxtd6B4h+vp3i/KOpPgLVQQNUPb/ldGwuvZd1rL5LM4FK8jYHhWbt2SAVEKui11Z1D89
IA2UTy1M+9oPfH93tT3ULcDAUYWJxOHIB70msRf+BkbHcGON8UNx9XhJORLgYZ9JLSnIt2J7K9Mi
1lR7ZCpPHld51hWl11wV65FTw4G02WLOG6FXOaC+L3mt6F5lyXxzMG6waYcOCcgB8uwJy5BCOpB7
3WsE2SX9m6lH6GOh/89yfi/oQ17r/gjP4v6mceKaKwxnSMBvzJ/KFrX9kWrKuH5FvdVpkpyy3xE8
gtJ5nC5VIkH0FkqOepCLTBTcMG+lBjpcrk0z8Erqc/bfZpaaKGCtFoxkMblzT2twaQQNyaGhawqg
RoP5Ha2fbDifO5jMXrZocN0AGXk3xMtuuWGCuTxXSatP+iflH+YYk/2brJHloXwyqQrWqnPgpQnA
Un/820U79awSiBo5ddrcDmUebGaFXT90Od7GRgLoPvooZBjK8eO6dC1rPlC+obfp8pPpuHKdTw36
MnL6kmSsUPqowEMfideh51C0NX/egrJgMkT/0TZavcNTsDDFzeeJqg9FjSKJ5t6RfR4H7phuY0OV
LwBUNUSbnIGJ/TkkrY5Q0yeVXkE6yemLkAExcii/FDi26HPcG3Qk/V8sHHsNHvIbFR9YcUip4Gqm
jW4qMGtSelD0GBrKtocb68xeX64hOy5dtOBZKcrXF9inU/Oq816P6CaQXOHJBPKOidKgVpqToket
BI4+gKsxPHs2IKUtZtBKmEXLsr+5bT5xm9w9SKPTsilNIIBCuoVeGILWqlLazom2bM+vo9X0krBO
ndNvLo+cQvi1g/bBZiKvOBKnItBibLX/AbzsCukRAjnh2Ml0IVqOBDQVy0HfypJ0UxXAszY+vDOz
aN//GC1f9H2LczSdaJaSQ6AgHLpipanJxOSrHMvr0fys/2mALoc3+nRnY5vPnGOpGipN8dYa0E2k
nlWEdLhckHD1YzD94Kun+cmQipjJVsSFhvlQlEtGsQ4BPhbL6U9IraGCtPL+Y8WjO5eWncPlVCU5
nmfifuYRSOp2Qjj25AHyv1HLJH9MjvrcaCS9lL3o7dKePUzf0HglQ1bL2nsLSLPOZLoxVzz7gJ6x
bWiGRfLlDZihOi+ezMhKi27Fbm0e2shAF50+YPVPNy2aLA6TbKicBjKb0xw2qRI52+gAiKsPTFPg
U8dRoqnU9zAK+jbjDzRwIQrt7DMt/t01m4uS2GxmSLH0Lk6/Yn31kfp6cPrbcMhnWiFPqHPjt3Qc
+FPxG9tu0fBXMK2bhnYA5ut82+kvHNBtH0o8RPDtay4qo/+ig5YcgoHBSAoJFUD+mncTpiuE58Ff
L21AdpA85lXNyMTDclpJP/G+ZoFMvXHm5xlwwpcs25GCVQI7fFEoUScMsKmcL0FBg2YH8pIEzuyD
6QSOK+JoQ6KHp5GC6FKyllPElsKrr8dGh3plNa2Ll5AjqAkxS0cdpi7O2wJYodAYbzLNX28WHTvJ
aaHSNoiDlSkcI12ngFNlRECVIXuq/ltE+yxbAfWnPbjpuhk4bQavXQHzcrkNzkuluBZhcwno1rKb
MJ59SxA3Z9Be+9X6QZ4keMWQwtKJGMF9dtxwrIIcf6qhMTiCbOUuIRfw3xk40sm3BVZnz4U06JFE
5N1CQytQpNrtXSTMRhf9UExkiDwLpfUbsaf+4QoaqJJJMD4ryaJhm26OJF8wUfKG5aJo6cYGg1Vg
AfuiYHTuPhjUydiOVZ6ptBFtIi99LgAhXidsGnwXeWJVriQ03bo8TscMHodAEVbz4pkN3fGhyAeT
FRJOKDjti8CsOQC91EA31+wh/9qmTjXcHEtPO9f9BaH0ham7sqX6tjP5uwycPtLxxwAVGKUHpYVg
tIaOQHAgHvZgf22sTNwACUGFbX7CVY2mwBFgcN+rWw8TIJtDw2q1nlHi0bNVUaPOxLMi4I+ZLrAw
6kNvvx+YxK8N1hngzNVusM8etWB2aDvHrKIcoP95AiHeZ6c94GcPUCeB/zlxfGIkPSjDPVraKRXC
RQVY4qGhd6QEiUxDnvzLMJHmrWEhKXNR+m0Vh40cZO5hT+H1CIoICX5Gl5wqy1FVobvg61Ow6r0F
x8hm35em+tSBH+NiUELsIv88VCtyqDQkzGpCNpc+mJYonjUoS7uylUtagT4AZ8w9IyA9kYvt3wse
a0I2qsu7ldjf1IpsuyUZN+8rUpG+ZzEQXaDQPtplcG7YWKYxR3c62cky8Sybb8wgoVCMqwpl5FkB
epMUBBDR/skWOV0lKc0jzpQ5iHDdVdm3zT9DO/oDMhFbYxnoDD5Yj0Nd52sGGN2n6bedKgBeLgJt
r+7cvl1QPI8Ro/z1hfkYmGwm2D2xm91jWZnGoPFN5y4tOgdwbHS1U9vkUIBKDaMkfPDNWA7Rgjf1
QXUqI/2tQt7D08Y9+nXWAkDdn1johlbLNsKwVW3VmHurqmFhiB4xB4/bRJUbQBB2YfLxKoBDooYx
rJ/BYKAqPkqgQaSJQVuxK96W6tcKTr+0Z3jy1kK48gDS7gXq6eL6w/pNKsILyZ7mDdxV6nAGz3Pp
DkSO2mqxWpJkQ6MRNSqsnyVvbnlRftxFzoCt+lVKu2ZsSeB0YJQ4oZ1x8cPkSmQgwKrYi8Gds4H8
8itPSDOzDUvIh9zT5OjNNMagwnww0YDNTIiH2CBPnJG0G1afFgajUXGe/H/rMBon3+hKAu2+LLnl
S3hRfUX3tgKrWfG6YI5ZyYHaJQI6Gv4COZQmyKCxkfyUTZt3A5AjCAszThN71qYMzy9ZVntKgu2n
L5Yzrdv+Zw05jZQiZGJwZh60vC/nu9Gf0NX6rJqnoj1T5ylmw4HM0lRiorKC7DxefpCCcUj6yO04
SnsYrehT+jMz7m3kCVt+5hu9DZczVtnEqv9pYS7lxaxy18RKpU+lyxPa4xHNFI6pMioH1rLKYi9u
ALhJyxzue60KnFDilRpiubOBsvK/1bA1oShsf3J54VefyijdmFKCFDxPQgCtXLmbUlXGgyKyM2+h
74xrdhNJ8K9DSGLsKy7AGTzsT0XBJ/mcyxVZmEPhvdc7IoEoTXAxKNx08CQ2dvRikSDKxuEHg+AQ
L+LGSwjkKSzE8y0Nhkgp2NwrDoKaUzuS7nTluxoEGq/DFXMV7fvrIJP1xxi+Ak7UMcT/LOvpd+z4
RoZRYGsmyqlpz+qQ6JpPZsATvJmEkkWeN5OtpGw9tRtYBaoZCRSUsDLZCRfdkC/gZ7QLF514i5bJ
dGmPISPB4PXqy1mK4uvy5gqRyv0yrohrjiAMgA3PXX0cpSl8m/OzGWNrVJJErUc/TgaDXe1SKi+U
NTCABXXAfY3G60aUnADz8064rxbEB6Rb3gu0HElCTZkzEmjM0E8CVO9UWgkBCjXN7ZP2dhPT5edu
o0edfKaWXGrXoyr9ya1A1a600xdKIBzKNrWvHaBccwaRgIfacgJezYO82lNLwgABq+QlqubsxrCY
iqHTlhtaL7+8u8hEfSX8iw0iOm/V33mhjcJkVUluxERSZRlftIqqAduKcV1ob7oNSMz7p9VxqG3I
4uGmeevVYhvN/zVtOW2QzRngoShKYghEDnNqjVNMLyRdciaIKMIxTnzvzF4rIoZwbEejgDceTLaV
76JA0t4t0WmrRkalzA8iBhMIQrmOgFl5gf64YE+EzZ/fdGwAolktaii6/442VVFeptZECC3KY5aB
p/CZOj3Ch0hET9pkBkHs2XJdIBiRL9FWQrya10/AihDcNq83IZtA/VdtsYfbiVBhKJIY3m3KpM3B
UpzI1rVSQPNOjL4MmHQFYqwm0rk/zCrJwGSSvYApP445kPkF6fW0RXFKWMweVvHf7deHmwxHEGeG
mAsinUVIXRxONym/22I/L0bLrfjQabin4GnyDGra3UZ1JyW3r/Ho7DaxrE/VeGfQQcDZ8cqkf77L
0f1suMfLP0khqUKD0XQlO9Co89+UDdrgFyDTgXFwFpoNOv6n6sPlK4Hf9W7cHuDWcShiMgu8K4J1
JF9M9h5Csv/arLXWNoOHbw3G0s89bUcPwzTCDY3ZpILBqnLANMyxTmueHeIERLSGqsog+6BW7cBV
cI9yCA8J6WZ7cj+AmSrpx0ozp4aieNJY1lTSd2mk+/TyEYQPdj3xdq7MYYOC79Bsc0lEwhPlHnCi
QeajvJ0INvnxyBvxU7Kn8gRW9DT+fJOGiQBxq9U8ZtR/Ilb0saEQy7p5xdh2FiZb1ohPW5vyNbA7
9OrcE91lb5ncxYjITSzM5Zt+nK84tGEAKqY647cYjAdFvJ4hWlOvtH+9Eu5fXUWV/2ZywMtlrqEd
8Jw6IhbnxfAEVkiB6ZAheUd3Jgxeyj1Caqbs1X1n2Qhu9rb2uRk9oieUJK9EL009b05GV+oSAlIr
M7+7ick5DzXfsMfQ+y3qGoNrrw5jyT3w4Wo4x51Qy6gjBKcfA5ORPQV0/fUs9opaK2riGbV2iH/z
930WP1fvm7MyGjMGN7JGhP/8/6GLR3JmlueewVOygtcdJKV0wEpUGqAxWZp4hHRXLaAVNecUla5J
Y/fDShb9DKCBPC0MH9T+1Y9ePAV/+11Q0pxQYysg4sWe8XtalcBSLAAPOGk4cEO0MYmqfQBrD1jZ
SFACAnPzPZ7Ty3lxG7s9sdS8ZteXW6OfRDCvL2QkF7Qunlv2OK29J1kQ/VydqugmVa41qoOPyqMo
tOOoMhiEDgd3Agvsb3i/ssBe425VGiQ/5XG86nIk5Zv0pCkc3PJILC0CzZ1ehHgKXYGRj/4ehGWn
WWIzCeOfe+R4zNO0Fas1P960T0F5HZ3pzf5iBrOceK/M+TG0MTnBkeYrFUFc08aykVhnp07DUcBU
LzwpnkLVrnbHHGr1ht5QtJ5xZ5rH3EhVVDYbTiKPeHh4aHC05BpxokYSYwA8wtG1uGJk3MhStrPS
8PMtQaStDd6phDmiblnS/9BniSOlFsZ6udRP2It2Zu3+7yrwk+9iYPhPnYWDJY474QoZNVdXFqFy
B+R9GlV3Dm5q0WHZX8s5CjzH7Fx27PksyMdJ1d0PErA3/DN4lZ5U8uD12xik/+CJEXYvSk3H7JlB
dRYl8ZpdmvHzYg3wA55oaQCIYUkNrcHikWWr+6yshes89Se37+l12mII5JquBkisNAq9ThwtFTGM
H365y0gCOFbBdY+aAEZcGLIWNRJnfLYS+lMC6iZAuDRvk0C3bDBZMHMpW+yDLOpaNRN+Mj5yK9vi
hIiBg9hza7ORtpI7EmUGMHmgQm/JIvJOu87xcJ5lQtN7j1EYR3mWnlZ/9tYMHDw/HLrSMT3Ybr9Q
lt/q3uqx5DWGjQ3kYTD8GgNiVPPZaV05V2S0Y4rSRUB7BkUCe0HSADeeC0IoElvTz9OrL8ngJifk
9abe36UrgP/S9aLwoyvDxuTxLW7f+c8jfqfPV7YCt7dCyx3qNwp4HTYvpGz3f2x8jdeMVqMlOoST
HhD/ehdI0B+3XL0Lv2MD2F6U1SrUAeA1HQzgIipyO89Pq9i0kYocjYFRxGyaNzBccjlbVOSYrplU
OHDXIL6+9nC0wY0d4lZrKDoobmcZ+NtB+j+3W4h+6ID9j47mIlhO1Y7E0O4Px1NHf29PkCbBYz0A
6nhYYPk8ZTak8wMqNWezPFHNZx277VfgGja7X+iSUBaxxz0zqhpdFgOfNQxIDT7PweWbKnWYi+QJ
wc0JXEzhJj6LXUZfZQGCoT3Y1NUASxkcAixFVLyNdN2p6MW13TUNLIR0jMZTu2ORQ1B2hdjPIL55
Be8qcLa2ks9KI9BNZ48wCA7SjQUz5tvlta4TDRVPKEtpH3L3eYmk0igOzpHYW5e2YkklkppzdXtu
+Zhi1N09rCQekhzy3PeTyUC28zjIRN4ry/E4hSpQjbiw6CMi4FRsZPb6WPaR3JliUNiUDDz0PF6P
ixlYEdHBPc4ewwuQVtQmglRH1SEHpEvNF+wF1Yf4QJyq1NQRDENguZLfoJfAasHbTMnnTDzyliMu
cWXSr3aD83a7UG3ExxijAZij78k4Oshq0L/6idT639muVbWp/2r5HFFLI5camM177VOQ2vM3HwU2
eQmtY6jPF+NhyNdlxavFZpncd6r2tPlkot7JDSLHDmQDwokBPpcvGlnuPlpNmn4oxuaoLcIZDNMt
tCEnBR/Epk1O9psXsSoA00lu+DIgHhaLvkEPM8BdYrh80Y5ZdkgCqVs3sW09eHgyR12AwSLO0dsr
7k38tLOVFz8ctDw1IjtHgweMOWuU9wetHg8c5cJGdMNvKXqj9FoJObt7iVNaGjBkX8FwtuGyNORX
WIJdTElLGqnEUdl3j9xsZUJlmoGoNV+pQWHWCNbi55Eb/ehJWBiIUcdPh67toOnSRnfv3ertZcGx
gDwJ/2tktJ33aEf1O9XgMiZL5WxKbEgq+tnJgTdmpLXJCXF4DZVwv+7EUgbESqEorAGUiXqD0h3X
UfL/u69mcDj1uzBmHPlqoj5g3rL5xwSUfwMNNzqt7T4pA+Hk15aQhzQfeljXiJiMMyBxDmjYSGjU
S5vg++A/3z4Vzx8gOILu7zUx6ystgXB2406JN4E+b/SpQWVvusI8vVgwn9esfDVubXfvwWm0iVzV
z5bV0PvxlNAV5R9GXRqfkc3RZ250GF9x+CFVlIIKMag5CRykBN7AcASuix/NqMqa+60eHtwQcDE6
5W8vUjEgaubYJgw5irhVbvuXypnM/VPCKuAlU5Dl4JLpbeg7PPbZe3DThVLem4WLEtZK5VvumziG
KpuduDDFdrR37zE+V51nxGmVBjWmNouYn9B99l++dPBhxnEk8vLwwENUDKG+Oxw0vcFCFODdhhYU
/F3TJ3WhLd8Zx6dE1qv2gPxY4Lu1TDnlIrqKm07ZtSRoeSjszDKl4CU8LhsGs0+fErT4UaeVj1P5
nrWScAJoD73JdBlpp6dywjCZwHzlfDu+hFOtzxdsnxD0q7j0SJIz5wiJ7UhwZbDm9YMefZYsNnWc
Jv5d4x5aMkPCqxC94OmfGCDLrpgDDk7GVG4lQN5k9VC03t/sdVx6XlSq/hQ7R9YtQKFayVEDEZFc
G3YKRXwf9aW5ls9EEPIFK4rcanigLl+QMcYdYT6IzE5AfzwFUI60SLCJYyw2SD6SMI6JDIHHTwuH
8CEIWAOFXDvut/05XFB7P7zqf1MNIKJnYKQtdS1oWiiKyDLVK23IFAWN4SaKIpYw7O81nzWADK66
9z1Uaa1cSoYfIiZhp9TQBOE8DrEvvwyrwGKxX+MXcIHKwZGRYzjF44jdaRCachf8gwzTe4hMMcky
JM8cl7STWAUYhdL9E2+Y86zLWQohOHoJWoCrvBKxsAbW5AiZOQ1oBDX+1jtyvdoTptycL6yYDb30
KlO3HptugyISmxupDvRYxNAz/iV02bd9HXMsyftLxh/9qF3miEEDx3ntCEDrt11bK7P1+x3OlcS0
uyCc0Rw/y5MnPI6Zp98PviNUxXaOg6D319s+s0XHBp6AyrySh4ZcC4sHCVPn0ktgZJaK9eBxYEYQ
aqqeg8q4mW6oZffbphhIByY/wfgB6SUmD0bTJvlrbqug21W5ZC/ieLrEcwZgkbd2TE5ztbNgcEbs
CCtbTbZu2FoC/v4Tiuwf/jJrWpCLH+JL6ux1yt0pjA8V7YSLbVBwrLNKRuyBS17uBp36MIdcXwzT
YeS4H4WxXrDr3UE0dj5MYSYDnFt5IeSqctIPBmAxzvmlbvqDEDf0yaI2gGFVscK9BMAUGGQEbnuE
xvilkMRYWdNH8e+wA0F1zjpg6WrgsghaoDJDN61bYOLnQ4jrfbGgjK5M1/Q/s4+xDHwVM1Es5KpW
Gks3gGp8bwYkaLX8RhXRvNibl2jGqNr+4u0K8wpQlBANctR02Rce28PoGnmty1uKRvoaSEk5aLv6
zsMT8Mg1MwclRTfJkcEqAb3Kkxex4QfLah84A/nSScYcoCmtdnH7tqpiIcmSoPsn4NzBN00IoOfs
a+TW0rnvOLTNx//dLbioJWvqHfAjkQF+Zg0dOCG0XoWkqq+Jve2EgmB5rWWtpKNTrafzPL99WHrt
hUmt8Ovv5V6sY1wHjpVy1k08/hNNLDHosicdIMzfCHRjU6h/8jqbimgWLmmqrDmczUyZV9Sn/zBy
Bg2DRuL1lJdv2RJxYY59tvXhN2V5m/YJi/LKEJIZlAGJ+yQ0Ib8mebs34ZGYwu2dtcXNzpIqG0n+
bSS2LU/DRbAHlOlZYGlC077fktNtkI+k0+xZQee6GtL42Fnzi/xHXOfpxX40ZywtjTAmXNJan1Iu
9rN2nOTx8RmYOmUJ9GycXWqoBkFivc9bhjQsyV9uSRYSkOChihDEqlKdrPYgtZrpDDYbLIbmAEv5
dXX1Aze/LgG0Mxt/4L7RzgBzvVPD8641DGPR45bsuCsbc3a554N9hi2ZZBZAKklLZiujuSy7E+bH
ZJIvO+hH1DXFHb/E6SFXQKXdPVwH1pHt8AHEAR6Eqmn5YbF3eaUjaH48e1eWrXBjv03I/NkYl/sw
qnl6ka1cubFxqGdLZznWOpwjrOjFsX0UxG7IKH/lzT4+rn9kFXKTIiOJjLne/aHRXhw/TzgCy3pV
wDnjc2llc+7E1J/88WxBFgJrQ0UrO3uSOPbU1iRvK1ooHPkHOZk0cXEp5EHKdwXJqTERzN5ADJnK
D+m5kMXznwPfosMvLwkMOTFGEc+Imq9U3QxSxirQWDrm8izpR6jfhT5UA/tn86OrtArUXHxLZwyv
T8PRXkMx+thDW7c9BWwtQstjIihFm+/FLIthdZwEotcx9NXG2BVt0mI8TzO0U/5zznler+PMwa+7
THQD2rvkvqykWY0A8U/UaWpX5/yBgfMwMrEPry8WPOOH7epRgKnLPPykwFQ0mTN3rnn21qJ5WFjS
0WEMCpSlnUM2im/XrYC5pGcZl+WXBzJ6vIkVc7mMeB4zr6OnkYW8Zdyilj+5g1sZILfJXRcUxQVG
YoFX/b2gY3ya+DYADQqh+rfXxpBvsGtKpy28aYDR6Aof0j5cQdE4D9NB4RIV9WRykjTGb6pbrhkd
SWHzQHf9i48O18YdR4QD3XfXXwNKkFGePgxBkTYc/D/77A6CUko2fTQUqlkPkXL65KqGWTZD+CDV
mwGSsdI0IyWXRd261l0fwc5W12jzM5/vFb9Ir24jbw5Xo1xSjYTcre+kLhGZBM3LxaGQs8ibM4zf
f+LGKQ9Y5qNsPYS45Wb05fgEtvmyYlWirTz8hQ+fdlQvTP9G6o5eEJVPqfgxjkCrRBLjs6k2VjJx
8n9gHuZZWaZaeGNZ0xHCEIGtxEbeag+8kr3/vffiSYfp9DyKoS5hFOX+3GhNwKuZ2juvcFE7zrbz
EcndN34FXIGLOtAg81jOR2ES/n1SxoP10/lLy8+QzHY1lbX45zLwURl36HwYh3i0gQ0nLcf0wEA/
AmQT3vcIQu1DPrrn1r79je0RfX2y844bRx4fzyEtqOA+V8AnlQPD4dca3YtotJh/lW3U+CsngYa3
37RadHCPFGaD7on0h5lbau3W/VYgigvs1OFePD67td2PLYPtpQXVEWW35a+DfuX8gCiWrZIsJeyH
myuMuTCWXjQCIEskmxz7eUBRJCEIB+iwkqnoquafOyUsxiaP7HbFE/CDNiDfvYUE+rsqSIKdfpy2
i3XWi0fgxBDARW8t+u3aHIHv6doxG/KdJTpiBoSihTLPMZvdQJDCaHlc+fVes5jDoEYWIHtk23Fa
3/ZT80hJnP8s0CvNjI7bCuEPzpSgwZmcEXf+nUHSqd8bs/51sHiMVipmMI9J+z7S0qFeklEBqzsP
0XE52ImznUvgbkSVGzfmHtoVTgrO/F8Rng6SGVq8A/4sACwupvr60tgHYWWxX7qXQjFtHQHHAj77
hdemerpT16HMpBGmK/VY1BKMb4c9ZQ4tu7r/XT/azKUy/FoN9OlmsJ2geo1QvfKaH5eJrDl5cW7c
A6odRQj7I9o/vOk1A5XHlziftNkbzHG9sDCkXN4nCgKYDWEd/t7VyaHGz6t4wDViFgPwNS0L191Y
k9B0Em2YWDJa/EUcFKc3jMsypKogvkTJSlPoMJGVpiFbjk7aK9wioJGgW7ixH39BQuns9zLLu3pY
jAUvRKp077yJxCVcOi+o0bxsKRbINkux8K1M5LvXX1PnThGKLjQVmkMVlokuG+KztnXYQMgT/i+m
c3lK/Rd2bVoAgVuRBiuSSIF6sYCArsC9GF6GYtLwziJ7beNgbaPFnv2bCtTrwnwdfw+QFDUkDjFz
QPyhwcsaaU0Z3lFKEz9WnwUFwy85rb8UDG3K54aAp2/gIaSspKdhHDOXw7o4pmkwzlJNMkOS5HX5
VZjDE7nvFwH9I2zG8eFGf/r6f9leUOFUxs5Cildqd3aoQ2B7q/VnKmR75fTim8e50ho3e3XiL9Af
fHUHwZ3QBU+f71qyAefUiimuPiTOvrEilgxC6X7Nq5rpJAfhPGLAvj68QdbHFBf/zzforU2aXDjc
/kbvSuL/Hew5xosN+WgPis0Iqwv/zkcwXUYqfxxm8sHZ73VtVDWTnYg4HL9l2TZdL8vcBHg2ke+s
oO+WWEw2z1cqZklTerWQ2cdVRpl0uRCguEph9/NsLWUlJ1Ze06nQYiJQ5RYSKQ5kFsB7/X7fObXW
uV2lvqsifNU7CiQ8L7HDuSAx0F7CUU6MlDvzXokziaHWy9PiOun8lkYYMU+1QTs4XhpjoSz+9Co/
aMP0LtED0jvxk6+4jwtBY4AJtCcJfnYu/DwFSIYY6sSLgeyS2axr3fdMUjJKrJ21UUhR9oKKSHCU
jmfXddFTC73gPhZqqNweng/SILrPbRDDCqUeBnpy1cp9Omkd8MGduX9h0i3MPUSeWT+Xoq9IAs0K
x5yYKp5l4IOZ5OQGYOzaGt9TAWFAjEXBVeaOwAiFD71PQEZ4RE2JX0LwdivwxYx/okjq3iCg91N6
2qhCN7Hsk3C9g7qBVB2jflb5g5Fhx60fl5MnNP94xjkqMUiJbTCFxdKP0OFrNKxK1I1IeFkkX1Vb
6UZEIejXS49vsNtmHt3smumHS6/DnCQFGiUJQSIqgiepzCs4KvbnOU7Yu4SKMiFxdIklk/NLJAX7
b4PrwmdUF5eHwTHbWMCajSEDn3L+YZUlrlLRrJ5qrVBborcmK+yyZ8wNKH9liRYfXtsc/20ZIFdn
4hS/5vRkEPJ4pG4gbdw7jFR8C8QLf4uyz8D2buIxVILXEhFIcfX04ywYyFoMG863hSrawLywn6/A
65eeJGIb2fjiPg84wCiU1p1ZGx2K5T36alBz/IlLzaH3JcksrLKIR9cQ0Bd1g1Pgcsg7+pOx9E1E
kKd97holhjLvPlnc7VSmk2aTvG8Hi5qOgyFx5LN3XKihMPoaZ49VqPdFUlhMtKnUZFtMKjBtxApn
INYdI0baYsPJsw1tmaZ0r9mpZqJTNg4XZOhPwTTBLOZkMlgPpOm1TaW4FlwWYkgWCP8Vk30u9jUl
ALJd/DtC+X88aINymIDwBNvrCL0vYAaq9BvAUhPHh3kH4HJuiQ6jLKf7V5w7WZyIKQaoCqa3NY4M
NMJWwKdSsGH7DefcazV/14g17+PO+muRBEIPTk4K9kro7dO8OwiO3wBiT/p5aqIC5rI4VSvLKdgr
gDEtQxhGLxk0jsfTP0er1bxlWwdFhL8KTCbdldDZllSGx0eS7ygih9BmcL4Jma77RW0BNR2Q/Z57
WxM0emotUTFOUeeJxILRCSLRrgYGEsaMgOraUeMwhKVDYF5noi/xy1+B4sy8hR6IzvZtv3i4rOM8
4BQQQviwl23hr6tUIqXFfHrsI443M29O5vXeiks8q5Gj5qgtJUezhS4O/ocweTprXRA1txgDhr/G
BgP5ad7lYKGZ5wZAGlNQUuOCv41lZ1OxGtcXkpsOShYDeC/quPt3MiYYaS27P2RcMvwoLS/DtNn7
0HJl88RGxXGE5hz/9encEH3Q1pwA/RQ1Keaq+70Hm0aXW8PkENtgV0VVVgrEd9BXbNeKLdz54hyC
ql3JJkjVmb359xTXkdFu7d0YFI3GiXhAdFZW2qwD1stxSFxmZQ/OyXSdYSeEkLlAp1naC/nadioa
P2TE2Kgnv0+y6mLuEjT6t7IvkqfxSHQWvQITKxo12mTzpAPoc6YGs3rOm1izZ8eKFWhgWM9glvoo
vYA8NwMUOQj31xlNZYTlf1U/pwGPc8ecqCzy5uWEp7ZHyan2tAGalvF+9xjx+vgodAZDUynh/DFR
LJ3ilp1C4lMJ4aqScCE71ou1ngGI9lmrW0pqIINkiy6yOcIpC2WLbORW/LqjK5HtpXsTcpkUIaqn
iVtc0F/uwcwZnWVMyAPWxgbs0bSeYQejCLKfEYu5ctC05vZpyKM3XDbOe8pbVb7cNNMwYaxqkgQI
ajCgnzKB3JrzOkzkM7QVlDAAPZYNdg7hqgpNR+Cd6hvs98kUAuKu5a1U+p+POXB5dOmg5HL7r9Qf
5jAwPzoGIRRYY0v99jQhv9GnLChisgj4jDrIhYNdkB2WJ1nFkIysOx7F7at9BEnERQ1oF6kyqxUx
DsQYRpLOHZn3c6wi7Ol9UlqWb1owQP60r9rEGjO0YCZzuaw4T+Rdn/VFQ99GAdCbHyOnbr9Wg8A/
eUz62cjAYpBCKZPSFX6jDzTh/YuXCCy2NPEJ1FMqPSMwi4wZNb9dPs93XreOsOrl+LalntFQFZS2
gvlI7Y1HPDJZNahSMmh29bHCt4jOg+AOTzzNNE79EXs6hz0mJMeCVUAy/vZw8d7TSXnGhGnMSItl
ED513EX5UeBbvEeQABLJWQvywcJ+ehPdwnI6yNN97GzGc9cqCB/pDzq8Pb3IKd22YeR/DPPRyK4v
/sJItiGuXtvJF/o+CtgXft2DI2gwqTPTkxuaSmS8quqX/ypQZ/OCX3Q2RFJgvoV3ACu1NJ+v+Sq+
EGLN0klYSyDM/JNb+XgIoMqRAshAzl6fZW+oTMhkfhKD/FHoWkmHMb25oo4n/VjB8GwKSaCEV//w
vZOgTdtnfqSirEGFLSTCOb4S9pKqgQ7J22x6035vq6/lSHhQakJBkr63mGWcWqrwCY0p5moH1E3O
TEJtfWvyOWAdedheWkC7gv32sevZLS6zKQtjdHjq5TPhfE6FMM5kDLCBJb8+3fqocVbq9bkxCRAO
lbyMXk4k8RowMmbiu0PT7LCMdQSzEW7IfDd4qUqYMT2srkypZm/Z8uVsGFk3yc0tZJXwM8M9ay5L
vmjUV4xzWITVLAeGelQZOZBk7cRFr0p4BmZwjXScOF6XqQhp6e743tjHpKdI0G/FJl2s+W7rPuGG
Ka955oiFfg+SshhFAmE+Qvhxn25CcnvtzJEVIs5e0hCMQaUvtYeXudcCgDkGaZPvnJ+yIFs/lTDn
uzQb3QxXeXfu5CFXNxDtkuKw4yHFz6viDePxJ4N8bhSu7QPtu/tgVAwAFNKrJGRcd0jRDc2ijJhO
ZKE/bztKCZ96mKN7C4mkG9XYOWDRmLk36rQv12vUwVgzDTKrp1AkFHY1oaPN2Jp48dQFzg9MAcpx
1+GBdjGN33rQ4+P+MiMnLjcwt7e2D6nMQ9998dQXyYWUY4/CAFcaXjDRcrPAi1IxxxZYWmq5s+09
h8Vc/sgFsqEp/uZIBgaPG4DR/HwwvWEs0RQLeULZLOGC0jglX1r9J9nluGtPl89Eq7bEynaoSTtX
UDBXSIfv4sxnSsNnr0paFAH3MmvBgQXoqKp/i0v2xWKIqfHEPRRGmLFDUcoJ0xi5U1TJS8Yaiexj
fQ9xqKeIC1Hkf/Uq0rJB1UMh7yH3CABjecSxtrzWe5aiCo2MlQLuidAE9hfa6kMLLvJX7aak1vKf
cBLvYoDw8xhotIiejshkXAH37dxmQtqswVCXnHlfzFxOdhu70WUfOxC9PGbyv5mgifJEdKeIJsGI
ylEM5ufhCFIpX5S54C1fSHucsrnYbUHRDMyjnIX8EyIR7ylsBjlYWaOhsjlYbiomcGuSxO60sbV2
TxE6G4yTJdfdcncw6JlioC9BWVmjl6KDBOBZCZ43wB+2/RqFRRCghAdQMJMRZYSS6V6LpnHEGxdT
65MXLuijN3gFl6AT96g/qC7HajFLyL/y8ApJv/zwrZwmvY0LVhr33Jf3c1VhIWh5ZaAIdrPdv1Jj
ZTB6hSn/HDo9kpbQ3hrK5uBYZ8Ge2pR+NkqEicbXqnom/UsmV1GQByZ6IAk2XaQnPNXsPLoLfxrN
JUsLjCGi/00qR52yJRMOR8CxYU1e+DQaVokEs9186LUaAxU349r/q06+TXjU8TwFjFkA2XRDmDtR
Lu9O/LgdYBK6PsZY3/NV3Ds0jQaodlRQXNL3xYjjmEsQw7J6+NqRYDNfKBPamM3L2Z0hNlvpv5h8
VuEu/bRQEiGNHJJn7J1xV0EHtsq6ScceT7QTBBHGifvOPQv+ToIXnUHUBvZXx7F/730HnCHobWzY
0hZyf+EFUdklutgE/HMvkj2xV74tRCu2AwyDKP2cPPz/9pICygjlgzxmIVh5ZlCx/NTtjYs9On8s
Xxcf1C7XuWRi6+EDRODljv1XWfczKZRFEJpwrx/a4r3oZKzyVqAaCYd9/ZBoRYw7JfALrq+FKto9
9bK90KqCbQq4EgMkDAlFqjXbEkCL4entv095rmYjECR2KD2y/hQzw7xEsi/hGeZ5Ao1PqdLaBeE2
bBx8UqMIfwx/osVyLBFa9XCdGTAqlA5rM6vnhJaeQc4Hgp6uRtizHfTa92UQH4/D2A0fGk+g/K5r
qeAj/ieMSA0vvLT6TkNOvpkaAhZzzko26a+ok8dF4lFgrAaCLa2NJyDFWuTdwFEXq0p1IIP+POuD
o9eVTSr5NOCYuNw4bkAgcV5REZW7RMjIX1Xdm7+0gMK7qTQzoHN1Kb+Y+hhvq5692znQiwjuj7aj
hIvmoYYmKr+MbUqcAxFTBZjKBKo+OjPKoG1ffUzoKjHqeZwWAR965z7BgYM2vApqZIteGe9BLs4n
4TrI+MIAuQNXo/d3h9bnAfVvpw8BhSwW4pve4SYLp5RizNmjt5dezTDEynRj6O9FJE8G1EJ0pKHg
z5sZuQ73VNwd6nR9zoyYEUYjWIF9KvOUrn8McLShHNPNRrRVMfhDOYzn5y8gylkpZayfOBVaSEM0
lfin24A242j2Kvby8quk0GVV9XbPPfMqrZTeEmNHA2rq4O8Zh8s+EdgDhVDEKtOcajF0haF6h5q0
YfBzwz8B9Vb7UbDqf6Hg/gS1hwwVjS87RqFyYxI0tZIflVt7+j0LyVhYnh33paLpeHQ4F+OrhHSJ
92RFUzwyDVrIXKnoYLXKCzrXs0ScjK19+Kk93DMZekvYQKzkX8G4SrQnwK8OAFts9UjDEH76FnF0
W2UaLNekLtkJm89nNb3LqSc0AnuTvQJjVyBUTUfeRwdT2rNUYKtyV7FYVw6pijsoxHJNzg+I+f8U
hamUBVeKGf/F3m2BFfA2lEvCtLYCSPcTXhQAMgOM3BBNbNnyW5CLwu1X+ZyKVTD9sLxGoB9tI8hf
bJE246J0SGHVGD4PITMUkOrMzDou1mGnhqQFSjaZVrzOt9Sr/IJMIkBPNfMNcJ3SMknoLrAZGRej
is8idHWHnHBjxSmhdlqtQo58Yl58zAqvMBbO9K5Z3Dld2EFyGk5THjcDBnGwUGBrhCKPy3XJGMk8
KSHXVcb4id8iX0lFUVDKChb0finmj/jcj/kjrX03D0KQp8QI0WIQiyF/SaWj0yenFnRs4YtWDNPy
jRweqTsvt2Ti1GLpReNvhM/0e4PKP/YnBEkZtHi3j5AkWVqEcozek6Y0G+wYzHIgW1nGbbjxx/75
aJ4LvpgmtVI8VaG565qhmsEUr+cevyWResoLBYqRBs/QS2HRn/oGDrBHr6W9tPeyc19XBmDOkRTm
/4x/kZCWT6SPG7wr23qe1b3p6dX49Uc3yuo2+SAKP7AjnlRnoxNGYSBu+4Os8aGXpOSHTB1S8S9d
xJgJldbY2WyOUfrvtcR2dH+f4/OVFLtnSJaAeQK8T58UBhxBjZF0IMvEaaFjE8RAT0gIDAIxecFZ
GkgorRE6VaRVSl3Doy1A2Z0BZFdRGo0k0p09G4mtr9cqL9D9loATm0NmIutsaKskdRA6h7aH2rPD
Hhb70u2Z23zoZJAuo8rYbCyLqC2/Zn1AkwZ5Rz9r9f+AW1T2HvZIovlFdMUxeoksshj4LWF8+KYh
8K4CCRvhnSeh+2GywxVOkc2EaHT2dm2egfrkitqgAMpGQaPKtxauyENqpEOk7s6n9jSjKDZcTtS7
6LEnVY0mEmnZCKsrd5Jfom5VqvR/IzdtHKVml35w2l55f0cOS8ZLPuDPtRlitCRQt2WBbMwbv9kx
fRJLAQIHydxBDo2aZ+kRf33a2mDhGQnjyy78y1Wh6a3s3dPbffXqTzVZOcRREgBSHlaCLzNjOV0M
ceYVOEJjyiBNHM14vGV2+NyeedV8gpKoS4VRgcNHVuzchjTm9O3o1SjpxK7L/FD49/3h+qsK0CWL
IxcGFsGgpMQ1UN4ozhOdk5zIM3Emzpt44iNOAJKkMuynMZpm39yQHXXvsAvAXrRq8W3flkiznCnk
KXvERWQRq5CujnvhI2iGv0zOerkQFZbw9oScK7zU71Iy8/fNbgnYI/otbBoBaGvE0KaPH5BF3co+
dUSIG0eW5kgFzQi+6KR3UG1LCzm9HTblqEXfw6fgnhpsqPtYXzUoaPvV72nfObBHfKFisiaqqqFO
zpclbmo2BEQOEbRduJG9kKwVmbLSCnl8B9Nzb902R5FwDu9VjFufUMIE1CrbFlMbkAJTBEBQOWFx
ghVYfQ81Xm9lkWq2qlucMdLEbUXT3kI3gvJFkAAKTHZDfZWaFK4q++jgK8Tkhwl+zzshZQ+C9BqX
d71ok37BGUn+JXOeGBggWFhb7itYgTjTHgIET3QPuA7QPj0q+S/6U6B/NbsLXu0mZKWeoKvwJBSU
MJtH9j41ZLHw6JT00XOuo0H6Ohn31vlMG9megW6ZWEBeJlJvJ7VSk35fNojJ1E+nkPdMyLz0jBA5
rZxo8nWqri77gMYdpgINsYImSYKdr7Be3k9qO2Ab43dgz8I4On+4w8FCtH5w6/2ZbrDoLcD00bOQ
BhfSa09vndCqwce9nwwIR1/08u2LkPdfF/5xyMnmsnonxoUZVwdFZ/P6h9F0QPgL1k+M0xC+pSLU
W6vnN3TWvfx82k7MHVdq5zQ/82tZMNRhAdEeSvaUkPgWUP1PCdNWhQ7ZuOTLQlb79gxfubc1Ldep
deQ189/HX9b1DAU2n7SWKYJOolF5lY2od7IpXoQNZNYiNID7qzJlZTCtM4U3VDiv/8fgs8tuGSii
yUxC9lMygNiNn82IcG7kt/I5QE1ghyIkn3W6YcNToRO2PbesmbtAYPFfQlgO8Lfk4ulo/TtXrxBP
/99wpLVBqigsZkJ9pFJG8png0w2K004cr/lqN65BUM57QOSdaBGctVkosjd+P2ffeW464V523KCa
h+3btjP8TV4CWQfUVL19MwOY5c48xdFkny81Wu6aLQXaP6gNZbSogPNpNrwOB5jTTJ5e/jL00DFd
0Ub4CofffjrChcuJm3+ksYUJQZStCovgcyVQGlUYEcNqWgT78lcwjlE7tPgD+tVz2TsPmUUry1fp
n6ErLrj8zgVt+nR5v1e+80ujB6fHnZ2rg7ITkbSLcLA5b1vzr9r4vEAH7fejNClgqaAWfE3bsyOf
OLQAsVL3HsvgRsSwHdBWHB528gt3qOQDFb+EsnXdlBgAX8oyAGrukWuc7SqoHqNXLLPDYHDaziPB
+eali2lNDm/V4RAZOhTJjVjYTVssE8LHleMAzGr+9Qg4IoN13ublSF9IJAQiDq9HhjY4pQgfWdT1
0MgwcmWKLRQ1lgQdw0YCyr+zh52B6YAdoKO1Kh1CPXKX3a7nCnQWQEwFIspKU30EyBgxm030Xo4t
jAzsrnWcGd7j5wHfXcuHB9dW3ynZZCFOfN8nLhch8y29dx4yjdH+tpjQdFo7ZaisWH5x3H1vAG+I
1rO5Vh9vNijBi8Q2lmGLl1N7y/1xvLti3rrZhzC5wHLi6/zFG1ikziYYvXRQXXMU+lqRlprJntxG
bxxD3ckMpBilNlSe0Enfik2eQYJKAMUz3YCekwFv64acKQCndS/Upw4m7WH4NlgC2/UviV+HfCW8
r6oY14RxWUu0mTA5y12HjpTdZm+w2w8U5GgIa6jxYp3BHQzaoZYC2iIAEf/4+NG65Nw8T3BVxfg4
mzrWQh5GZs0QKGKfS/oFXjmwLCvdaONfcTcSxG5kjGCLbzGn3RAp1xbXjv9G8l6flAWopJGR5IXe
lBJmT8SjAy2Wpd8C0Igjku+n73tfqTa0kw2jp9C5UDz23UN1PcKTWzYOYRK9wX7c01aqDALqcOBg
cYmquAYVaYRGGgNcA/2IxfdXMZ5meKU/nAo6Y6MWXy6l64k4BT/tkR94QoXqThyKid1SFq9m9W5S
SzH4U3hgFeVVldkD5cGVbI4/w0zcvQoxv0fzLQX+OewXIoG/Uc4NlJzkc7+do4pCrx3MHdpFqHAd
kOZH/f6J/R6+x6oDJRHNN9ANTNqSd7wr3oypffjFrTN8dd2wjgJqxqHU1lHI00TjNM4h82H2NB15
HdJQWoA1NxrdPm0K4pEYNsHwvW8+rw1cLiaGsr0Ge5hfs8nlNltYI8QV+QX/phZG0JzXYR0PQ8Um
o14SLPQV8pEamFzHWeiohEQNOcHpYZxrrCGhkQOMiB9DCGCTFCK0kwUpNW2/zZZm0dmHA2iP+ckr
JwVNXybbG0k3NtYFN7pwi5Ym4IBJodvOhJSCNbWCFI/F34n+vmP2r/LNMGDueJVI6+5Fo+BmDfmH
7ZTevUKrs66CRtW9K37tGI5Gv1BIm0icmwwRWnScPvM+Ck/3nHFCFrAhW2Ch8m9EKK4gCchVU+D1
y+TZ50jwVvHEN+hZ40j6g1K9pjfkZylBrXKExCaSxTO6+66371A9m7bczdVWdYviMpmesUCQ6rr1
YIJm8gele4snDHOVRsfXTXm6gywJf2wqG2DcbuQZLYX2hpRLvnMrX7a3UJYemYS0Akz4JmLQjrGc
ImMk51JKowoMBJkgKLflCb2SLqDj70SzypLT3Qnzsj0ClbRVL+R8UeEObsxObtMlgCxjVW1ZYPx2
yQsMzQlitezpge7Zm56s9MZ/sfi1gXR7IPUNMChO8RiJVUeMv4L45v45BPdzRos3Zf0ot+r+5H/E
ZeUPPKUEab6koksjCqdrGi/F2hmPo7NA4OxHp1pOo5cjmsclrWZtrZqq16L7Z3+4erncqJqEat5Y
Zs3NpwIUDch+AcWWpzfc74UW0R8/OS/2OwIzLEJmHIqdIBR2RSFIgypk2xf1+r9UmnM6kcChlTyV
tCFRRHHB9DpdTm9fQJ15h2PseE1SWy+fNTmIX6CVwYKW7S+n3WkMXn2GhIZ/hkRc6sC9eZTEe/J3
AuX2Cfj/xOmV98YhuqhniVAqEob5rlEoHrawugvzIamFOxHu1JMhZ/+UwiKw4qr4KX6MB4Onqte8
/2whHcd93FEUs7lKECxfKeB22ZcgSjOj29asnwb3SUdK2ft+L1HCFYRnF2HwNBs/03AUj0idP3Ei
nghAZ2vaoF5rg4Vp2lKlXEFo4RohGp0m6vFCR93qgvoNYNQpee4jGShMx7gx1UdSsq1d3qfpeiGc
E9B8qfSODJBfqVhRgZyr3I+AMlnoG8YPGwrgMAUAaPKmQC3G5pohwRwKGzHPIXg9hmTNOl58HEkv
MPUwa3Ro+mcQC5RTqxFednF6io+zIUp7yxAfQVCvayzJcFKH1RqkCNcv++2+y2sa4wqm8lp9anrm
Bd3oGgXiAukH9ks38geQFsSWknUlPEjuUOjIokk36lplEqNZi30hoPAxys3We5vEaTfJo0smgsuw
Parsk6eb2yuS83j3uTZ9bDavYknW8Y3q/UBFMJ6anXuipCM3S+UCCcMTn/UnszKFFrvVUIOYEELp
8vq6chyhTjowIVW2F1uHTxKJiiEWqB4r8MHoQOH7QsV525pD0s0IaX6w6bSPBxcjmbmzrZnMZy25
ESP21w6r4PJgJ0NyV4wi8BOsrLcStyc/oIG1ABIaTeSFLInYr6q4DCmxHKGwQAfn9bFsw6Uh3B6k
2Jn16bH6m3N3nH1tvimnlQ+GVC6dT1jOZOGGndK4SXlVN/r5BiGPvFUKIhPk3r+Rh2amAIoaPLH1
OsYHKNIpgWCymclTux4edMNMyFXfYPsUfqUBov8Hi5boJyuki9FOV5Cu+GDOdw6fQZX7CpxHtg2J
gSljq3U09v0FkkHQ+uJH1eVW9aXNTYJkAeynyHwdzrZerlGJIfwx0Q/eWJfZvf20K+mDgA0egJaZ
bZUdakFEwqdrdWzsxu+Kkw8Uo6nBXXYZF6+HcejyDBAhDgUe24sEVf6mAgvDfFOHhhNRhlaZ7a+T
NA5uyyEOYHnzkNcqhRycCGOAi+2QmnEeFvozEflS7vUbJ9X+9pxjZuxaQ4F9YHo9pwCB/CiDZ67N
1tkz6W4tkB4gcI+6UGOWkCiBjF+Z0NKI0tf7IJr05eoeZmJMxB2X52LBG7IPFEo9ScyGkVh5uddg
KX2TM4A3ha6TPTl2IpRdxFX8iZARfmGoL+DIm5Eml+0k6j7sJndFm2tZggCRDSQUuGTc4hRCMOn0
0A32LcioYv55Xosd1YdQMCJyC7+GTR38jn/arMgj73Y42FcZOTI+5klgt339praXg3vAdGW5rsxE
79ignGy4lOMJ/pkR7AWNIaik4gu8KVGFxY8lZ+cd952S/jp9xTLNELvM8IXmnVRYElTQcO6TjnsO
ZCXPqQQ56HSVdcML4Hi2Mo8nyqh8tI97MIwchoSrqEXmXg8Kgj5nb3ViaVLjP0c9xk9/vNLdjNjb
cpQhLboviT9e1P7IP2PSIc91rAmhrIudSPBEDmVMNvPThIGzjNV5DiJDPHrNHeYL3+KKKINoUett
SbsdBpJd9qVE8AfnNkN8YdRNoQmfaGTlGCBleZxCos3EESvLUlbh9SzhdngRUJwEdj++u0Wla6Fg
/pkaQCFB3VuYSwXVBRaQCQ6eVaa286FGSy+JGT4GJLKg0MRtIFi7t2y4yBPIj96nVpntEEsZQAuS
iTRq+gUOTvm+goBAu5v6/GTpoqMBuKnkYhDhILSB/hrR1NSMSbBZYV7zTv71tG2M0DnwSywWw8/X
pebEz0eqGru5KR6/Q6ZlrCLWbo/eOwC05F5GmMDyvakwj8OLgp+KpuUrdkcWdOGu8VzjjFp/4egW
MIX0JIBqFOnl9teT2AOb7jZkqIUcoPLXu7U1xfyrv23A0ECdouPXwKWeLS/RjzAdHNde0pNV++9d
OHsNO8nQ6/woAV8+QU8ym1Klq7XzqMEfJz0e2xuEASHGQMGInC0tZc2HcdCB4NQXOwMZQlW5TvUy
X6tn4PPuv8Tqyy07WE3vBOalP3WZDxNtN4y6BJMovJPj2sysEYt4mFautkFfz9m2J8MhWKqfj6mS
IkEr+IgIud4z2FiLpZ3UvgsBll8Ldj4zMMbAUpDNbGv3qLJ3f5U4i0VRFWG1y9DTFv4sCzfNQS56
PCiVcr52NI5FVF7b+jwjF1mnhONXQ62Gl59X4XzwisCu56x3AoEbAv7ADuJer7ZhXipdIg1w7UZb
2F7v6F/u4z2U60nXNajBeoKuw79mf785lDzoyk6Hq7uHWUcRVMlglejzB4iRjT1eUePUYRKppdL7
qLOCFgs1wiC7Ip4ldFg+x2V7Y/5lvfEpeTkgrSUTcSSN3UmNixAaRXxNgWO3HU0At3wlkzzj25N8
WtkNWLbfQOkSA0tuUAChtClNy+QWMyJ6VysSQRlOEvFHdXaurUQmjPR5M3sAAuYP4TBzXGIWDjzZ
XJ85c5uQNhI6kgroWHqtWnIpgxsRTtBFxb0HMkZ3DSpi1R8h2kWtgqI3pfznxVQAegXynsK2W+fz
fnag81jBFJlp6XWfYNDVnwR4/oZmqIqIteojG9ZSfxudqjnz9otZ06/ySPdTHNXvyjt9Egwi4dS/
hFBT29wHKn1PJI0RP3jOC4MtX6SoCVQsNJDpnpB+az8X38QnXP1dUoVtnJt9GTXZw7YcdEeKD0mC
nZ7I4Oes3UhxTKCNz9RFd342CKWukxjdAh5sGL48u8qkOk2iB5DWzEiwa5hG17vw4Bv2wduQK5yD
6WhavCWbdYnABKoOaQy8qKTXYPRd/A/Q3JGCoBf2nb3O2jLiBz+BmxKxEHUnAsOGwvqyb5VQNgBq
MgibG00uzGBh504LidcBodkzE2qvWDxLqm0F2vSZSch1kI9pGYpddbAZfStVx8TGk67iKPmP61d/
90heUXgQzgMrpyY2R1znzlqy/SohfOhPTyv4H9UL6UGURBBfh2Xsby0N24ODSLuDeHfveAZvqcbh
XKQ0tiy11syBwnkHG7+zHQdFmxuH8ZGe5DzpW/dKTUqpu4mIAXjmFi9qwtPPDEVrEBPc+f9b7tGd
OX+2fn4BfF6dvdEGAY6U0ZntZpXvO2tp80c4mfUS9gyodxWUqQ81Scd3+Tw9H/fCKb51n3gZFnwO
EmeYZdAFzGlplqe/TxbWRPA12M/jX6oZN4ZzzrwEIFQapePeqETIDmITvxVUYjqjcrXcuRraxIQH
w9eqQKmgVzNoSqBi/GW8enkHr0nLiafdoN7rordvllxv15aCj5DfMjH3UWNA2cT6QzED5vgM8e+w
+M8nVCLH1ljQX/VqrYINNGWJdXDNxmKOQt9VnlSuZah4Teqf4p/vfIBJ8drGM5Nblv3TN82g/4D6
1QqnqzhC6ZiFg4bForE/hGT27OuDzsr9yvXIotyx52QGlF88sacpbCdtcR4A43HzvM5cUV57jJjO
cBbEEuMvIFlX41drTl7baljnYICwJ1D6S4EYPKnKBWVlI1xKAudeiJHTZYCRBtQwZPc7HPlYWJVW
L3saC0JINSv4/86fHIa6uJY9VCgbYqGAUgPRfUMP6Jt32HqMLLtosYRPI2fEucBNexx9ddKwgN0t
idOkGXaBLGlczhFIHymCmGnomWR4xcFl7Hh0IBRWb+r9XtL1ZJF97w0/F3z2Ddv3fhZyOou8eW4m
UWIVPaZf0aHspzW4PKJKMVem+2IbBi1Ve6bTUIK2MYrGgF8UU2lHP0mGVTeqqzRpKvmRltoas2ma
m/HEMs/IABGJypOg8/3vzHLh6wXU0tt+D/jkJQIpPfEDr/rWS8srFqswctOBTRmQ+dTN3zp/62rd
mPFUGbJ8rQuzUWpW9f/9SouY2II4tBULL97W0BOt92yrWPCxDlSYM+BjBnqjpmb42XBbSxaaI0Qd
sLFieKiO+oWonIG8fXqHEUzPD3VrRu6G4+yu0vbiAP7c3ngwrRlcU4LYBqa6B5U5IG4BxN3Q0+TJ
FyewSQkbEO1XBwAz7PCZxn02/lznn9+cdaqSY8ZN87wBJ2qFcmrWS7DX7h3QXR4OMfvP4NkPA81j
8DkX0BSKSH51Z7kyKW/Il8XH4QifdrEZ+X2FBDO+yQ8DFT6AA1dWrY0o3RtcPuSjYKmJFNqLO4fo
QZdhEjbJd0jU2UW9P1vRNwdUe3tHV4UwmdUFDyN2Loq8MCZdyFrdOnmCxO+sFKQxlVB00a8wWIQE
6JQnXu8iCsTUOa090zo+bdEr/jOrZGERd2/xVUN3F6Fz1dis+RdD7WjqtmlLj7uW3x2DLbMgnCdp
AUXgTpzCm+NnaDBXOCvYieKxmrW4pcNHwlTDqEcf/1X8t+jdbJlVe/IqGWzz0XprDMfspOaZ13hA
zdclIq6Tory++F3K/dMpOKGpGNnd4tgGfiAFy7XcQAT5tZLOP7mKpEXCaj7YGqQ9FwabCW8Ih3EZ
YB3ZRjOlfX7II7UbiIglPb6sLcOxadAGe0Vs2aJypyQ7jklR53EAQtnl4sevCJ9lCre8ys0xq62I
9ksyRU5JTeIzaP1Cu0RRJToiNTMqaeDOjwIiE3bvlYkLS3WmNeaMJJWzvg04M/T8Vf06AW5sCFrF
9cOMs3tC00Qkrt2JxSaLlswkb3HeCm1kNa8SrVUn8L2+6RLqFpCKPWWt/TA2xJHi6avoHnwmeJHI
k37eDsc3pYoCSPXAKI7WlIylm4dr9Cgu2kOwNTCo+r4ndWkxSTvhsnakyxLN7+9ZMhdG55tzYgh9
WL0Y65I3FG7rGDRhp9t2tFoPJ43VkayIaywwxAU5pj9qLQgAnJF5zPzzqWaHjXPTCDhYnO/Zmfb2
3MPBohmqijNCRfGgMP3wjUACbEPnRkBffjG4uJMeUpBppfHDG4G8aCPYYukr/1SGet38sY7tXXdu
14iugdVTNeSx0NJGk6vFUSgBmEKZXtAIGjZvRO5IeUKLNgE1PbHMAmK/IySWKEnKYTCHV00Tpci2
4ArWDxAgrMSmx5+azG2kGHhEM5WU7TNHWJApqHT/9Z55TV/sOiRuiK1SjfevSroaD12X9t7/2C/n
RcTqdDpsHw29IUSdP/IkvZw7SN6SobWaor88z2eXAw2MCiexiah7fCTAyuJDnNiRPIH53BlPHiTv
vuies+nxgtqmw89YClV4RIi4RwiLf4jHbA9HKNZy9RlKpfcQa+ltP2IXuv32uPYxlkIFZyKjL8Ya
B+VTh+hxDFccZwYYFnQhpOxeY5DZ6U4ejiFYKVtYIRrey33mamocmFu83EsbGL9DWRjW9i0vADWS
qv3SCWf00zQB/F3ZvS6VE2/DCM55xOtaLEYIPH9HHzUMyd/SLti5poTT2WVHoprHoVB7Y1JlVTZJ
pdf63273iEw5bEzVSgn02xEIITDHDDmGER65dSuwShSXlBZzLlFAaHGozJ9d+7poasZSPND7kagK
vLcgxlka9t1jJ+hQi17vwLIT0qRB/xkcFCNpU8l98uHfRKF6XMOdveMQlOYaNE4CJFUJEoj5Eogx
5bXqPpzlfwmuVO+PvzUCrxpgUy8xLUeFmy+bFJrB5p0ejFYXOll66iotCoyjzXBZmXYL18KspDqA
jwSkLNDJEsjHH36a9a2nSuxr75k8s6i9Y3HtBobob8YnOIQaCioWJiD2K22V052r5z0+VbiAse4I
LqcGV4L+NN+ZjFJ8RmfpsPHTsuJVlzu8oE+H0oDn0jCFMieGRWQtGKK0DC0yYMidfT9KWg0wyBP9
E1oRMGkaMDOPTer0CHxo+OHSkQsxZwMPMvtaBeqpxYGMYfoCfXhIVmBzre/WQdPvGznZ/l51+sGK
TQzyJnN6Ar7kIG5F/vzN8QlBaWgfhaBTc7+n4jTNF58Fulruh8J21TVhFm1RON/LROouFJ+DDM16
Adu4dd1Brym5tgxUFC4mvkVKsJRwVgiLTsZdog2IJEWVPOqzpeNaxDSO5GwDJNNDCc1sT67JKqiH
it8vfmmHRxUXycQUQNHkhS20WGqyda8JgOLcPs3B5Bq/v/W5E2YflHrNROEbdyf0LOF0rCKynhIY
4SBxkQhjs2H/Zppomd5VTPFijIu0k7jO5E66xuMrfRt1JC8fbCE/nVZsb20XPeTH4Hd435XekVVD
Uw2hb0+m45KK236fyMJMwBwEeBWNeDDil97vt324sG4gcVrj2cJEbZro+BgkC+ZaSDFDJCx61GpA
iDH5SNRRn+90PIgAeGpNnkQUh0YlbXGgHF5KIusbA+nulM0bIHL9XktF1paaE+aS/g3qkw+dnJTG
wm77Uoydoto/UvKH+AzFDTqUDbAsw9SINgFVuVvqFSTMKOQSpE52gQDlRmlu/vYRtWL7lanrfUZt
7/DE9vqH/Tbw1mBGDryl96MVVxk6xR270Z1uUbeskOhUsuFWlSXejQ1iuRsNNEjDHomXHEbNKUja
6+FRHg4AN4yu/tZ6QvIvhL+r+FlWIgmYdLJHORuarNEOnnq6Mf6l+PVemJmQTaFCw7uDYZpQDBuO
lg0904+DdJXl97AweZUZ64eTG6uXcQ7k2UykF/eztoS+8bcryecFndw3cxsYJEClhmNV9NPp+B4j
zebwgQf9hn6y3RatZVAflXYTn31QniQfE6pHari6CvIogzEnudAQF1vuY3Osohv7NUKFhAjSj4EN
f4uE6gBgP5Few6K6SXNsJOnKyxjGxXmv0Z/A1EYTMfDlxLQJ7J4gHCgTYPqqq6HEcPWF5C8DHLJ3
Y7Uwh3JjJVb9dobbjJlVp+Za1Xjm6rGjpN6nPS/8tg/dYbsdEGENdN4s3GUyOQQRBIfhrABZ+Ul1
2DU3hhthjUKFui92nuf/KJ5lZbLdeMtl1War/1e9R3aHi88s6Q4Qkg6+l2edIOev5HFyJGbPDSg9
afS88Z/DPI5krfIqMGobxAeCoRfZZ95y/UnbZTCeEKUdhV7nI+vJUOE549YaXSGewegYxtwOQ3W9
bHUJhvaGAc5hReNwECGkOx68F0hKUQGq6OfYh9vNMNJ6ECSWQMc3USqTyVmf91s4DmsmKhWUT/Fe
0AHNZtliZMJR6NUOJmVxMmvgBxaKcS/Ig5v1Vdw7jqKtgpYQCPo3LmR/dmhsfBaRMaMKwxlbKHEz
iJfQWRUoVB1xXOdTzVVb7csJp3U/ENwUz4nfT4LIIpxgIYTQnKAJrB0OaC4uh9SSpdDRYjHH/NB5
BLF8fYMpVBZM/52cq+8Whr8vnjUOB6rkdqTeXwrLJywAwzPJup8drwdI4sQ/PxYAjIEKhTL7PfBW
5MgGO6DIxE21uVIiGtStMfYrzJyV0X1FNQb/WgKBLNLr9FM7ghXEMbkwxFukRUR8aBppoyiDTckX
tUfkp6TXN01lkPhgsd6Gw0Z+SSnyEqStjBpnJBTwCuc5iahnTDT9MgQF5POQlA+bPAgtHUU0qDGG
mHonDwwpUxPY2PLZRXpARfYS7IkxIGYi4Q195brypfSPABfUPRW/ZB+NYlAGLp7WI/vzSDsQVtGZ
ngtF6vGq864/wkXiaLLzEqV32on/U9OsY2XjiAWWokaiaUrIFUUwPo7XSZjtInXiR7O/14DR0pWd
u8vobdxTXVS2H63Ou/jYXWtStsRUosAUsnuVsVy8K7hOVQLYRlFt9uOjDsLp9/GnAu5q0XpZnhUy
vhO9jB5wlxvbvycZis8UN4L82XJLLmhtzPzaww2GseVRR5HlbokDLX/igoUgmpDR40QCOXBlAqdr
SFsk1UsJLtdTK6WXPlks+wCes7ty/19QTNmhtSpT7dJ2jgwiMKPPr7vVj63Isg6+8XlrvK+ri14Q
YKWBxmoGaEJ5EOQkub0+I+KibtDcF+XKlKjHXF/bpl0zIDoNnLmNyv4OKYcynSOvnlXUEACKXu2p
1gH3su+zj3Ds+GUpb7ACyC22jMSyE6dVBvOIBMJedHHYMmCh/Gba68AWmYk/vUTXcjUxDPZg8H/U
cb7Z0STFXZdVVd2jD5ph/M3CYsGsg/x25m/9CLijzcInnTI4cwWBANTxkSqhqnLyMTRM9cxSc8NI
r8zDHm0iIZ3+/gv3TK3hjgE9pzg6VZINgQqUd9Kc7WWxntgu5WBUiZgWU20zmRJB/kHmT+BTQuBL
wfY4xYiYDYS9PyeNbgyw78No9xw6uWeF6CcUR1VCmCsxmPlhYtnqnvSXiMZNsOnuWG5mpHbHshr3
vZiK7bxKd+gESp4dAZZ+GJBe6ZGX2X0OEEmbTdeu36BHOsPhWq/hskWmTOmEjf4X+2exc+Knxx83
bO4YI80zbJAjCKFvG1icP9ZrrRM/5v1F1pH2xExzj5at2YgLUcijmsl47hPQGN6hACzhB81jAldV
JAi0E/5BwFjsm9vLqd887xBSd91/3hIsPQaLTVYtLf6iXzIvn3KDYva1Y0OnT10Qk2WaFED59yYg
47PNEupuLWx+WDOTB9EW1BC9Umga6/4dZWT1r5Hzo1ORcO1TYt57Yjb/H1S+1p86c/IP56XuSxlv
R9r0aEAs3ijeY99224rAmKcLj8xUeSULvUE7fAs5JNMqcIY84BE3N3llIoFSJzuWrsgYujI6Uf1Z
MQkWdP0yiOm8RkadBXpZH9FtIHUGbb0Qz48N/usd3VC5jMGNN2yYRG6z7FAVDt2189sSuMHKFuGP
Qraj1TM9iUn0qI/Snne6l9OWucYO6Y/injirBAgMRSMnL5ogLPk/OmGvi3r6pIpZwyJhziTZXN9U
v3NBKT/JSGby5TKIsL8+1I+WL06iGkL/6jjW6St9GwFfhj4WIhrhNVC7ryZATM7Q94xik66R0gB3
qZ52KO/s12czKrfq093BqeRZgmv3HylVpOiz42V9KKetY28fpNcYM3ykfCG1gVHvTN3Jc6Z4Zwrv
aNlfkkzIJDf1c6rI/TxRVoJWDKQF9ElG5s/8GacPfQsFYuCdXhGBI5SRIgW3Tx9GTHM2pt/fEdEY
bHI72RTJqGCDk96oAG1jWCBwdNmBVs7+SZ9Uox1mrz/dlwDJXLBJAhTlZW3Wb88UG3oyknKks3n8
uIjjvToabFT4FSZ0NpDrpNX2HEk2H366vc2PTGCg42y3/bngL4yp9TO85oFBhFEeluXGK43VVxRD
xQEinIlDW1IIy++aKzx/mA8OownhS/Og1bc5/sIwcqfNerQgCGvUozH5wRSqC4oiBxY97HmWiU2Y
B88iJvKlE1GatGblznE+LNej98bE+PhUnWD7+vcVYR7o5qVktdBWtHj0/zochkvq+Lo2NLO0YvdT
1sAjYZ+nm6/kDC76njz/uYZhMHO2nd8QMc+h86yokZ7lriQfk3YMf6KR61cq2C+VZBQ7C/b76qZH
66t/9ryYiqft/PYAXC8dHqvmN8g+h8R6k/aAZLyIlVDYVMlYBABaRrUkon0zyyQUJLIjpt7Vyf/i
uDijNEWWZnRfOn4Z50C3A/ZyyJ8g+ySGknFuO++iycXd2zk+HIl0Uail0Poye2O8DFj9Pqdwnk9W
fKAfdRzbaTyWfPfLaGsO7h31Topz3cNVAUc0TET9Aw9rCkV1nIR4hhJJ7R97Td4AvwFJhxYs8LGg
umFMz5JstU00IGr0caka0IEVkuDZ7cuNZAnrbfA543La2F3zlSWXjES8xYOcr9awplwtdQwUzeFK
cWTJ8fp5H/8lYm1FzN0t/hTj4t87KKSZlQKIcoIDxm/L8KzOxn9HPDeK9QjiRHdZzSdPLAF3TroL
vP0tK0VhjE9Jc4QKnaOe12zZ2YEtfaaat6Xfxxca6KpOd8gXzRNauEDt0fzlQ3MpmRC5i5/MN1SX
FbxpcNqbri5fMUEg3ZLCQr8SsVKL3u+fk4jVwFTsabx78Ym8MPxgudjhpjU2n9+VYoWe1QQhyJ7e
5BK5hd+HhT0/5AAQAfRUuGDFfAUHyNLjTp8ba6ClzMLRsDcPAtWs7KKpo/ug1QjqWJ35LQXosJLD
YZ8aQaJu/YccE/QGRWSBHaWGk7sWnfbdLGiRNTblJi8HQJjX1hdbhZUrhwte2MNHyPfTufm11tPn
azCcf9Bwd4EVDcYlSqZKO2t4hnykwfQcj8NhHhJyo6XrBhsHSBUS8/Npq3iBamqmdU4xHJmx4TUG
yRLYfDrIgQZPpi7iw9xKlhaHaXXPLk9fjLtoK+z5hAad64zOrENfahbxJDXnTPYramiWdDRJRO87
goQlphyXWcy8eTL3pP1FX17LTcLrscRpr2qEWeYsPyp2LaRmDoMSJAdLY8mTxWpiPx1r9OJ9r6pT
+HjlNHOuujbqTw4JBwyB2eyPb96pwsiKS/siEwFl7fOHlkOqiaZgLBXwoByi1PhdqEkThqaYz9Cx
SvobmOjawYxs16w47jAm2++Cqr/XccB4oI6Ic2sMktezVVhv1xoDcInt0vu7Smicqi+4YwQ9sz0L
6Pqvmd8Xp3hZ38Rwj8LUrtGiAomE9XSetmn9DHvHHW7Pp3c+3ckd10eSb2n22EWso/4QOvjFDWun
8pV1xIzuqR2TddX2BCMB6+5PSITDCaefTdi+s28hVZIp9Y2XrRfd3wlStTIKWbp4uRbEyLyH1mk5
2lS6Vv4a2VWy/oXsRIH5I3ggTdhGh0GpGSUfKu1sdZd1+bn3LX9qfZAR3Rr6qaS+Mza2Eo8rShhn
2cW51QcfO9Bl5rEkNT+NO1/5Aksd2LE2AOCwH7LEFGKtvfcSJz/WUk9wxDhE56MyIvQiEdNk6vbR
FanDu3CLDefEVUOaXM7E9sbFM+fmnyLewWKSeSaaRtJtaaPDjVGcTJ8rFLZek7twAJv/PsJUNvm5
wNioy6pZkkhfVVpn3GC8tiIe1LtA65KS9+1LDWMnkw7GbG8miFIVUhA3CbTvz2vhy4MaajCuulZU
AvOr1fwEG78fAS52S/MitOgDSY3C90OFy5zHesDUhOmZAfQWkBaartRM6HYaXZfwsIeeTdDfvfij
a1jH1zLAeHt1rYNJCGXpD6v9q1SXLptUfMNRt+P/2DEdD1bQlW0ZrYChcGx7wYmRm3XxL3xVXVFR
Djrtkzh3VOVVMQa9VOkW5RJGEWzCTbPgYi4m8SqnPd0YKKpQPN6zZz1rb++r00DXOQMz0Iq4LDfD
DbAdxG4tY4wem0nbyYUlJ1g5S9mz8F8V72eAIFFvnL6DDTOM8uYjpazV4FYUHtIxJJnXrLIssfbt
KqFu58Cia7Jzt9ebtUAXJDdAyDHcGHgVtao+vO3jUuAsZ049+hrdp2gX57ksDGiEsrUn2hjuN5qs
FVZovWL0867TiEPR6jTv+bK7fdPtHDlMnrc75GrsYsY/+zf5NFMmsc/KTVI/SIeQlLT8neLoUNXy
KLfPvtDAjeG3hUOOZ2s9Itd5gf/owAry/3M+ogGWOfEXEgEDL+AXDrw1RvZr5l7UuEGiVEpNo/sd
rTx+NwyXUqto5b5nt7048KZ9LAFNJmlPx72mWvUn4F1CATMk/iQb09x5WngofSFw55a4vV/UbPEF
85p/PKyhYi1g/YO8PMGohRsjIYe4GpnzrHqWI9XLleArY8Idec9W8zt3Ov46OpvGUVRIdtvfRmA+
eUeCokZcv7GhbrW0E8UGZrB9zZjqQHgfAZroLn3/3iRhokqyy3mxpuLiQSMc4maF9khDDZBD50Vh
WALtVomseBlZWy2eYogrEXauHTDTHrDjFqSjAUjpCJSPJ7OaViLYwpHKnogxMThtxnAbpANegtRh
GYYrrbGjqbiID8jac2nhF0B6EXWrMLqIkGMavbTDSO71/OZVm+qeowJpZ0kUe1BpQvkhCwHkW9+5
Ao1Cug/wN1BSaaluFpLWe3FTi0Cw8wWvv363v/zjD6lzC15CdKis14bbjyoSU1glUla+gkmJl2EE
XGG6fJK+iJ5zDB8Z0sGTQSGHG2V/25aIDPtHeAbgBjj/gY5Y4Dt1LzxPH8GxO5vDzoKRw8qc6Km3
ACkZxygpjHiUnKwBw/WVMNf5Ir8XtvEy9bavef4iYNCWy32MVN0NVp9hGdnaT2Fe5TIeAmrJsukK
xSkCSo+eZFUid8tGlbBE/Frk15b056QKviNRrdFNU2VBUyebjc5rkNsb3/icYR6NsRHEv1rFHn2K
n/ra7cM45OAbGTalUv1QHkqjry77Pj1OjSNHHLHJqDtc92TRCgibcthyne+y6Exo1eX6DVOALopE
2MPSnOlrNngp7iS7+jsT3hecM2SRA6KopaRz5+MPDdPIIxOB18a4DQQL8XsqvP+Gikjup8zYLE55
tYl/VwpRw+Aw5ceoQo5H4BecLHeJpn1B7HnheAXwH7AmJzOznbQRF7RpvhHEDyucRFP55vKe2dn/
eCRsPFqNzu3R85lyhHvKWHHQGs7tJ/zA6cWaUaaYjsK2hQULgxX2ltWczA1WZYCTAjskw04U+5C5
5/xMYELzHdF3YSYMlqvuHnz8hZIAy+PdIFJe6Hicge8W4thNlveJwjRgpz7nQi5+V+PP/x6QcZ5q
QLNvdBdcllKKbl/ymi6yAkRKpd8ZuJe0gN6tiSyLaM7x84Ff10YjlReASUthhc2THmucNJJF5i1v
SUiON45tZFXs8GmdXkZPkk5rrTkWZq33z/uA4Ek3YU77pBo3uvHLBavtSsuOJQMbPLEJpcgejQZW
h90NEDeuNFBxDQyHxRY5rsjVcFblemjRtXaX9n0eVFE1ThxH+SAq4jIqotZir/mEyHJvFcPBqwTT
AFht+rZpFTLHhW3J2EJSr2HwPzipuMtSFpWm+Eet4PSyXp2RhnDKeLhtrJXBonfextCyvAL5fAmo
v0MClhFQj/W8e+m6Uym1FsdIPNXOXrIVSYE+7ojkAui/dvz4DFFpLLSelwzCRMin+wHzipJvRu+d
bYkklwqhieneK3fvzBIIeldmE+daoS4tIz6pg/mHqAtarNWeVZ5b627sb0flzHiivX0SHkG+rJuL
18wKaf/Ide5vQ8mQ6YLAmyxR8oL3bruL0Bs0f7ZeCivnIVFgNaJFzy9aMUdKd60iznBg4MZ+zRu0
F2XDSBR+I+7ogfqpq97MgCMAnl+Awi0HkaRu4sTWA3dEthm3a5d1l277u8WNn5+vMctNQ1QNFdPx
mMHh+ss1Xncq4EfzN8r2bGmVs8d7ZiyhVF7BL3vicKNSznypiTV6/Ynr/RR32iKhxGpS7tsQJQ3P
5uPxmt83k/vnVEClAFVJ9SAo0oJXZ6c4835OdW8r4HWpEdHHD3CzOMrIchH0/1c8Kqn8sLU4wO0h
Pcem2uAyfn11WtcTAYtwggpjD0nmn0yQ8V//g0gLe4U+KMvl1kQpn/f4byVhNBTpNp7aKKZLwxXs
VuGijwO+uGWjOJdzMULHq6u+9mjG8jgyswFW0nIOpyEYcArc6ixZT40FooXZhw4teHwHbCWgdj9Y
qsnP+lNWsMyjt/xxcyrJeLTbqSjqVJIQhVxxFY82PdidDYPJ80c4L8fJ6HBol/ew/w5J1Q6SoNND
OC8jseUfIaG+uk6oBmc9nKEaLHc87i42ezjHrXHg8fe8xfOSedwiC+DN6LNXTxNxkh+4wEc/XGVU
gT2BYFalA+nNEK2Y1V8A5bsaKh9BVAOPXRdor8Rqde9sPmrfRD87jHORRfYxWwlAETaEcOJKyIKG
5Cwvnn8uIo2ztloJE+wkW8roQAUmOi/3l5NbuhQ0cOwUSQHjibFNrpz61xVhMJbyY9AU28SRdHJl
arREoxCbPsMKwvVPOVMR3VwOluHANkvhriedQpWzmyJZmavgo5DA27Fzc7L74F8ZokmE77RbbBfx
oNDbRxMO0u/1P2DCfi6RT5DHWDxuwvT9x+oQJfF/WPi1NkyHuSoVkRsBEtvgZ6TzqA/2kX2r4mgE
oCjI/jmtZJixbUaDvBGPfaPfy2NG0nnMcWyGHXnTj1/GMTKBd/fQAgtSgSIyXYG7h/acX/N9Y7mE
FQuY490wMcb3GECHbGp059uD7X4jaWeDi48FcxPqVgMeaGE1FcA1i+4i6MJlwj/29o5aQ6rsTpN3
q6gjlMfVDjpnF1uiza2rrVD9A9c0cd19Q5cA+N0uFCbsLVKyenh3UYSz9r2YqspAD3WEz0GSK5af
EpDyMrecI7/qVhgcZXqs0wYyXcbtzMVwjBeWxYuSom3c6DhjXOr1jOv/76KlOqSzrr+t4QZ+grUo
Wnwt6VxJFvR/DyE+K1RjaY4O9TGGdyi7q3ht9IpMjMFI5Aa5RR9heA/M5P+JyFJK5IcshLymyeXd
qApaWSwTBdrC6lxHVKOSWLyoVgH2UWUkFJyXHEp9yrkLuaspSc13SdsOl1V3xrdP9esFJqKqYYTP
UOhS31zCfZi+WsHTYL34l1JT4pPMYTMMqu9ze+VyK9VKye6d2cd7/tCPncusQmwy5s8MAmFYzZ6b
zTS+5sGPJrF95cZ1QFcXOOXZFRn88rAZ1weMV/+Ll+EpoXEj60ZJk4ygW0hu5zNtCFQabJD3rXJv
4bfqXQrzW105KrNe90zj3sXdUvlOypw72kcNUt4oKzEcVKo4GEo8JqGtn/CXz70GA1kIapcrgkvT
k6umR8N9i4ACcAHW6G46xSRVSFWA+EzVS52rSPi9pciusoyzQ0dZK9/KqK6ihwca2CEm8OlEzE8i
M0Tv3+pkSDjDucBXpjYn+A3Z8898qTmXpq3DAtqxBPaD5BmvyqOItLSqGcYid648pOOojSWykvxg
U8UNgfql4jganHf82eqAdwvcQGQgcscHHVIZrwXSVXpbENM74nFmAEvTtIlLmueww77KkpabArmu
OPusj0UM6KFbIQfLja9rwfympP6VzXy3MMDpY1fHLzvzh03hgXq0I7HFYujxAisoPVSHB7IYg3C1
uixNqdJo6gVG7C8UYwOP0HGF7TmVmoMG9mqI2qvydJQsH/0m7/uCfHxam85q1QLRoaYyPDlHOGP4
8Vx53Qe6ksJ2reQSM6uM2/ter1Chxpy8Me0yRG1o6AI+J7eq6Uxs11w1I783Z4TbO4bRpIJD97HG
uYDX5G956qh99xTyWFqj8N3iM1opyTHlZRiJx4GIeXMtPKftxrtpXK1OUOSFJU2zDlFNs5RKIC25
LLdrkKHAWzED7ne2t0WVORM9UkPMUWTQWu/jYTC65xXXq4SyHpMXs0QmJf/MTo/+v9g1TtEaTzwu
86akUwkRDdnETthdAnZfFQTqBtHDZwvdEm4zxfvHdNXJpNBHmor+6P6YQHjcq8/+d4Ul7h0LXRi4
Pz/3kn4ZRcwwPSpr9oaDFYKozYmhV0pYPU+Ef3HUVZW7DI/4WIBsz/6um70VHK0UkOQXy9GrQnj3
aDekId9NC0o5HcSf73sy/ns4NAJj3E7ggklD/xiN8TfhYPIRTvfHItoWpgS0ZAoOg4j3LOwdRgEp
7wmuY8iBqVVpDU3erpq9fnGa6RJT7gwJJ/B35m+P7itG6e+XCEqITuW0I1FUOz5McYhTTA3I7Hzt
AR/JiDsAfHSc08ENVM5umd25TYcMrdMK8gVg30p1nOZ2WJwxx29w/glPtioLlFOngwfGxo3DuqR6
xfe/2A/2MCJwxd4xdBU9TubuJK4rqdIdDHizFfLV/Bq3oQchYHPlkTkH32JTYif8wsLADeUylIuG
HUzgMSk2jLEXPQfSjkzBu12z3FxUzJzst8LHV/68g1Srrq86D8FJQ/sHjLoiSswZdWQm1E8IwcZ8
wWxv6NPyHakTuDgu6T8f/bn6Acf+qGTk0EkPixKdIHlouzb/WN5Dq6bEX559tM2dP8F9E3Ne7hNT
hiCJTjzfivAvd7ivqc06XU8btuNTvvg0Lm6vcMsx1ct/5HxzMs+3Dce12PZdv0PHTj9pAinA4+u2
S5vah6lyhg7iqwaPCtLkzEws3SXmsLBGGHJcFIVFbA30t2FyrerpzC9Zxld0KyLV7r0XVSfzBZQJ
6+wWAORdc2cHxHxT4WRT7dlxQSeV29psmH7mee61r8iR9ParQEMPpyU=
`protect end_protected
