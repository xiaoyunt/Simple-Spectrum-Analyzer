`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gl8oTb3yK39LjDQS0B4PYP+vte8cGiBpEmJ9JLxCkI04rBQJe5sCt4dvUGvg1Ga0GoPkN0BTvh6i
v1YMWuZiJg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LV5tnIhV6fXU4gAQOLXCxdxya9doivJt+Y+5yV24zJ1I56Mu4gOTYyKzdDBlwz49as5fPNOvHvtM
FEjflUU6R2Yh76tXBr2An7Tc7qdcv/WUX57JWpXSPQfxdtsoJzfNEA5lf9cFyHWa+eE27NH4fCIB
fHvZTqNYCqZpO8hMEWo=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CtefK+dE5tJYyIkOlXrI1GU3HbXkaFgSREpPJj1NZdNualyVqOHiPJK5xJ71xxO6zkXYtBYfzkxn
9Eqf7SpqFizTSC3YZVNAp0ix3wloJ2xu9/08YGAzwYtrD72s/REOd9GdOS5BW5KfXcLDWxJnWFK3
mjj+cPJfHeoGuNLu6gH6HD/lNP6geaOelYYVD/TVk4P/j6qWfCikFKKuomVo3jbRD7F7QdkJDCeh
d5Xc8VxEXSaKIjFRuMTWZtjAQjFH5UpSMVhxV/fXhvzSM6V5P4QZA+memX692B8GYsTFU76iMlss
d7ocDlaRWbY0BTXFb2HZNfGcl+sqYKs8PYn/UA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UTuJ2/FiXz7w8k47LqoJjpB8chaAWEBjYpgn4jj1PBd2l6Nj6avA0We0iYNi5AJkwcUofxaNsFtE
+sVWsmGPk/0vN5Q90wbwbfGu18ni9SqWiSNRSUzzfB9h0bol599BuMG2pbcdYlanUIn9oPi4ZKeJ
2M667aoQ2BTcU/o1U8nn5wuoiboeNIqzcJS0jj+j6J5UYz5aHgwMcFlCGUwSQuAp+2VIulW4T1IV
NW+4iXCF7wife+1/XS6RYcYu+n4km8U2A8z/nLIuNXSO1T2HaR6rR3YxTorPEFUQnfrre1FxRLzT
6pi4dXPFPyG1bXISdn2AleLyNN3VFQjTEgHwsA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FMUkchj5p9XvgJ9tR5grSuP9aw5xa30l1YgNWO9WvtYYjYtQnsPBns5ryDL+PXPqQYQ3i0NvbEVZ
mN4H44H269BdOgH+vRRI3SR79goz8NqADp1QSv06wD02bUASlMq9aM6Phdxmqoalzn7A7dWDa+nU
2QokmpYQQylaKE1ZbXrz6loBY1IeoaMxbsQcvxJcI2aG1HO9NfyR9d5i3K9UmO1t9jFA+8k+GsKj
kNnLxX6I0J9fN8wKc7D007S9DgoQs6+WuCL6CudeG25OH6Gy/uLkY2Udzdpodegx89FgRLo92dDh
+0eWKh3H5TN2vtQ9mtD1iH6zm1l1IqnYy2G06A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IjA88m1asiYMyCqMLSP/pVhA6mm9v8t5bFtEAMOvlQO8WTy5Vpca8kFPPuhuf6voqy+zwcLXRU9a
5UwLvCxgOEOo68GA3l4AR9WaPmcxPTPUwChO8zkHIDrS0eoDFMY1OTr1Lv8pbJknphtPExopREwk
KuHbtq4Mg3zw+se7q5E=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nZ0uDa4zhbQfoZoNpOAKrHOsOrOlSYjg5j1zWlifZ7mksZmmo1GUwbu4BrFKsE9nPAJUOa85AaS6
3sPqXGDLUL68TzDI06mN0/idhoIRBSJNinUfJpw4Ro9h/zNx1E//RfaHklSArW0rHrP6JnabQq/E
ywpKofyKtfWBjZrTJqD+xFD3BsXO9W35e9lAY/pTqzN6C7dC2o6xELYMw7a37e+7TEDqEPb1kk1i
VC/DX7v1veomIkT4wlTej+pa1pSQH6uN/huOhLuz4yEz/zZdnoDInKQyuWaZgdQV+2dfYBgbf+po
404pK0Ii/DBBTh6IKooZGzVmsyG/5MKNX6F9vw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1558288)
`protect data_block
8XHGIUnHoEXMsMueQ4/I+rdsBKO7j7VsaFwm96pNH5amFSr9U+1Y7JYBv5bTKhhKoH/xYISEYCab
uu1JGF+OfSunTx4va4WZ7YBt6rIx56kZ/AZVonKXpHSffww13yr4XaWH1TYKARvcTZ6LuafY32p7
HFYdQjpL5Ca8k4IrOjXKtHUb4zXHd6x/sPzSWDtWtjkAaAYLRWplhuahOuOANxdSLNcNVeRm4EgQ
bQakq0aciVFr7vQ1X13qxtO/fTbwNZnlN9Ogerlqbs1Owborlhd+XcLEYo0Cm7hSyFaOhPIGMVNQ
DEyNJwzhLi9hpeMIKESipIK2J+ZU9/NTcNpPqY0EUYEnZlcPXSjBlrq5ZfDzZB9ctRTRR0iwHKIE
d3Eq8Mt/53FJhouRbtF7EafrflsslfJ2iNminaMmrOKPfiCt7vUrHZuPJhpqRFp5YYuui1HWsDha
q6nICl7dXBMy3Bob+TcvPGaxl87IPReaj6mIvoRe0KAg7US0wLIVeT7z73WM2nnJ/9BZklx+A2uW
TKcek6ENsT2xxKJ8CW1ABi39nkPb8Ev4Xnd117OAQz5hbvw8Dlw1rygjn8gNJ/dWdOZ2DR/XawtZ
eBZ0PcR1Rx+pXvMQcbYquy5Ge/4iiV4k2Pp+LYYLpdpmStPr4Y39KqLJ8yHEOvjp2DWqXqwBMm26
ryQ0Emer0m3r7uiwtiWfTsOrlDmrzilbPgmOyNg+akjGJf3LiTirfz6dEuadfune1727MvpaepR8
NY87GahIXUa+RrHwyiz4G5jVst9tbSsfv+FB3Vi2aXbMW4HOjjs1P11YMGag/F7q58rX3swCCPHs
wVeTaky6E3kSoFoUM1G80/fhrFeQMVQDQs4xMMjjejzgpBLFf1IjxqFjA1rs6imIPzzahw1RJKPE
hW0j5Pjwmtu7Tyd+UUzr9MamG4FT2NOOuUwvhoFkiwDwotxFVMU0HtGh5okK9gSgepxYjYl7pDlV
WPrFWFJp21Le4lJZCNaXj1YtEMeCZ+VCOVBjBxNFn9z5pgsUXetYfz1IdwFkqQjUca617NXUHlmK
gK+NAsF6BZnfezOsmgNhO5F9KUSVsGhA2tvFOGhrFoe1vtHMCsvG4956Eua4F/tMG6kFFcVHX9bh
tfdFyqXGARBiBkQpYUjHn/Nb9d2c9+Fw24S1GcaKnsfwRgckDQ1qqAy1eRoy8EHo5JYnPxZdYPlR
c1YV4IbxXiL+yGhX99NHdSJCShd31m2iifLPgUn5fGOmewe/reTBqyh8FMI3pesZzl62FHnV9g6/
qcMMiI9rEZXs7vMdu0TP3iWlJ/pw/nlonn2SUocVw6VCIJS2U8YhG3Z7KO2b8srIUG9cyCvYGsvn
16WWD22Fb9NwfxFpCKaSraxzfXypc2lsGM9MuyQu7CVP7fNTA8csnB/2mPD/+2xCGYGCtvrKq9h8
SMAUaOddyJ25HLfQ5ZZhVhKGG3DWC4qqj4Fc9lVrqvWNSBvScZg3q3SyfZGajIXzCCaKsGzdxwTc
HeiAUfsFUu1kcEPXOMf8FgX6VZSI+cdgAgKRHpWjesRtOn6gp/H3j3PqqCbIvB78zT/mcreXazE6
GU1iaCia11KuAIQAZotlibXEGaueParqz/znABtHvrfuRMiGeobLR3PztcIFW6ix4uMbra/EvJcu
Id4r5yxkzvYrHcMg9RLOKqCIUeicS/87sHJprVfzIL9auD4EdPah0r4tpowcEh5q0mlfUz26L7JS
3yDdNyomPMVmxnr3eCZxCOyhv8wbfes72MpfDXLsyBqyXnGuQJRNsPURSivQLPnqk1hGIGq1cYK+
FaqijM8QzyrikdVEL0c+/OovEkUYFXapekP3qcynDu686puSdKUy3IlDu19zj6eaekITWBlWuwIt
fpyZQMwyP6OWgQqvFGRei66X2WeaSi/5N5vdl2gOs1ToKwtSEJaMrHl5p70XGg3jST16ShMtBoXD
3Rq8gE6QFmWCV9SefKM3TtWBT3PAnW8IlXkFRbNyUVox5Qb8DpWUcRjqFSfg3lc89OpaygTkTnqo
LHvqLeKfr0fXBd+UPoUjDsX8bwCqru9TAR8BCuFsRfjukDJIEQlUrfClh7k8UThr50r46WIoanDN
w6/JK6eQ8UMmhq5mrOO7Qef3Cw3VPds4ebmsbBiM0CMcAIv6xe11TJeYnyFqllcuG41y3bJLR7q0
4Kt9FoTTUfCPWIBh/kptT8pcrAEvFpiBu4wsWU/LtBswEbYWVP/VikRiZHoePMGBsHuWwnIFaxeL
HR+km48G4H6Jlh304hYhZviP+zpiqJpXJ/h13qjVQ5y3G3XR3X7N15jnNtet6nDypi2M514psoIE
s3eGpCgK909/wE2vGZyy7FjZkAukjbB/s60g+pbsteQ15BbjRAMf57hOSgUSKAOtyfd/gBWRNs2B
adYN7VWAJcQz4I3PtPaobCP6ecSpDF5LjjmbnG0gWyHH6qA66fHjG5/lBxRmGS8OlumlyGDSx71l
xtIPva1uK4lOBxOQBQyijifp2riqLOKyk6d1p7w13O1tmLcRmVPZmhi6htOqYiD+0v0inV7kohtF
H8WlAzM/Xfdg0KVGK5LOpq5tVjrUEOOgpX2ogxAdhzGLE7ZSyVOuxAMFGj9l0ydIWiCk7Q5eu4GM
thYeO7C1Z2Epsbr2whBysZ+9NA0uav3XMME3WYj4QK70myl61B2PLgFlNS0OhS5Gd29RmqRpnjv8
EKdwKqkERVvzCsE4HabCf+H+YRr18t9LllZlt9m7tRilrQTs74l40zTwOL6O6I8uwsDngIbWYbhe
lP2Ab5Up0WTdgTIJfIkhtRhIaOEAal+rqx57mwtXzJawvF9n59lsH2Bs529DHV8LtqN3963SPsqH
mi9YKN7GXHamdlA1wrwo+rNZFm1b7kFwjpWToewWpRWfkI/bi9qcDY8Kh3VEG2KRtopR5o0KJFrI
V35iXaLbghbZhr7xBH5h0De/Gb+n8RKbBavF2veIFbWuLqhmD+gr9cD7cx40tcvqGl3T5Jar0Bm4
Hbm3RXVHqjyeFETC6CeG+YOCwppACc4kKzx55BYinhcwao8A/LTUcWJqzXijOOw6BEhWgC56AMKo
MixwW3aK2QsDtxbbBVD+9UP0lBjUgf/6BHgLPQlEaR6K6RxI5xVAUBOtG/vM8OObZq+CUPVTrDs1
Dmr0GyxfvXzX1mDaIJI9lzejQaAh51o5iP611pjhBShDDFz27cHy/EGW+vOUPQysNsX5pYc/1TDO
JhlwYN16t1xyJcIUnLogtRXDmyHZpn+AUp0N5uw2K+KSYHH1kQLU8mAkmarnaKigPBpJ5tAA1pM1
MDj3G3Zpm4k3cbRhPacu3cBa5gVLEHCgN85ElTAdZZZcULWXWndBKH6Bs15RN2+LySm7ievELVqD
B/OZLP9ZUvaF74W7kPtM6M3XU5mNydh5nHLvCowRKSjsrfWLYEhX9BF0PU5tfP9+V8t4foTLYNY2
JMR6Pf6PtGc/S7v8QaJAdgF7KMkDAytzYU07IpHxFr4ZffpiDrJ25Ilu3gRP3XpTzk7FSXNR35IZ
4a+VJ6PD8RmK9toQv1dv4ca5Iqe4q+3y9K7YoMG69uGPL6Rz99T3fHvY4Xx6VFhT4iYZPcsBg+qI
CzZ60z6x/S7tCwsWbNiYvC5ADWctsq9HeIToz1f8PRL0fVphezpn85iT8x3itoEseiiTDhb1OG0r
2UvbSCmaOqcQZ1gLlf4/rjchkZ8EQ5WjdtWerhfhIDMTIUouryLwCKyqiA1bmMxM6jgtoM8uBwj5
6k0V4wnvCnKCaI/OqwWy3OAspxWBjv8tmpDmp7PKCDVjDjHcli7R/11L9Wx9/ODXF/qXHPvXuPbt
XCmDqbMX1t/3PnO/FWMYdIPbD4nj0sne0Kqv8/OEXz+23UhRoJqGINBWnusw4VJccT7NDQj2A/0H
/YuRSlI28qc7AjlmeZusmpWZHT3bxX59Ws/S1rkNhPGOlfGGFi+ZAZYhST0yt0YtvH/pPLkiYwkA
w/E30N3Jbyd6gXvMnR0GTub/Qy/Uf0g8rkjDFkNmeGaWJnRp19FvBot6WlO49wNuhRRmpc4vJYF1
9XdLf0GgpeE8gcxARh1ed4OS9d9yfi677jsvuio1fOqyqcRGZenaJdlGEMbWSXe7GPJWt2hhwipr
hPYH9MysMibTf+Dh+kzS9kgSq/Yzses2go0DE2azJNaRJsRC7cA6cHNc8b2YBA5b+qJm+23EgnAe
nD0oK99LGIms5W3eqNpZV6tyurmx2S4IdI1mlflES15+ol3hPtoh7nrt4p+5udMC/Vhvc0Wc26cf
PWbhb32eK40eQBP9gE4c9WHX/gUWplaHRmJeF+psNwSj7fBj6jIWBoZWAGE2QZRbn6EsA7+OgI5b
Bn2YLSLJpzI+VPxgG2bWhZwdxlojVQ5JWm1Ub5+mcU+6xNFP2SiWFVCpEoS5K8AN0JgYlCytaCZP
ZldSCJQDESZHdHg6/RPQUTZK2DAyb6Z4OnZveKXVmMNIm8CqJNr3elSa3J9ykpOxR/VhxPSR+jLR
4QAGFGYwm4VGKBqK4QHHDVulL411a/4Z4l2anruB6RFm2m2wAJjH+IKk8jWMLa1dTj5ByIL234VU
pmixopL2rf6YFi8312rZylL7hOl7BYSQ/djyPJN5234mPnK3wHSstytszV9xZVkqDEqrO++uyUoD
ACvC67rG3zj5nK8MahJ6Di4oZRmQncDnGtQSZV2j29INTBL6DzgOP+2pAVeEVeZtMcV68kNvkTq1
SzhXSzOCLobLMOuDqDdZWJi4VhzxYD78Bbhh/MU/HORgYXJeKNanOYHJKaZ/0wrGyy5+CsyzKqiE
MS8MLtu5TeTl9XL0Q8HVQ0Lt0c4kBrU2Ffd9N5iHOMFcF3vi8FbN27I6ufITTUXyvi3MNjYPARu3
yBwaM1KNHVKLE51HGm4dht/aBNd8KWen/sgJ5jiZCCZ/JZD6V0RnOQAVIOO5IoNVPPBPK4o157KV
6squmTBYueQLu8mKCIaoDcpY12QDWCRLf+g7owNg/MhiLCIvfiuIV6tPVbEQ0F0N7vRHG2EiKpW7
FvgEOkGZHbHvEHPH+IpyFRoYcnn50cuWKhXqDJ8xdWwHb/PcMFeVQZzOY2j9ilW7r5bDdKiNCRJc
Ywu80Nm/n0sNhTCi97W53cS8tYT/M4kd/nYCokGkpMQFHaRAISpYIufAVR82pq/BaGP+VKqvWoLE
x/ZwKmLRahQrlkrBrOHDBam3zmEYvJua2ZKnI/2DMhXo2YrCf+8bDvzWMwZSayVQXIjnIiH29vlY
5HCWZ8IO3/7Ik7UbS0F7tZh9jYR+vfFSGwRf2NJrXoztab4ffmsXxMc+ARJ6SMZNERkdEl4NqL+e
YUeyybN8MAidBl3mX5ZsBFEWP6TuLtF8VqDN0QcARF967fqdOHaHmx/RcQ8mjxacJ2TaSYwOaHM5
/vjgeZSrx3K4PV+HIceB9z4atjwIElFVDgucxxPL55FSdmewSpbECfgmekwW1Dd+IIhEwlC4/Q+g
rnr+XP6O7Hliqo1Uf5VOPsK6E53YAMZUjA2l8IAk5GnIH8y0IEJVRIxmChArO2dNp9PG4G4CHsoE
wLMMB+zx6XCo8Yhihc28O6NEw25Wi1qBeyyS3Hq5pm5H1wxlm0Ols4/s5eE98eG4RYa+vEWJDnUs
4hM9sRL81hR17AfRdm42MWgGCjqFiAs/OU19tQJZ0qan8aOo4VHkYkR90gE9LHVGskVaePCH1fno
n/n7CDRGZk//XbHqNknfVizs/6TV+fJn5yrwrpDTxBEUq0RtAOVQFUDf2sWkjij2Ed4VLlvY6tXj
gFWF7gkSz0fkf/ZzXgitPSfVtZSBrYWvCPRbHlzOK4k2yRnoSyzyVxUNa4WnO9wzjk6e1zkC+uAh
X7GTlBeitPkAZbQEqasxnOVP2CEnuxZx3XNgQ2fpMCgjTJUKlXRjSMqmtzD3d2dmHNYhZo/DEr34
tKqH2gMdYuQlYbO/YjqB8NjafaHGWjOGmE8sQFAJNBbFPf25HeGY8Tefx3NWDXDI22P+jXg8vNno
c6GRH75/55pC4OElsykaLqAHjrQBOd5DEdSYZRq64oF7i9yBj0kmEVi3GF0Yr44mcfpztndi9Kvf
c3QaqTkNMS0eg9yCQWOy6pWsY0QOE2AUtXWr8QWfiZIC61yryj9x3UJpmMKKbdI8mTfPzwZa3v+G
P8D7MKfIwe3gKf246PHMrYuc/S2YVnRGNWncYr6GeK0zzHyPUJnKQk9eNxwnlL86/nuiA0tqe5zJ
l4y7kuWQXZNevulGLBzplI9RwD8uy9iINwkG8w9ruJwrqD4G2U9ZDJMCArHTnK7cHOY4oe+gyyRK
zU51ng4igJyiZJEmnFLWT3DUHSyZ5m/wcMl+lHEUZhg46/ifS10Tg6AjNvDtbyLSzl6MR13wpP+2
p1fQ1Sngk6YqGOSTRASySlRnYEESmf4dHUlPGVl/m1MHgTs70ubcHfn0pHVdXEX093jCx9+xBm+f
tkEEqDX962FzX1+U7VFm9YwK+WZwpT1JrdavUeh0cesSMnH2nIsOHu3F7Ro4G5RojUJcPO8lnNzP
7zjpUhw8KMH7DC9NWjI/Eh1lZDznkU83DD3n/QzQgfprgxbo4jcL69tDU0Li6f3YHuCV9WotvBz+
MTB3gBW6sUM+u6lHvUnI88BIvj8Zo0JxY4PFU1l0EQTjMSElsXKMGgEGSrk9A5KZOEG5+iEz4uiQ
bS+y1BkIft1YB8pV3R4iARbpjGpwQnTlEQLJYDY5ZC3nZAEw8BS0VD8n6Ht18qvnYrI6n2+uPYgb
q74yUlZE/BkJbBDyvujfmFGgE7iye6DJF1XDBe6fvJyprN/qXCka3e79dPOw9W7JNYFb8rXDTbE7
fWd5MXaUclo2DW/Fa+P9mJxUGH55r/oWZnodKgO8dvP0LC56TsworeSPyC9JeSsIq/W1lYc+SpoH
uCJkI+NcYQWJckTv8QzgJpWXI1CdgzwPVQfcTod1Khhl5yjp3jptnu+GE0HtSYlaRuiSCKJDGjIt
+YBILhhd/YRz83oFOUAxTGuQ23EjXdkaIzrnm89zMHGT4PqFVGdgRLP98wrWq+CsKp8wc4OWvOGs
oRtCsY0V+7BhU8OE4FXw+v4ICXaY6S9D3oNQXl2BU8Mx5gAZI9p6F3rQ6wtvJjRv4mpiNcCly/4/
s8LrcKNizOeV1/kFrr920nPGqJ2PSc5amZ+PFxwZ8OV+SlSqUJ+Nn2URXcIfLfZjr5t3WY01jgB8
gWqV4QbED2PkH1xR9sOhVcN8I6EpGXyAAmwcczCZK3LQyJxsBYqd1Wg4SvKVYTFYJ/2qwoOIek/F
JZ6cgf20Ckvw7zfB73/2MZ1f6W1iF4Zm9sRhDrV7AQWiS4bqXlRaZrsWBfKuWLiV/CE7Zv6TzOdi
cAjejJ8O81qr8pVvyeO3i/BMYK09wTVq2HX50AsrKn5zH3wdjEiATs/OFYxcVPSKT4WaF9UqW0vH
LyC14pZlbmbAdQyKWE+UzJzDsOOyUajVqtZc53Fj7518OAxKL/0l8UaEmgBYWGn8+EIuSqd62prj
PQTSpuxepCABI8ChkbPZ0gG1oZTbycVb1ySj/n4zVcTgGjxXcu+OR1aMLASj3biudV+bcspssl/+
nr8xKmCa0pncV2HxQeLZnT11AhCL6SpHcuqagI1pQu9qBcxoINL1EdQN8wzFn1PDr4J2mW5WCvS/
5RRt7J68OjKUMK14RAV72Vg35FqwM2MOEuFv7nt1pkHgHwQ3WCtxp7BOp1dS+HPcK/KLXxrHMD1L
GJUI3W6NqSIeJfww2cVoODC5rvN82ibAOqhGm3rpnc4My97Da93t0udOej4DGo2HVZ/lvfpkODTe
CoQiPOQmkA0GdX/6X6dTfDTysC0iM1qWJwEGs9uJ59kiHnsbk+d86sLxWqWt9BN4tAVBUUj8f2Kq
8uBoqc0wOSP6FqODqPAdulwYOeLrYCYGsn741e5fWI1XKPA4I/gfeY2jTxCJpo2I2auNvQjRZiEZ
b05xjad8ZGDWV6e2Yb9fKC3MGDLon5qX6y1+m2UbDEJV1CgEIq5NjyxOxXXyjARRciVZAn4n+VuZ
764PvIyowjUW3YF6kRce2Nif1w6Lw+CURDlIiUPRjlaCk3Rb5L0pNC8ex3gEqYmuyIbsNL34Ir4K
VNpMK6ZZd7vYt9p6PbKn+KXQXx8nHKco+TR3P5TUpVGvrpbmRq7ucGcEukQqRGLcTPrlkNZ465z5
WQdvp84HxtRbpWQ4fL+Hs/reH6lkpNQv+zkN0QuumgrFZZsGdN3hZLWG33Bvowrs3y6+liaH4OJt
CPUz9SPyMqEfIHdtl5RhETRVAhiFaqcAznzu2VtcIxbmbw9AhcDZdI1fteLu8FWRivGevvQVksJd
dd5d+3Dj+hGQg/DTB3NXDCvXJZHk1krkrz9aM1xqSzYvU7ag/YitH/WH8xRXzhWpBGVrtgr5yWFM
RdxKxxwjgSiSLEuSUH0FvQBtSHjrCPE9pGBv3ZXjGkdMk8bcu7jDd5MGQCUSNazGm9+xEnLFr+PC
XiKLWuXgVMvKlc+Y9Uqunp1fXcZD7yTKRWGyjwlAxyPjO4TnDUZlnuOqPGyNtuCwNsP9pxv4sL7j
bEApL7cwrRoUar/DKZm3TuUNoWKljRAyynVh90u0o2ZS8y0mMNLYWbsoiURBl9YbMCFkLprM4fof
wRF6nryDgwyOcAn9sNK5MSVz2mudmNghntFM1oWt1D2XnlKIZPhZoCs23KBxOrho6M5kHrVShgqZ
lZ5Ro9+RUqaEXHGszp4ZO7zz2OTvHPN4Ls4w02cJsRbRcQuwserJCXLMkkHDOquF7nuLZS8mMb4M
DMT5gbz0KjtVr03tvXP3TcbDyBRN0QsRkdwV6Ndc5QB4L77wI3T+/j4Lx3AqQ7/mk9baEjdIyfB4
Uw717RiHbiwWvZu79pyXW66ZgRFA0sT/o2hdbBseVzyy02JCa44dksFdBSnoivkBhWhZMPPZ4Enp
+PD5K4ck7J1K/NrXGeNaRIUnFazFHKovGDR/dRwgLM0xfISqVe8bT/sVICc/8lR2KrQVckX98wv5
MG/8IFVOXUA2hmtaaX0NKmPtk5TC3kD2FtT6ZzPxdJVeb2C4vt2O95pHL9tEmkZoX9m3qNKMB9QB
izh4MIo6UeyVUN1gyu9W/AtCACxGmBmifEK7hjXGh1LTvx3tnD/CI8/yIBlgYSQcsauP0AotTMDR
QqS0VtgMfIdnZjcgUFQpt97cMtTeB0aNSEo5atII6zh2HApQa/wNnlGdq+MkLPQKjkdayU4Ggz66
W+Ml4SdFn1AFFMPbB13owBbBXyiH0aF/YhjHM/0uya3lQMROaie6kg2X4640mRK9Va4o4yO7eV7E
QovxWa4jxREIBS2bZq2OsadV8UlRcC3hFMGuV8vMtObQPUfZOX0YeDLCItTzVk2e9alDDz3Fx8kQ
cUnLF5RpwaBotEP73WIvVh3lhVjoRy8W3k2q36a+29cJzbVlwiAsf/bt7fZs/eqCYFzDwblC/Bzc
E+SGwmAzC2+/6pSzAItDQ2BttYQluBX1ORSgQVpgB+03SicLWAlgXaQV/P+rnet17D4QORzZr8Y5
0L5J2b7wjoeHzZEX6vJyBLkJKKbBhAJHeTwzjnw//BhB+DnPWKdVKGC3W9bSbKwHL2fAT7pKzFLV
Gn09WroGlNf831HHl6X6sNQKjR11YC6q2wovnPCJ+CTwCjQcJ4eSyzmKLoY9zvV0o5vJRqS+haj4
FIL3geoRXxgXO3el37fkbjti1AxOIZ+J8IuTPuRq3ud7UbpSLOl9BxWTrHONPRP2nba9EIfp2l5E
W7owm6ZDKNlGbg+2gkVx/jMaKzsq0GfOFI5XLsGnVxmscvmS76XhK2mJ7I9pMFsiXx1vD674nhhk
DMmYkheIcKVhsSRhwcT1pE3a7O9UxLk4hqJVtmJj0UKco/FpesVm8zSNC5xFc3XUL2SDdv0Jq3Tx
s1n0GMwoN4V+d+GUNI64Qb9FT9yGXlK8p0XW/eN55+dM98Fag5WAy2Hu44NHpohGU+MwCZpWGZZZ
1UOoQ5KHLAsffpjwSF0YlGMXq8n6gqgK6Xmm1QOBpLZ1jDCJEgzLi00c/N6BRV7Qkbc18nYgGLo2
z2+RHFp68R1uhkTmXQrwLYBhC27XaewBq39pEWACW3Y1IkNlC9gHRUy155BcUoEenSmbt2Zj8a5R
oMhr0fOoutHsYY5Kju6DpqaW8sIlE7VXF4vIOjc/9IiObF9W5+XXHpk1hS3D+Wg21T/oltsV0qYJ
xoO5tdFlQAocegS9GDPNQYu9Bg9bbBQfP+YBn3PZYu6muYVLdx104IMSatqY1LfmhpMKX+ObGpfG
MMKPwOTnZ5qJq0m5If6ZM+4l27tIxsgoknU7EQPiTWDNCGDD3998k1b8/BNpdkk6UBxxsefj2JMN
eARdhrxWNJvJf4YW4q73lcOJFLfMKRbwEC/0xevEtmEnxVptRjJ+ecX4cikuU7uOt6TMvKwJCG33
bJ10KuL6ECBkRTsXq6laDaByW6Z9sncANy+TY80PZeh7NwHBSZ5RJbtVSi+fF6MeWzbVgMEbw5TW
IAYSgZKT8JGzvA5xZs1SD4IyzKyt5xHqCgHPMd3ef5NRMlhNo/Q5xuWUWuCBfGatMxSkXhkL95wl
jjVgC89rl2HWBRpXsuuCb4CT0YwfYgj8wNruIVjaMSuCDEdbS2G8FQFtWkxc5a69lSRbqPk9wXOr
t/0NVM5d7YzRjT1BhmeuJ1PYa28lHtbdC4FyQzcckkYjGCAMb27IRo4zX2ytteAHLPvM1i7RlA/A
VO24vti6Zul/Qo0k8xWENNQSEsBfawg298czcTjhAZtxQHR9BxqV1F2xUmxkvyDmNvPDujmeNGXx
uL3EVxz8qhniVnEkcqHD6yWNCpx2qVuTgXFQbQAUzjd4hDiAd33RBQMJm5hqPNqOkKYiYrfBLXfn
Fxx01411r7IpiC0rvPbnVpmRMHXdytUL2JUQJO8WBAYbdXDq+blURK5Njsu1I+JJjDOILNg+lrZV
6EozXZzEX6HIvXGUt7P3WprFsNsN7RUw15FsiRzL67l+IVf7xDaPU1IifmfZ5LNTJzBMY2JJBK61
oWrq5MX28tYG57ZWoXBBxkMdYlIiqgv0NnXJrwm5sUHFvXlsaD3HXQcKaSVACGsE3VfaVOFrIvwJ
Wh58AKeberICzgC3eUgekazabXGJDdq7/PvTPM7/OQbnsj8hkWL/fqYT0dDHml2hm/IaIiMgD4uj
SBHMrdzvq38hnVlEa6gMfiweNxWwfdqil7Eal0ZwtJV+Sj9prgENkSDnZ4L2MpTfJDORcHuvnqvZ
ukJWyfTtbE3RLiK+ts4fb0bfAOGa2RCvS9Rwb7d+FOuXnDDj3Wb6AncJAGcbXWqZmoILHrPB1hzh
YsWg7ZM1dYkj+AhcKuUm0N7oAbVYtFObfJiVq+P8NITl43ZiPFYCQIOJ5JkZpTN7oKQxKzR6BVQD
KXzqXkOul7IK0SQgWSvJU7cALyAfw23jmCJmro7UqfixH7VYDvPGKkikKl86K0iHEPcLqZ3ImGFA
aM0hplsevk5PdSQqYjKJfr4oItuAy95OKKnEQLQh4uN9yyURq4U1MggzO8I17OUQ2fFZ73ydIJZw
WDsIOkGxQPLLANeV7Povb0ir2mNulpT+UvAupq5dHaKbfI2J4DwCbd1vOTykZA5F2Z9eIVlLTJXS
Smt4TFW5xB+N2haAMAjb60i3kSjjt9PERLLSj76sQDKUrfrrD1SdeNlSj3EsO7P11pkFCRisi+NL
xKMbrkNTMHdn8jsQE38hWM7WmsVmFGQlRmagw0cyrwOkr+RsdFB0Mvw5Cu2Mn498ER8PiNKRhF0F
fa6hbtVYhtK0snQMt7Yk4SXmtZ1PDm4qwjSGGllMH3Xk+7xBvj5Fjt9zexOBwCU3fwceCb0/rcne
TnEXE20w779ph9g1OIhDhjiVrsOjN0uafHAasNHKGx29YDBF+4BF9ea24qJekQ6nMzl7H2VWztR4
SiNKlMvS32A9ez3M2sM7/bWugsYwrsvTO11LGgfqhdXEe/hf7Zj3XK09bVhBvCD997NAxTEYEdX+
mn/QrvaovAXkBAgescJ8L4oL+2N47/pTUh6cMOlMkBtQi9vMZNXseECo8KYzPjdJEomgdpkLj6VU
LD9FLOrsC23+lbvsseAynohL9wzeAhwlxHYDwU622xlXdVgBTWT3N8aQTXrm/B9IRojff517XOwi
LHzK1XCX9fZceQdh6kd81tNHYqRheCxF79dVqk8h32eEnGe5kQDUJG4S2sENN13o/jvNeyY+GVKq
XN1NMXEmJjI0pr4u1oOBkf3C3B/VpZKe6bjT6kE5GBZCTF/Svf5dbxbhzKZoLB7KLqSVGTIMk1l6
NY5pW2VGpVKhCdQ3zTGkuHxDm2QoJ2EjKVneDIEEHaQMkgv5FvngMme3zfVQ75Ijjrcik8GNetar
07lJXpW554BLVhEL3t9UfRX/UG2MxC8BYmH9a2IGA+EFS9RsJrBmzGSg7AN6jnBCPruuOxB2FoAz
RvYqousacpCnvAFLGgGKwbjBcq3WoMUzNTHocQEMNpnIH//KfLWTNxZF7aUPuoN29ElC9Q+QkgBt
cL9cn/FMynmxsHb5XMTAzT8EbkWbHOECKbX9cWGPHf8AR+rIqBEMq6K1qW452lh6RnYYrq8In3+u
0XLYs8Cr6PyhTUhjo9XMKLsB9JymKTGLDa/slK6eJQZ3eoMQqmAq0SksD4uTd3eumk2PXMk+hcAp
9jxc3/Ig/V3jxnOSwYuYgV5PJfR7a/GdJJ66jUBXMCy52fZDFEL2qIbM6aiMel++j4G3zuBib6Jj
uDq2kkWun7Ibzv0Wa4qj0cv6h0U9SKo8PSnpFQvnb2/hd26NNOhrLL7e48m0Xuwk7ALhQc7L4Cl/
DYDEkzCxH+O9oadIUjKP/V/79HpWEktzi04Kxvr5jZlF5Of31Ae8W8daxW1KLQkzL9Aw4WBJEIuP
McyMrqjcdNyExHxBJCYt4tgCIyvqB7D3cDdYHJcVHV6QgAMkx3VRHhnT3i5Eneh+gSaYv9iQBqwo
whJCj3naglEM53rDJBeQvz73GDUwNp6aisvJor95GAEoM9lfai3exUch6bzsNYDfp/extVLAAg3T
BfW1iniqydGpiIfKH/yp5ZYjhxlXKoaFOkQLRkea9+dyq4kY6yGA29gIAHjA45oJr6cr9W9/aV6D
DeGTK5i03y37va1ql8frszCHSk1af0udkeVtiargFS4sM1m6+Vn39vqPrrJ7d6Ta5s55O25UjI7k
ExpJyYcZoN87zkwtGEH4pFuAa2ZAKRcNJTicJ1MeKW0aKkni5wPfCZDK8UIJtaQ+dn6U3ZGhPiDh
wBz84G+7ETBXfjoohndiful68n9uHFeNtEC7Qb4YGICYfd1Z97pjtw8XlxTLHNO5JXmsEGCWNLXG
UfIX296opsq/Dx7/Oa3jcFBXPNq/aTQn9dDAzV1sUuUa+Zqfe2Gu+SiSnHOllXkTHDlqX3hjDPyG
CkiuZJMEMtY3WUJ5/hw+H8JOtiIwehdfsc9MnUIdgLBtcqoicl4lXUgFQqB2Jgh77GBuq3BV3Tkc
O12po6SvpdsAvL562kC2CjsQ9vO8j3JJzrBNHZRT+IobcIVBzrmJwU5BarQRs5roPqwwkCSS8aC0
74KnwiCG2LQQSnNx+JUGDXxAgyfFZ52HsOmBhSdQ9/PQYvcSv1AnGzuD5MX0u20Nd8mBJsM/LhQB
GxRFt2Ya/y4Kq3v6FVh/BgcaNRrVousNOWC1HOU0CYHGd6rgxzVmEXvPbWNvdo2jf2nfedRryBoE
G7k5YB/1ymd9g1Hr+sz6KlAcIAnq3dwNac2NNtAYEXiQwEYASKhB0ufZ/DFNmfb/B1jyvG3f6AyN
6tJWheWcD9wfY+0nC8ES/eorMFU6PQgKPyyc6XRr8zko583EllIX0dSqFpXjhD7oPgmmAedeif7k
DNrdRL+bneF7MDrdEOFiRTWAgFcA4wJm8FeyxgiIF0YK9QAU0YfNcTpOcvz9Rz3wM+XsngRRWlZv
sn5f98mdVMRqZwxYbuj2ga/qU+/kF/wKhLlHUEEqChzHeOzGDDtG1ZEM65fBsW9LWeIrQv1ywJQI
xslo8IGJ42rZRb0kPGr16Yacb01jSc7uDMXQU2oUPUnuAzGDw4tPjHT0Zx3HA0UvrsYpfXRyNOFH
yFbZCX0odPBV95po58JN9l/HypWwsf0Nn7aC/DHRb2NR3Vt/ERFjxcl3exh+3AuZ8CZOa+Zew1i3
wBU/FdzFoT6x66fmy7Vdb3nfA0baI67MmA/jU/be5VYUYj2RJaCupUPhrwA4/2F7qcQnBKtkThf0
++qUUCojC1JIrVBsv9XIPjlhmbHRwBHtmC/ZaHPnFa8Nf9lOv/jgS3d7FOwLRi9RgtD2eQvI1shP
snpJDtZ8meU2I/H7sE4kGhn4MVd36yIGL571ApDuO0qoNFCpM5xXQ22EzlHwr9ZuJgujoNgC2YIO
H3RC8C0lHL4B/iqL4nyn2+u0r+tKykfcaKbe+Qmou1GSOYhn36ROCJjXR1tWwqgEu0I2APkYJGBh
qvFtYNggOBw2ErnEzMz5hZ1q7pE236OPjgjfTG/mkqFiMAEVghqFho/nk5/8+k80sTz+78sI78lx
eg+PexJtZof2Orc5yZkjIYB1/o7dwyOR/Au+iEWyH5cJt2sUBtWakbbofx/cdfE4QAiziVNxtdvQ
qDkycHjPNlconmtvz3Ixthst9Y8XPOyOiwKAdPDUjbcGP+2nIzq+kU/Ynxtc1WNq09IIx3s07lHh
xBs2Yp2GdWjyZRHypwv3dpAP/Ie5cAkPCxKxullp7nDz0krvezQp/X3dzPJ2rYjVf0x12sMNpKGs
SYoA5af1Jb4jgpGD4x9vnpIxiQMbJ6BngT5J5fTKBZYjzhMah998KWaMxXcnNyhyXdwsSfXcX8I5
zqySEnxLaKgOI+3TNTUiaFSw/vvQs8jW0HxBd5lzRTikwTwxauHJJjY3yhW4iFlzo1S0r9KsmVEI
hdPyWRpNSOOjx+rTTpRown1OrXKfT/F+HquIOVXL9cWAem3mju1+LOcjEN64bGkGjOtzMmy5XT35
gD3bA2lpFISDGFHpw3Ft0tvZRddAAgONgr/MFaB7s41jweOp5Dg/u/SheKspR6wbqllnO4Jz7ONz
EKho2HCeaPbeIPCx3Wuiq1ZMYsheUeQOzxBCnteA8jzdnOVL4jB/wdn0fyxkMq6syMhsZHe2jAtR
87d4wtV/GD+JC0MaG8VgsFHCmG5cc3R2ObuNaVrHgXO3Z9XBM2GLNJb/N+MhM1C7BpBGquVgEU/k
lsQbjObEAdL1Ah1af4Eka8jyb44gwcxyCnla9B0feXH0Od274KkqmEHYmUE5oy9H6z7SXsRToYmf
7LVP6lT7xdxonVnpxFmhUDn+5VpVP1b5OyPJI8BJh2waV/FrAGpBXfnx+ujrDGAQHn6vVoA3DiRY
uKMd4NB//9FNdvo+bfUqnSILBy3fqLrjeHwXgkRgvc5Sqv6omuePEq9c/FhUY9Bs3kdBrkKGbJ45
+zfmlx4eE9eRGKAJklHGszkxstnnv5y+kC1RCRNs0zvxwF20nmG2LuPAlEqpDO3wtNyVZzax+lVS
4sSLCWXPHT/G0jxK8cSiryBdThjj7JpQrDWm6msDq7t90SzVGCsywObgWxDYMMAZs80Cl3bLycVo
vEeMus3yk6ibXvvYqmKLlo8/rjpuBMHXrx/TrAgsoE785eYBK6gg0egu5LPOTbYT94fnagYK898b
lUNWvNqm9WqLp1MG5cBomxoR2ADiw4ekeJ2pMiVfkPzeqv1+XHC5LSwf6/IcAaHsNI5zydfKXi9N
o2Is/btm/8q33WMTtiFAJ2JgZY0jx+dXWGXPfRri87fGa8wiXeWuNhe3b4k0hbrZrW7jAOg858L0
ESeTkL8KovLPY6Plnmit5SzW4uI2zWluZ9fTTRLBAaOt1adDZVe0UpRWYoZGM0JBcP3Bc4L2uX9O
4Nsb96ZszJFQC0NLWjpeLWp9gaPrGbMdm0959L34YFhsAIgMYVPvf6Hk/o4KioDvxXddz0x5n4cI
mWsT+wB3jT5DSJLXV/5Ma0Nif38CuHaF5HL24VEAGZyUgzUtseq+I+A6IMYMgU+ZjqT/GiN678jT
M1STptFP5BQIFXNMT4bvRxvxvn2fxuyfzVt2TY5oLWkyDlZ/nW5GD98ZRmvTU3UaeDcz1w9uD/fg
Gb4HIpJkZxRuZHQB+vqr92xJOXTdaKdI2IxUGx9kBX2gUetapu53TsYbgyEIO5gG0IyNMayfh+ux
lgYWO55vV+L2GWa/eu9AzkYOKzhKbBl2mUwWtfFmz4Fg7wemopkh0GaAS+aevlpXDF4Zs1QDkPi+
SySFAX2NlQQpxr0Aqw+YUyym5bXlL4esw6PcpdkSZHel5RxPVcckEWPx7XMMt0VzoFjn3c+4gtoC
n6hsW61R7NlLFK2mjNRMTnQkSTn0pgt0LIss50XzWTCOAzP3pbTxk9bDvNMHjGD3no/FVEy4dp5r
Y/n4um+8dQf4U+NNXzxfozfWcAgyctdy36vOHjsWErobhd3hGM8FfVRhAXD8Sy6WBir8uB3+6CcX
mH3+2/Dc5Tbw4oP9FsTyrgsBWysBbPOTXivWOXF5g2nRa1olEWwF0cKl/wR8bBPFWgeQ7XL9enrV
KPiCMc6kyWVU6gfzKTve1DGLPBH19IR+0cu47bycGv0hqm2EU+UZR5AzhEyI3ytvDoS8EaqFy0rx
iAs3hdJH0xnd+BFyScwfWPdht83UF5qaNI6aSq4STn84IFh81JmlbpVNSUUZ3O0EpX8nIiyuZ+Gv
Y0Y4gH4Q8qItRD+6cqwW+0bQoDvWQMjXg0el5rseS4tzJF/rAvFs4x9f7y9hAuYJEElOihGQmrju
kkgXyQ5aBFk0j0Fe9sgZ9l8HfTYAp7Bb75Q7+ZResm7w7QUdKhsD3nCW3weSAVEvy/DNmZb7Ng9J
iKnqR9ydRdl1SyiUvoOVxgkVsehzAwzwsqzvqon5tlcKAJXIPDBqcPUuUMQcnGThA8Fhli1qGzyJ
A+8zinfP9RUNJF83HIQPAqDyZqo+JcsE+kw1I3FhdfBkkALsmuwXjln/mvEuIGKB7H1+aUdv2rUy
xj98WASDKe+9XfY6YWT/C2SiEsH5Cd9l3wI0OjOqz5Zxyq4O1mMGkXebBCISFXL1qdIhfxTF13cE
ydY3YA/6WN7dhsWNfUIEcWpekHwVJO/vq+OUi0/oPA57JH61LZBHRR7GRTyYaxyBMx5KK2YKgeH5
leaHjMEe71t9PBgx0taysTsI5+SaWy0mZLphaqC62fBLZYbn+bfWf2LrLp01/V5Kco1PJ1wA9At6
8dZUwWcGm9Qf4egP/Na7TkyfSKhKmbMeibxGkMr0OKjG1HGftvgBy+8dZsRxd2AdRyB+djGPEp7q
WUrSHM/LyGs1lM08ek6sWeYww0ujY68Wie/tMpUkXCbjzp37CVZEXC6Uk0xEEjfkgedlFEZQN2PZ
EpkqaVdWNYbn23bVe00GHDCVa5vXwSl2seKi3ZNC6/noF6XX+pDRgNP+hfv3LJ4Z+4uWmjpsO6/b
oP2lFw0+Iwi1LEfQtLGQE9guhT1puMqbmWm7GgrF9KUPKpT3htr7leLC6QSEx/m5YZganzA9aDB1
m6YZht9v0uSVBLVXceN9gC0XDWb4oc1N+ACml+7d0NMisArqVlWMRzUELwAoPwEqmIyIHUwulYkP
96zqPkWhU2S3qWleYH0yjQBo4RnF5zTjm8JoIfuO7JkKCbfPnS1QpC7yAlc46JBWBO+yghhflvDv
chETpRGQKQIEqei+yTIcBtBTa46a3um41E9gdd4VoKZC18ru8Zqa2Usrk+JWlT8hPm7tjnbegwV5
cMbgKIVSPrfnb+0G2+I0QD+JdcYysdpfubuiaAFFNU8iLIx964bmxNzIQ7xRlwy3/vX5K8/0C7pt
pYHeQ9n3EUTc5WSdZh7Wv47XiKuf/a215MAOCzIDUrZ6b3s2p3LA8wb5ihyRCZnLcFFPBC3jldLx
6dDFiB6LC+jc41W4yIjQC/w2NY4cRK8mZ1uoIFlqiPgFH3kWNCp79x4ugNryW9XcZ7GFp2MeSoUk
XsFLGNwDkkKHiyjWxCj2oG+mJGTjXUeIzD7z87nY3VA7r+SwOj0EjbQDjhwJIktslF5j7dPJEJ/r
i2TlixuQK2IeajpEfmvrS1w6UewKJHW1YIz+kUqqwqQFycr8Ff7q+xZgbEKcpANO04khKWFQ0ZgW
zkcC/pzn/msY987U5UnmyIMGkhHSEfZyAl4w4lj3c4VtMDO31CPvAFVVLUtamroARDA38sHOBq9C
ICroPTRFz8rV+y0fyzGOhXYsgJ8U5EhvboyJ/f/LMFC5XUOOS8OjSC/m9vzVAuhMK1bt2V17TLLa
eOoJk6rXOn2sGO0QvWrG24zpLP+pqG7wpMxLm6u0ivkoSgND+Ou2Nhp5yK81exQwVOqg+hGt2Mwq
tnHLoHQdzHls42xBX7MfsROCZkM7g5A+NsQxe0WKuJb2qJGQpXLi9PPNHyjKqg/N+E3IpZjJRDXM
3yeSMSqvX1pq2QM6Bimwr8QrnnY4ulbSgvfuulFrM7IhmPrvD93dGNXhNEtVcK2XRxiVrFO0vlaB
CXxFN2ERlxKDr6P92W3sESIo/ZNZ7J05Z9YY1FEasNE3qKEzlAeNa6pMDbIDTJTcH0wi+3eOxkTG
/uowI22dh3sgm7MNqidoa9q/O5t7vXXXjaz4HvMTP2431SGqcz8fusEHOnEgnE+knuE0U8AfdCfO
/hiQJls1ZvMWN7EQcbrEntTtBAZhCcD5unpIh2u4aZ8HSrD5qPxtkGACiPH8PzvjQVbhE0FWPxLk
a+vhqqEmxwJC61I2djon4Za/E719bBzgprntqirN7fLixtq//HSCUgoqG7D1qucfPUAaFeeCFuFu
Y9nuqwai9k1hxTx6vUOqav/rp1l4rPAzjNQodg33J8/BvCcucSIYKkC9TZM0UO18f+J3dlUE50K3
oH/k/5YCYKS7j6mr6QVnwFR7CBBFUlbxRDOixxsNIqYX06N6b/oO6neeakkjrnd0LDuP1z2NumaT
2Niy3z64WPvVtkjH12jI88xKVNIQKhdfS1kNkNvovNtSLXAMELoCe9ZSCcJ0quaamrompeI3IZop
xD89EyTGekEHLK9FuCjtaOzL2pMKlZLTobfGXUKWnjUuArnuOO7TTv+E3ZkhzWubfN3m8pqeOJ08
oD0sd/spyhYbOK3C6W8t3kcLTw6AjGq/06ij6cband3h64o5mKXzYJZktanbP2EDNumpnxKrZ/oU
BuV4afVrkRugNpRjzjjv8dDrh03lqT5vC54VydlhvWuUGaosy8kiPTDhfJKr5ZsZ9OO/rTn1OVH0
OlSSFjx5Z4bk5iEbckmsG4YUTWMvy9wEyNAItzMv9vqPcOHIlQiEF+gpG2OmvAS9oqLEdA4tWPvw
u/rx212O/oVU6RIUO1Q9jsi69S7QQVO27NW1Q+ruXXHPyhi7tEClt4SMwAoRcaEJBtnl6U9GGPvP
kyN8TUV3tEUEO2TODpGziyYNycvsV33vCdscWmNqfrtNw5wDFqPdUsw9kiiQLrULqAm6dWuBr/lH
ZVXonBpvd2ft+PE8WjUeo8hK6EU0W1Xf3W6R81W88aVm8YeQDfXhJzsXh7LETPengKqX2vTvMAeU
MWltCL9X6skq+h7Pmer7zX3BqIo7+xI5o2UY+nNwkdzgonSbhRJYosR7Z3PdzUskIdBxQrrIk2Ia
A2sQK1s3xWes0ed3JxdvptYXdfm3JI9NEaGYhbywCT319CT2gyr2kdn7zZPmmlrMtdogIVpsY76j
Kb1turwGfl7bFsHPur6jA4GAMLEx4F2ih/DoEyWJYmK+sxuuh+21KE4qxubFt08xRPFevm8fMix1
fEF42jmf5ux2SZP4DX3fzVcfqTcWeqhsuE1n9EUpIcFMaYX07YtH0f9dfAyHro04PFOZ7e+S9js/
Pft4l+MJAL0Hhvy3A07uzkzQt18G2f+ZXESLqe1Ab9TNRhQJ4HMvuNDu4m7bufOyKfil4KW81E6Y
ZjTDlryHf24nA3hySMtCNONzcU2CS1CMsgxlgGAyjZbkmqYP5zwsgcax+KURbJe0cgVQcuNgoIl5
EnpMm/CJt+cGTCR3DqHvYewf0WoF8R22CnPbHouDqlYBpL6NHHct4cHRQG1aq1x9yPi2rJ8CWDLa
Cl7t6J1c0KUhvW1ZUy+4Y2ZZoq73MhwprRaF06j6zfuBRLJ2z4EhGyfKFBpLHy+RYsi+b8AuhuKu
844L6d7N9aziTSTqIHsUWNDiaOkMOX0KGR9+N4Enfo32P0atkyPfUNR4YsMdxmeociQXu4afiwrR
cc0HRAMlmgJaDuyauIfknDjmdnk+aSK8bByVaDKmFeOLNmCNbLFct47rfbGsrUbUZlDkQCGAVhjj
YI0RCADygIppvgILnpqFwVNB4mtUv7j/S5rdSX0thS7wbBEcGsWkHtyR7yTi4DoMICz06B0ZPmsK
P5MAoWavtUW6MkS/4e62oj4Q4If6PAOMz+JT2vHSx9vVt/x5JOaNUIa5dDH8X2FVbLujeDuOmPiR
dLxPLfjuOr+zJJKK2upPQYiks1lJ9qVk5tQlzo6xqXj4M1dySF6kjTDuOsRi2hgU+8oIV26D/mOe
wc6BXd6sijKQ2VGKJY47F7tCmeHY/P7EwTx9ltQRpor8+2vC8BVoPFY3zXI//jidPoQKzc+X0rex
rSEDh1y0NxNnpFVFLMMMZ8pi9dhQf0+hr3WEOzKPvJWsHe7xcPPhpzJiuINl4m0nqV6jenSpgtL6
FP/46F/NzKrI+fUtxcWObd25E00CM2N9Hxm1f4BRChIxHiHVpdMPXMMekq2hd4OzuwGXZQwE+dXY
li9i85IfufiiCBpGAHVcjjX4RzXAAjVfNYWltijHEW5IuBa0noa+/f976DmxV3VOJuZjB4DYdx9y
Nwe3ZFivF/9Huc/nnCZxWsQiTzNqP3UKDwWwdy+yAcVmpDGl/IUM6SnXoZwHGZ/DEnO/G5L9IFg9
bdj9/dL3pE5eunkYC/yxgf3Xu7j94Cpqst35dZYGIMHfz2vnIX90EIS2w3UuLSC1PCUonysZHCP8
NeI434zvRx2L9dNILOK4E6YySEfuM0OSXUImbzusCCBwiNlqz73bWPIBwHslS7N81+qDmTtK6D4s
IDC5v+dKY4QAdWOSl3bCVYYg0M1DOmtvCSEtcNVqCUQm4FCYNf8Zpoj5WpRfi7abj/lWF93qZbvN
GcmN/KullNyOT0S8iFTPF2g9tTDbJ+fyWCkVRLDUi4B98iY1yo0xJPMhO4QvUFUgJ9+CALHw6ZHT
33+e1as0iN0U5bZ4855OK6iqujPEWkUqyJASsFwvqXVN5v9l4+AqSDp9Dy/uOpZ/oHT/Ls+zNYhH
/qigWSAzyy/4qu5FVoh6njaVy3tTGeUjCaHGDjbSOxTJE2qIuM2xRyZ17hfPhdw9pBmwRgldHz2Q
Ax7BdJ0BZ/NjzaTP0ICe+qKfbo3MTOzzrT6CyB21TQYzcevaFRKtodbjh5xufNW5a8fjh7bB75ka
gN/O2dLgqE1cEtWa9tfDJm8TnlmzHeLYYOGtTaNW/gLZZsODaLVdeFhQvN55pRmdbEXSR46eofhw
51cvOPPP6RuvE87ZxCLPMZW5g3T4BsYk5vsnzZoSeqnOenUnxIBfW18/tYGCWwoWqFYcjP+bTW0H
jFWO42HSPRo1mwlHFk41rgx+qxD0er8sY6DRUvG/wo2w55S3TIkaLU9uKJQPHiGXgDF0B+6jokIj
7Wnu4ZJEywOloGmlqhBfUXU+Hxn+FtKhiuLmEKweettJnCQrM7ZzUJDQuc6Sea/7Tu/AE+SO+4av
KevRf9PXh8rzP9sVOtMHTxFh0XdMGjdqH4/oK8i+A0RGW3RhGIgTuWzeM0Eie4B7MDXEM+JFxgrD
ycFxJzlXyV54IY0vZDkBQ/jsJ/hPdDpyLx/w8T5FE7vzR2BMC8bz8VdAu477zEklxr1PuOWsBuY0
y0CydV7Bc0OVpdIOBunXCSbZa4+bqnnQ/Wtr4tBsUNYr4sHjzPTu37nP9gFlyjMrVZg0PZXYDDNw
YDE7LLR6H9biJZxHVv/fF1w6yGADST1ZOnQC0HG+7ZiEfRkK1f6vHOlTc6HS2LkFitxjxFGj+JrY
GKZ7Sg9ma5i1NokInN+tt9mhAnhAByjpFaF89aNgr0ueUxgVKhyy34nAUUVvckKjjPLu1dv+Dcl9
g1B8KMsFuTOonV9eu6exeK1F5yFy2ZtYqRB2e3ONrkZ5TU6RI/cBiMKEKSv6Wl69LTDL3sk+t2/T
HXfBmxedxnWAo0mQcm01cEKkGwNUWdf/dI3tu+sC1Ry0wxUmkAyUhoefIup8mq/GkpFzhcLZLmSP
CydqbdCYiRS0dHCNOrYjY1ITC5Wxcmb4WpxpYrvVsnZAEHCO7V8n/QBJrpL5G0Y3o1vlEoeD9nc3
mA9H2k6gvu9K7eOdBMN33Bscv6x2+mr52l0FGQ85vPH9UB4Mgyellk9+e1EHUuOcJ9uVHCYiraGQ
XQUGA1FS0mR7Ma8PbnjNaF+zi1CN+2L72PyBM/bGFseFV5kIu1R++pMoxUSXEt1aimakXD5QBY7o
+aZTPyfHARHfs6XisJlqgz6uYM718aAreX7udTwAbB9igHMRGxi/1kYdtzDpYuS8sIw5R9SnHWw1
UFBI0GmkIWsCtNMiBW6ShGBNNZVm79cXXZ1IKhf7CXo1e9zAZ5riRPOZ4TLfTZt31K424GrqnVMm
Yjyt3wifpAo6Gij7h6AjuxEbVbd/BIJYzl6nptXs5xBVvf68kymQEg+8wpu69LPLNYktdPvk+KW9
IcxDIZMkJgY1k2PknqnYtNe9YyU/RnY6wp/PeIOHJDhbHWOe89lLxZppuDciAa7nJRl2siMI9Fuc
nAFysPVK802nww+RpEsoLwCNyvRGv3/0m0G9B/yzwMuf1aX9RJTaBi7AZlPsAzbBno6/OJMNzQzR
UIfhKhEz0pmZEzg0HDaYo/fzFB5Zl2Mch7LEtZ7cBY6LUabIULBro+PiB8uhFhwbu0eS9oDq3VvT
3BNKjWWc0Lv6P9entLwq/HnkK73yLtMNGUVjHA3Lia8A1yaNT6W+XwFiptALILYobf6h9wwy/xhQ
eFgwrXhIcLDzRXUYkpJCj5oD9MW/olNPn3poL8kdskrEzeRVlD/Y4VN89wvi6D0iRb/DSwqsOYHK
umjCoY6YimdU4I3HXYQS0caKHoQHypX/dM9NeDBortzU717fVnBHgMN4BmIBZZrr33/iWpQD95h9
GmIGo+qLufuiUyfvEAoORx81WFTAuqxCYhHeYsYTw+MdbhK1pmZDi7+qE5tXVClWgyUq5ZBWeGQL
XlR+XhyGsJKwfEJlpiGCJXln3J4Lv9MDYbkh+z2HzuFFzKMhNq+qugeQKb97rninA9l6LtTwQBrv
ysf/c2rUDc7fL5Ik56RYfzSpnQU6A9os35Bz4qhQHpiawRyXELKfG2jmy9ZCe3EAEt5iPsaKchRd
Tsq1wdxgCm8QnzpQxa+mLYfS2K9f6/6F7N314Zf4nI6VoG73f5o67FGh+RhCAUUMiX6B6Y722SG4
dJadGNJm8mbFglGn68FY0cwO55DDvGnta2q23Wj9mELvg5Q60s3LvaPN+W4NH4uCzpyKVFj2ols9
cxfIEeZw6/xts3ywulQBa5IzqVW6Nr8l2hfbnPjbLzVTGbgHp3sTVTFv7oiQk10p4xyOjbqtisUQ
HaBLxdC17PA3GzG5dOuPiJE3Nldu1K81U0IHtTy0mglhd5V0TfxsFCdgMkuhJrXWgo0J5pZcJ0Ym
+scYfEjqhw1p9rnlgkS/VgxFkzgqpqXDtyheN90KXAvsAiXXt5YmBpKBLVKR/LhHBY6qd/qohXNl
Sk+6vAmD3uObRaCeNb7Kp80ttPuTsb5UXJbqlL4My7kNeX4P25+clF/2OSznjtETLMBNbFKq7HbG
kdV4RtTb1/Y/AMjv8uInSSwtIHimGgGHfxXThOfapwIc7obcpjjqhxgOIhTA2i8LMrCWHnGIEtjP
M8UtKUq1Q8H5WpiO75GIbc0TSlMzCN9d+5o65IhyXyazBeFpebVgrm5zqhjEN/NbVeECfJKtg5vO
W9zmbkYebiygIxkNlrilG2JsWvit7pxJpdCoLuaR1iExfVKiMPrZtAUq7ghx+Qmaseto1F+jWEVS
JGXUFd+ie8oYqkEQOFfFtn4FPj713nKLcMIOQ7x7+BPKnjEmMdImcmJMNa7Vft+Rg6wJOAm3DyP0
c2u9QcvFYJ7z0eIneaR8UmxQynFUsPBvpRT76DRtp/W/iu5Wma8PNP66zwxqYXMNvXUhc82SqQQv
ReypwOeKNjwrd30EaC6qyUrp9xBiIoxqEJk+6TSF+O+Ev505fyLRDTdWUsuSxuxwft3PJtD9qXR5
34psWvxCciNGDpTZvVDvQI+gEuFYz4yDPndBRLLAOUhKdq4XQBQiBxmYPefd6dwTssjsXuNgJcFl
ZAbQjPDLsbg1KoZnSCO7F+P5Lfkp7oO+ubMxAmaKYvp+DK1x0S8Y7Uuuk/thV5wvYFYOMfQtDHIX
9LreiJp1RSeq0mbmjrR8llcFxpvvrGy4Sw+W2uC91Fn1fpUed1XC4AQ9dSGzXeAGl2gGj0nCQ8Mu
0AukGIURLnspXenJW28LySemOQ265ZRZB4wNulsfvtJqFOUM39RzguIwzu4lWIHXP2SEnB7INux0
WgPDpMuzqgnywxC/1+rYo7bu4QXUu1WUgJXTeGPRC3gSnxAv+/LPgKAcLQKNEFbKHDLO7Vi4Wltp
raMSvmsnI9Ep4Q0qcPJZ8djidNpIcjF46f/OQtc9eJsTPcn3zseonmolyAj5j4whVP5QvwPtjQ3k
c/qEy1qm5H5W8dNEbvI2I+jjZ2kLPM8kqRx+snNngCpHh35EhkHWgnHDsZ71KijI7W76DZUqTWid
cHwWULrfGn9/3UU824zl7fDs+ssOqNSfVJTZcO0TNyRDTq4HBtnhokG6W1WGtBupuxMwD2EvirI7
TE/9kKYP8RYxIMYffBrQgyd7wE5IBFWmbBvaXEgRXeO7rvMfnFwjf55sLIjHFbwctZVK5L0j+bzM
x+rXKdIxkJPXZ2ndsqeoDXF2r0sqkZpRh5yFRlHWffsaVlVUzq92dfhIauoWQUk+pzYX0olS98gZ
SFhIzOe12tLO70GrXoG67ljZiPULReDl8tuBCeZFTWCqeug4cFzngQNdry2i6nRDfWKf8GDj+qxd
aHPba7wAMaJSHw9R/kAZwp51qcuJnLACxA21ds186VjwxU4OwXEFKoLZKO/Bx1JZHaHEW2kDM/1Y
WCouuEVS7WdC3Dup6Fhge0g8MwW9eKuN6bY07nn5Dl3Zu5F7eQj7t8+rUrYBV/cuM4KqvGU2ojBy
TYkOttZHHmIp1rkRnHtiEBqiGJ2/AOKLbjTKy05caAKBeTe4+gOZ2pjXV3h8jkCDxnDVbzID+ysY
wlQO88mhLHTUJNt4mhintP/PHpPAWCz2DTOAl85OyFy6lGXzP5pCOp+I1erhaEOCtS7gkDlI8vby
3kQxqBWvFcS7J2YGNiUtI87cXc8AY6Q7W5e7/TRyh7jFIHqDsipbgZgR3QWhYhhn18Fy0KZ/1aPQ
lgyivtQesQQlXjhGwruc8fL0ItfBc8Cu858h6ydNY0wKdgwr1ZPCd1yV7MQXIdAZg0RVyqM9aOQK
35N71rrQPjq5Tis3M7b8fC+N1mxcuCJ1sW8ATaKhuri+DWwz38nfhaM9ccgx2mJHSmFfbjjfa5Z3
G1sn6hmvh4nq4OJl/lpGKQLWRmgurbctIk5vXxEnp456zjdnbS4THSlkyRmqshq37zqNOWtA3dxY
Ps8/lKTllS6/rzgRft69G6EW8VYbQoSi2Cv57GXjCuWiYBAzWPr2fnoRBwsHUJQdwsNrfATsG4gX
pZxx0cxURq1wBWWZNPbT8ineeoJMA0klFxxw1L0UQScVZLc15QAOS64OnfKyIburBhGK7us1ya9Y
8kihpyozsiWROrYGfTAfRv2DaK64owRELYn95mUG+QqffqM4oc4XDayvq80bfDvabf/HCuj0/V/j
tcM6pfv5QeM9pl3cwWe8rDQZB9hDvRS8Q/YGD30vSRaFJMCQh52PzvUYZajlgV9tYfwpQTSKngJf
EvGexIXU31jRVmSbZ3VryuU/PZSlG+JMFf5WB5YrJGcdbAdenI970phc3XtAQn/jKSW0oVcjOLkr
Ne3Xruqvlt7+56HSy6zXCljajt7kn99JnugP/EkHISfkma2LSiDIXE6eD5VbzcyiIL5Bd32BvFcZ
iYqXgnJWx/f66pLQOps2mjQVWiY43rIPW2Bvm8Ou43zjN8u8o3NUyF2C6tIvRanZH3jeCVx4g09+
RibcNhpiNh/S2uZtW/BfDbCEUGFo85O68G2S12HeX4UAM3TAXiCgzRx9f2JEGHtlrSWHsg7wz9jp
mUzXKIjrQcogeH7d5jhlTqvsf0i5+vPa+NUC9BM4hqKTbx2gjtgMAxDAqcd9GS1v+oyAK3Uo0R3Q
oId7iy/Wj+CVYYxH0aWfSUN7DOrTyG/RdTPXAkUtQv7a/5NT3b8mYgl2avBwVCpstWQsAQJ5pwZY
lrhxG6EQlO40LyXaKQOw8vLHBqOHowZGsyGWyWvxSazUX2IGl+oFxmXrUrYV6nMLD3c38nNdDje9
OTRXmVlxqHWzP4oNAGlcsSWd+Urn3/5ilyYaHpYvdg9aJp06W9iAzxV1wWXQXyJNlk4lI3io9t+s
hYErNWDEYh2+B4TWQZJPoXTnQ0KttsqZXphEXY4lE85Jh2tj/1P6eDznro4y4xbICnM+zpxIb6aX
EHkPMjuWDj+g9itw2to6E+2SQl9r4dl4RIZdphAC2KOsRyPKeKrjCFyio5uFSz8UAsICCWXyD37W
QYkKbGp1uX9kxVj8zMeLmy77s6YaVI3R71QIwRvCJhhcv7H4Tpos1K6hVVGKYVUdQGMVHu5I7RwC
0iTqj3ByXzpm700J5MlntWkQMKAORT/MCqy1NhccwNC+hP6uyZPJMBp3jnQBP+B5XeMm1GRzqVrx
XxNyjq45B8KDOarQD43jZop8IeCQkRFPo9djBzKC+xpao1FSRIIGkF+NnZq++MqfVrtdrCN1Zzl8
5ttLOPCrymBdUc8BxO21ffDWFs0ryG6SQy7dE0UWBX20X3OXPTFhZ1tb6fg6cQ2tDbGwOabYgUel
qUesEMCzTUTI3N+s6nTiCHC9wpG8poSzEoabvRZXJGYQzWlmtaRgfslwtzBMtoAvnc4LtG3eNV3f
TxLtDXOj5zc/7UnBYtFja3SeuPem62wJ5d0lw5oWCuv93XwP8NP+Py2tNxdQCrnovNVSrONUq+w2
dLsHSBEriQNrEe3R/blV6h35i7iuGxwFmYK2IO2uRPCFzoxa57Mv8QYDwcgfoJfncsUCAYpUgrQ7
Igu7RybLY0Esi2Gc8G02muO+YXT8XxSMsDDLEEoVHIACmwvWJ9rfrZUQ2emG8vaW1L/q1vXS0Qx9
iIdpVPzjypzaxSRrIdwvvKUUapvCtjG84ZpXGXbLcoZZWpkHhjox7xBQmSOugwklzaTlIYb+6jJ6
T2t0QIceT+BHaZwN6zzGLB1DrDLQF65WXk8DALu2RC9oRkf3g0+acLKHD4POoXUq7AzDuAdr0qrm
vZe8C0RUp1P2G9T4OhDr7gBTxaUQah3QNM7wncil52nEQMqH0YiPGETqFB08U5lQIm8ZhR/SglEk
SJ0BrHK+p447z1kCcLQdeunSOhRnZQmM4sYIFkzTtBuM35bZeKva47Uz86foS2qx5vhwQGtagQ6O
EIPyfdGCWzJjkFxsBhLQO5/FIAibtKFSfdg/c5codCcuQTQmjie9izOgffqKcMasubrggjVyMOK2
/4y46OTyiDHdv7GRa0EBagCGsZdvk+8xDQbFrpvQUcw1oWNqrTLehLEDCwSUjU4R0ounxHIRdWQX
i9TsLjpnT7t9v8lCk6zyYPQc6FJqH78a9WjnG7mJmqVngWZVesFPbTlm0U+BlQsUzJfG1KXd3Wtu
GA2YOKRvHqFET9uiHzz46OUtQug3vbqpBXcL5X9Yf01ZjBvoIcjMbDnV/hYNhIT5dIndjsZCh8r3
hC1bdrcDoc4H+GuJ5QVXbjFw0/r+b694j0czPB3muP9JLQFV4nXFuZ/SYgdirMfeLQHJat+AzL5C
0bmEvvdEjCGmjqSmEwKq53rN7hT5h4TzxiJJnDK2/oK7IdTSaw+5vj+23bDhTIzhBKHMcjsqgMNV
ZOqCtfToNUcw4A4zSwsNRlcAerNwt/0d2vDAbHM2gM2A6wu6NtmU5j0x82/f4efBy2lUYoUqpzsK
sBbf6QzPjoLm5ie0T0rt/Shk8hVawylccf0JFWT+UYtYi7FdrpUVICRpzfld497sP0SEQP7fKvLJ
JU4LV8BAjbWGH//+I9A7BPEsgBuNM4ivvCPzoC2twavjnif4LHhQlJHcQKVuaycd+7mLjRu1OUyh
Yo1B5ZDYiji0I6y7+AwyS4LAFDeoO2C29AAqszxLBW4y2QF4NCNt9q/TN4iIcPlQn0rM+eBVx6At
6WmJtYnu3kONcs9+8ulHHeZB73sxz1yS12PxjB13uahXHg+75Qovp7lB01Hu5qoPkYmkqi1tuk2S
LqdqA9vLGt51TonNmhOOIqtAaeaniG/tSyUM5mv4kTHKxualBwgSHvNma4Z0ha8BYO9HFyHGpKA8
5WQ9ng+FTnfMmdGjj4AthRFWGN1WiiTBh4Kn14ptg5LfI+EoPJyoA/AZa0vFJnpA/n4EJ+kkzl+b
2O4tWaxU6QqMv95zkXs8iKEDWC8uT/b5E88a1idkuhgxPmlW1vDIYWaMHgat3nnb4kDq4TgO6R5k
FtJzs7RNQREBE8A+tP9kVLWOwOmvuMOLohzSDtFLsZJV71oGIJ25B2wn/0gO+/8eeJW+TwIs5c/v
3wBDtsDVOSeHMMPEGYvg6HxgBVJiribX7Sa8XaE6DCuyjy73hYOVNhskvaPy7IUYVRvxiuvsh/R3
RGpEhm2D9DKRLOJRGzR/MB7uJzfc16vyif2tV3oNSCgY3AAPTXA93TwLf3AQ6ddcQ+QSVSQVKLnh
2vBskblPQZYfYaIdD8t5TKrcJ40T8W0CzbqGl+HThrH07Uo/irXThf53UuPeJCW6mqsnmT2xhCPl
r4fgpEsuxfd3h87F29umJE3s8N1mbdq8PVNRVSM8su6X89kyVDZOW9XzctLddQIxZWlJMjDpeJhk
GYNOUIc1+6CKpIeLIj/Msr1xD4AgypKmA+n8yyIvIzUJCn6OE1JFKVGfbM6x9BMT4nbufvunlkFm
Qm6gb/WCpSSg7UH/CUtj0JttR65Hcoewui0wR0JYhjqlreTftF/cQFZRaKcTFy47HoxeqxlSyPw2
Zp55t1NTHsDZ2dz+Y76fjCYIFWFH+l9KOieckIHfjEZFGBV9HI1xGSmz3XKrKQqmunKsW3jrYBf0
jBhbU0rGE/TrrmrUuH2FNSSWmZZtQvtL9NW7nYKE3AJdnVBMCsghZTEMOBq9z333Vn3KbrWcUwWO
HMykPGIO7VcHC1/sHseTYXaZMOmS5iZ9gNXF42aUvHpU/qZc9EPUmZaoI4OvJ3DjXudsZ1aoIMkA
IyL5GsMfE4QZrzV/3PODRCAYmyXrm7VtIQ3QVO++gF9dVdIFdOJlpQiWWeRklhYbGXKpYb9D2LL5
+B+3/dcHnryjILb8I7IWk2iIjlYXWcq1HIE2TWD6OTWN2qzhs93I7fi6uLbUAzaogokuh2wbTOjO
/Mpkcst1Zxn+0VB6pIgu4EKlqon0SxaPbzwyifgPiPHLfSjPw2hvYWrk90DgLTEjvJfULajVbqyt
RDIEv4jq5ZkXP66QQlzgHhqTWOv6I5aaZzaUcPm1tSd0FQhRK/sHulD+tr/eZ6ObFNOSSj6mCuwg
SE7tIJeKsA/rqkl2u6ZOsuarwdlYafNziQ1TeErT+lE2lINkniXvyYpNZBzLj2E+9QZbD9f0rYUV
fBIuQsTs1iNERT3fmzVeCsGVSmf0tCJQJsajvF4cVFmvGv4vlV+qboM66xbjRBwq2o0F1DcwWTuZ
O3s/b9gSB4OkXlZ1t9Xrv57hJmLoS2vI1RGKtBODyU5JDBL7y6KXnZQrTT8CU1UDdXHezwDXc1ZL
IBh10eNE/zNM0m3L/WXKSEEM4S3RqJ8wROWUrqfy0OwhJzumIv+DDClIw8YWZtuIkJtL45fM5TSA
6cN703lK+B1lsS1fWn7m3DLXJB+8x3R0fWSb1tTVo0kgkn7yXVkd+i4ZpKLzQyHz9aS1M0VERK2y
3iBWiQgO2dbyZcgdH0tYoygD/TLnUbMynubfNzGh435zu5ktjieBHQB9s7jk40EX2j9cXWn3xQfA
srgR3mxn210nKMcsPm46YaOvdGn9nEZ/mpxXHgc3m1A5Ig5quf23TYakwATO5yY1BcHvcAaF92Li
jWxJYoZsx6pRMnHWMrQcgvLEwnkM53rkjmia0ktDKYcYAK4Wc0JLvVYvRc7i5geEKW1eZHHJCFif
ZnHEbVPStNlyTpr3cyBRpebDlWbAwSnankyRTrWYcxKeYpPz2OtrQ6Z9P0BS4ANDJZQvsgKsO6Wn
ssXUzCKJee0vxkMfc7fhs+QyxnOy8ykX/OvRhJ12FUCXSIOKroXLl272jm4xeFcew0y4rQxrIBVe
tbJMU4bvSeh7xxfx/a+9/dkHlhZV33rTP2dOVBsTk+pa7a8c8kzGiyFQpq1lVI83IwRn9OB4eo8i
BjVXFb0XfxXnQdTNLtGmk2B8n57jAh7eu72RdT3EnmNHlukVTGsPuWW8g2xnoUA/XxHxYXYVraYk
CZ3jmMk9qKZJUFQUOV+4uHiSljrxnBmela+0cklxJmQHSLVCioeWcf87zc8eQBrYFac47pASoa2G
By6M9I4eoJgWtRzO6otrq0mV8Gg+5IjYgKV4NHgek7pY12sqfIs1OSBUU5/u/BMM9VrQdXHDfVzU
9+FnwN/wCfDhVoN9t51iQnqZou3A4vmuyzaI84MCEWqE1vfAYUHJjV0p2GK35qglSGnRLyDqQTwQ
tMmn5PQsWDvK7w+N6P4wpSlJ2w4pNNsg0swdfUBwUzuphEZanuiqk8myfxccd0RohUW1f+T2i2vz
gXBG2jAe1/l+m8D0sX0oQS2hoTjCy7Yy4XO/Rj7fUKMlVDF/W4xWU9cWeURGGcYF1m5TEGh997GD
D/Hez+EA4rZht7nQSzJYWyh7xXC/q0nMyeKZBrUxYOlmx07bJciCxd4UkFV1Z4Wq9gXFU8cyugzQ
dcgfaCVhTkaIl+h6CcXJx+Me8ja9vBLf3eZVQiyjMRVSbjWDZmDMJgoqoZ/LuOdW86y8FvdBSQnC
zWR7Nnn990DDBusUWZBsU6PwMLBCcAJqPbI/3vq6PjW96/VUtL815NmEHKRsiLW+Nwx2LtVEnCLd
Pv5F3WsEO51m3wm/46RKU8veYKVRw0qRsX47CSgNb80XPAxhoJmGA6mdwbMD4RdtHXqPykRMTuvF
/ua0z60QydQI0E3dVwdBSMFMGyoghuVuRNHaUClmK/V6dbkchGv+05hidSyiolJZpqSnh9CVzCqc
/VKruT/Kzo4hSUBwkEPup0FjdoZx13+LsldezUnRIVLZLGZ0Q5KCmUTfedekqFUf+7HN+Gtzh6uc
laysR2DcH/Q1QuR6dtkaqpvWhiFL7b27zy+KTwGjc8cHaInh+iHBH6JTbejCWYTc3pTKMDuC2XD0
4cp79sKK0yb1Ihaoom1V9hc6T+wmqolwxOkMeI8HII677qgjQWhjJMwCCgoPz142Am17JtTdflyp
eaV89YUEHdqyEqTNv/S0n5Tm5fvi2ty/Uhd9zVvEOizZMPcfRYPrPrOe1RFC9i5KpWceUgq9iBx7
sH7dhefVdVn/kxVkhO1Yg50dgigVl68DgXKHx26ci4RufZqJ2bhFgDAIF796//Ahj99oIvVYccU7
iXC4p9F4W/NUbBzAYREC52VBaiXj2yX7LpzNwuh3Cdk3sYpU91tWlKWjJVy99KpDXuJCUjCPvm0c
GM7mKNQY07MTanyPeoJ+Xv7GbmqbcJreh4vGzN0yO/eztO37LhxWBccb7StOsExDYOWIJ9MWaDuj
XUPeWFNRQbCIyjsai8d4oIRG7TTnxmkFccRQfBY/wsxyym9yBOSriUahKNM55naktHqQmCVozLPA
UjgYwjRirkIKYU2ir2TSG3naH6W4QAhJgoJ9p0EGmYuLhcsd+PHIU4Xcr+c13HlMOXVQIdHKmm9j
7GP5lUGVvNtfunD3Q3qf6fI2/ikCuRs++jiPu+bMwQ1KWUCIiG8+SNG+XQM2ZJ+bHv2o4hOl7z6h
7vgvlbcoogDHkG7n+OAjH93troc62kJDxk6QWQa6TrUb5MpRrIpfMufw6eYD3lBXHn/fWloT2DZ1
Mk7yYwL1gWfiUQob9FiVBc9L70tGPOpL9RH98/LIZbVy8eoo4nU0ZpadljpbvvgOX1ujHpfIYBLi
aqDRlbg1auYwJIjdTcJh4Rlv8Ovq99n+eNbi8DSCfDvJx+jUCryD7U48gi2qRpRdao4+kp8m1VvI
vNpPw8+oW7fPUp57lqzfCCmNVeUJRI20M2a5ukPtBwd5lk4ZcziBCJ8gRw9u5Vp8TxFU0ZisyPRc
UARzPRbYZKEg/EYXVWH2gzEbfHT8CmMIkd9+L0Jy4rvzSs0+P1rA154jIlE6rqJK5yx+Yu1cspo1
Lh0s9F5q95ojubRNn45mBzW4qo+PEX7nEcf5rJtPPaBGd6dirbbNOeKwIJ5LtD4M69jwLYiWg1Ed
RSYuCHmFsBabKmp8oHeuBtzTcD1KdL1MC0+m95iQpzbFYz4k7MZZGv0j9Ps4JiwsS/OpQX2Pt7Rm
jfrUt0pde5nH8E3GFlpIXfW69oWiGZF6slHK4tV9U47H1zL06Dg11c0h9ANcGULGoQCk6HJi1UwW
u/hH7r2QpPm3QyR5FY7ybiY5BaX0DonXf6rUK16kJbsyikdEMMQk83cudhy7dgNX+J2jop4yN3Se
md1BsCI6Hth5crWJnDqa3eMOex3GzCc/gv5u4bnkPToV7gIXZ4eJ7QbbcPbjjUmWdAkUrayfcwnI
S/hPu9XV4HWFlHebAoWacjZGddlxSdkcZgukjSJ/D25ARmVpVcK8WFNWndsBHB7SZ0gFilymtuab
Ol/6RRkhP/V/sXwRViuCZtyW6VsrZKK0TJ9SheWsRuOHjfHQoISFAlqUnyQm1lGbS0IVBGS36jvX
iGxfe2q/hz3QetDeNm8+Tadnrzy04gzcCP0LK6UXBbLKlkWG73jnqFVkLFXPGttkWwfrPQrSRgY2
KCIsp/Glcp0Fc6HGlETxrgQsrrScbp2KtUZ3uMWfDaP9rME9ZNQicr+0umOeyQHfpuQ5m3YPQV+T
Jxdc3uVHX77Jo+zIC19U2mAbLRJj1GGG6Q3GADfd81e1NlWo3wcpxL+/rvC4tP6l8C7ltFXixDFi
Wn9svm1LMnUENneL7M9EZt+oE/q+C2PoL5Qsg/hLIQY9wHcUgrzw1dXqS4UYzVSYo/r9fOgkEvLk
zHQ8exa4JoLjUxEfYhYWqX9hwaIn5BXDgLscxmeWWWAw9Tb8agoVhDBM7dEHdXk12xLFw1UO5rVk
5ULH/uoK3Wya+UKtc6Mgr84sshjbGemqVIU24Utn8WQ9j1gOq5ijrCP4zgp8KQftagMOG+hAEMPP
kjdO4XujALgWO9DUC6LWJa69P8nqypxnm7Of+jDHcjEWxWhD5JpPp6e6gvPGm8WkgXQM7yBPCK1v
BHWxG9YbDj6jJXq+G75cBQT8RqCjVGu5vdqVkBgfBOSGmllgjenPB2CilVwvqhb7NAJFTrLeejGi
VCPXLaMFD4+KZINhwbdUSyinidY8JYNKceeiwlGt8BoHpUXlfU8eioe+Yw3mTtujRBg2etukO45f
TmU628eQ9V1YaPyPFxSzZ+AFV1nKcC+WeCp0wArhHqxZ2kgLHjGMV7IFjR3jN9KUgAsWgdTTleX+
/5nynFxyCXLyeqd8EVxBcT3Krx19H2oBIYIhzSvSiqDMo/3nEm3wjMf5ttwXMekOdXi3vkmQzFTz
y/PaQ9EdTUTjh+yX8qcyvGjVcZqVuuhYRcEfRJ7OD9VOW/MTvTy7HlSqoIBIKR2nM0iJn7MdGlPE
eGD5PQeNISU8Fsk3pOtZZ8UrpPnU/N7LpatWX6RxkhOPmKmnyeJYuMqJXGmwu2375toQUluD6613
zEhNa1fY62MG0/w6RD219prssS2IRwxlr6PRbhUXURdfldNvQajRy35NB+8ioZJnj6Yr/HmZ+Rtx
OOq1c6pXv31Cy7NJG9rN4jAQPgcnuiqJgZg2xZ4GYfNzTzSarDO6t+24YqZySf/Jfea5v6CBaUfk
bWPEWNdVeyis+y/zidPpFGHsIM8SOsuncgxKZLx36YFFu+tC741isfHr08o9gfPDYQkVnuJnEJyB
70BXXKblAEI5jgDhsSDMrtKU9M4oq8SP4K72Ev2VwP0CR1GVMaRn2ZvJkAtPB2uoGJGyt5Yt3uSX
bPAAFLTpo0OyFKjL1266fDJ6rZQMhtXJjOUakjs7z7WXVNjTG+8PtMUN9GCXKcRPvKTJN5pv4UWD
ek1JZhFyOy9/l9VqaUPMHXdmKPHM8jUlmhfj/nO+AziZXe3H7bZ0xiR0RJ7Ym/OhGxnF5sr1/2Ke
vFYTXWPj18M7gGPYaidqtYNhKj913tr5glU7/f1OjX632UOJjy9SmtUi8/icDywe1pmylD5UmJVm
s+n18WAqjydVmNT/y/+UDv3+/y/+jvVfyAZwU6OCLDNlx/0AhwypXa02OBalTygwfYyEqnRGf9Wo
f2KMPQZd/WXBYPW+022xIbIxMSyTG0jLIi1Vv2qEbdSspXjTNoQCx0vlgRSOlzJ0UPzEoot4S00O
+77QLsldNxXG+oJR0UDUn7ycxynySauFG1fofcfwuLb9wcZMr/M6PICw0iXLNpREuRykGQLcw5ne
OaClPN6UV2/XRIOprSpssUbEeaS2u1XaHkLqiWzkycXx3OWBQHu9UFeKCUaoPwCN+QBs8QZND22P
nVguA+OcYYg4DvgMhkWe1OPqKIH97qcpCr0KLuB+4ILtvYtAXP91Aav5jmJJ1RrM0gfYTFnf0JWe
fCaXOyiNHureMR9w5e3y8vsWLc1EHPTuf9D58M7SUlXaTO1NnrhBb4yAm3nGB5M+NQZWa1tOSCBS
1jT6NQiCor0VJxAUBxszJso1k/J4mmIMVRuNkAFVFb7o1NVhXoQ4wFu3xp9C/052rafBUP/SN1ay
4MJy9PCZQ0cLbwdHv+rY6O7EpabeD8bf6Cx/bV7LUHfg8cDKcEoeJIIHGRYnfjO4Ws2Cp2wn7oKZ
pPFCGuxJvhR6OA+qO9OtCmzZPUneaG//8ggQrQYMLS5lSIzvW8C/rtYys/vWZmJtEhR4QYJBievL
TjRfYwC3oJMM8kATufSfimgm6Oto02vKGC+V1W39KE2eQcJr0q23GjO6z3Sdqa06/AWaKzMkr+Wp
Qemxx0N4Ewia8MjJPR6R0fHxa5LoSKM2zo3DMa/quCrlZu6c+nNP1ybAujoBdniQKtiULk5+aery
ewnTdOHlNbxDt7iW2cvn/Jc8NvGzDJaKIvdLgcmbRmEVRarYFqRQXKBYHbHO0mW0bwNs69eahIII
sU2ubteWhys7XQhrRb87id1FO0j6WeONbxAJNhJK7ihFrQUSHonE5o0jqwXQOC99t+vy3Qe0acgG
dfv+JMyPlOUXBFrD5jdhjQpRgTQaOxs6MiUjSYfTUI82ZklAItkz2mwgm9SaKAXpzjG0ztpay+EZ
9Vv9emzl65Sd4nKd8wY3iVDLjzp1OLouzdDnlDnqxAtYma5FnQyJyNcm8S8ZijBTUxBMNJgPhUSY
iujF/E01jbbptV8zrJfJEMfw5PNVkm53kuoj0U7lGuuHMeOEWoGL7bwcxizObbUh9CokORQDbp+V
2ySjMgfOHOALPWfnA+bbh+Pwpx0iCB/FrczJ4+KQnh3mSwbro7K3gnJXlNnR0oq/du8LXsp5p6Rl
JaXm12IwevwdFoUS/kTXLCERo6yz652kOzP9VcFhss5kLdPwxBZZuwe0lbwQb+EPvEgxmKredM1K
qX09pcwMDcHba4jkEhrEGDGAqKYBkElRaEogeYb4jh9SsLqlwP35MIlxkNrqaVLFLNIt1RgozsW8
+UzzjEy1c6Y59bGeZ6K8qCiXuLgzlVI8jrytS3pR+mDqehBgW41d4ig2XlYtmdwP5KLMlRQAs5HC
e45aC9s2iaEYoycvM4hPS56BHCkrWARuMgNdNSAgK3KI4vejLitvgIknwksuJy6mihtwTqmLAgnJ
5l0metyLFsj+3wflm5kuKBMyiGz2DVoJtjfujuCB0QGYSu7xy1yPCiTwEAfuIuCJ1Ga33TgFbWvh
5JmIBbMwrfDN/aArp2uT6NxAXUiejNffAE9NQPwScwddmazbF2Tm1CWAeG2sB9Z47F/kX0oAj2hl
2l4GReC0ZXjpeSm3rafrxm9+R+ZxkI+YUmb80KP4WJE1f1oZTvbuwWusgguKmJjZNIVL8rkDB8Pu
a9xFOxrAnmI6L3lfZaXeoM+pB+O3R743atW7HUxsjPTAqH3bvs/xx1dPKTdnNWAL65+wKG097VF0
DcBlhSIvoijgreQMKmFSxpNRSte4C3zwgtRV0Q7ipvT1wsJgje4v8EUf1nFrKn0Ah7f77fJ/jNQf
xLaVyqT5kk38wGKHZXboJ4xq9rt/mZLUB64Jcg634jSS9KiNmWEsk3YRQjwXMwEcsGe4306K81xw
8e+2y3IKSXWB9yrT8rYbsniFCrW2SH2HvKSoVFYSY3JegzT9x4txypieE8ysgxhFr2u6UVdT1i9I
adOopOjuayOoqXi2QL0n3FpoL3mmvCLKHQrGLD71liuFg6raHEoz7fI5S1H6xusopU53dmz5VgKq
ocuKiPFOYnA6TYEINfi0IEFGnrtXP1DDps8zRcG2CF2mipdT+WBC+u4e52R9mzBkuscUBika8tCw
VaLOsnxgEvuJGcn0SHa4A1aSh392ODlE7COAIRn0xHCqFlJA8ByuaT3NBYGx8AAclVKwLTc3mt5I
ajYPlhsR5wEilc3G+AK/B1bxFGKXph501dLL5MlZMHi569m7cMnLuYIq4Rs09GK9IW/gTU6H1KbG
LyXJrhyvO1vZwXBf7IeEWm+BYiKeJ0Eu4q8lwBJJfts+gYhycNhlErG/OKELARPqcEzCC9U/7kLe
tz1LpzGHmOzoUldz8BWFJ4mZhdc7BCy6tcaT4XjSGh4RL34AMQmIFAw71+z3p4tBo5C9kO6yHxPl
hhlWXhEwH4s9bba/jtofwtp9y7QmrVTBGSzSg4LCZfM5m7bUOR+JgMgchNiGjnXmHwaZ33RI80TK
VK2OZQvH+EiGB8SeSV04sRxRzoyoRjEbTeiZYet30dMIkzCMGnufa5rfYVa7fvf0bi7g41ejR77w
yr1/wjrZ3Ybwufptw1cT9EvSUCR7qp1j4bet6c5vfRSNexEvePyxGGEIKrVYAMPrPtaRAWJ6na8W
ZEQ/K43lLPeMxOYGqjqv0Gx8nk8b1RhTcpHnrPzr+oai7qH/43nRN3HIHrwMLsb5Kde6612Tq9x3
QVNUnFNDOR5Y4O4hwUX6g2QlfY5wseQRrCDimMB4YieTyZfOPaWwzSkkLmarF5eEQShTh85G3VmR
pmu67vWn6nNd22aZ+sSFcWUp5epmt9aDw+OmRsZnHiMDrqbTwTo8MaI9Q62FWbo+D6UBsZ+0GZC0
gMinmPG0ueSg2qb5v5KKCiZQOlyaRI5x2+FU8IirrTinwSY8ztwC1W4JersTnpXp1+RzsmuauDXd
HUf2+rNKXIs5ppEZEqlFDWctBvKCTa8AMJuXXqK3ZGYTj4Zk589sI7wrGAGb+OBHISEbR6SVIDgd
byOVvQSN9XHR2b8afoxXg2mQfcNwI/4U6ANiLuE9XBGZ6SIw4wYIziyo06Ab+CRuOJA3FogicWni
63AiJqq/y0f+I1LzuHkYdAjo4hexoTE3H3jrLq201KxfOTXD6qeEL/SenYuojAM21VPzaWNKuMOy
wItTzO3tZb6/GZo+Jgy+6GTm33SDrTDpsJuMXGI2ZT9K5E8kaBI33XK930NuT2QTX/cEF+If4DLB
OaQ4L2T6gtueTlvNSErUuJ8YZGc8I9au10KR9m4mcwrpzRKTR4pFFW+1rxz8RwfNjKSQerMDFTPc
ls84DF0Fu6n4Rq+BFthLljIQG/RpPrFz2IbBYfo3paOblKqW3E39lh0lsZjhwXGS/DVfE5iSN3r9
FZKSUjVbV/F8FuaPEu46/uv4QEDAvuN7Zdbor13/Tc30zfZJY6nGl9Rluv7RSMOkLn6ia6JEMqEf
Cjv8bDkDH0I/ReQes5+nVsSJ1SrXJ7RaQFgpSx1dlUBqfi8aY3cTD032rCaIVPfaJxpsiVFn3DMY
RD9g6b0SLXWfZvxVOI167KjSzxUY3OcYJM4BMXGIsaCJhocw4O2DhZ7bPTQYTzAEXlJzjmelu3/P
M7tiH6bomWXE4OU4SzTyPgRXJSKh0oTmJgJHJnTmWtcX74dg6IgcIdW5PHUfL7bvs3dp0tco5QuG
8IHNkWvaBF5GiQLsT+WnyZaWNRuc0FXsSuLOIkdskyhLNdz0rRW1DoRzx6NhW66BWQU+jeSdnRxq
W2Ki/VmnbH6kbGHdf83jxFbPDSru2bJSuXGqvPKtE1bCj4qLY0dSJmAP9XKZ1sAquJoCqJwHtqbj
3KAW0Pifjba+gidinAEpAYcGNCF50yXSCCg3GrvMN5X2UrKebERZyXD8z04+GehnU8MmcBBAaCTx
LmRi3LIL7k6lRQNqFDOre201G0YAQBFDSFpcXmBZAhIxIYj1GKZNR45TK+42uaEQjJJv3Qa1e6qU
GHPDSek5ALaMC7Iln8oQ+iDg+9MvE1dSF8kvE2NmNlTWrwX6tO/NWkXsYqvyKcViG60oni0SMyFM
vHRNXv2pnbJp6fXXa3tgTAA15hvkMaxuMKEW9k3GYOvkMX9VZk2aCPkCTc02kmIt8O8tBMXWpnIo
2uYAG80VJRUx5dcgK43Wn8XdnmMUaOrW6cU1UhmvQylSgAip5vnkgLAvLJiaM14+ok3pdZazl8TB
CMBZm6K0O4t1sIRXoSN5BozcwD9MbOVnpbTTX20Ri4J1JVpG6aEvSZRNqjtZMTW/2l69rRWF7Np1
2fJ+4uqByidkebf0FbAThOVp50ZGNtxyHhVbxEJzkJgM1pa3N3VuxMtXGa/1EyVeSrEfFVa0Fwkz
plEdHRyaDye4cHnHBJMmw20lhX1P2v/2UOv+i0p2CVJVMuoCp29hqWOjvI7sGBYoqFKZCTg2myTy
ZKUJQ7cQ7LT/27NOpFK2ebWVkKPT+Zm/F6qMjtzEa31k1zk+cfWRQxSY5qZqZbmMBncmcMysRvab
reCWcOC9cEQiTreLj4A8qpJjh//VGFsjLSY3oDUDHLhEmY3bjrrWvRrtUP/g+BxF+ONkQuyS2h4a
EoEj7WdUuq5Is9dnF/ZKt5ksgJQnSMz551deenvdRN29/JShfdCHFzESIiGQhklvjnm1qWfBu159
Ypi7DgC/BeafUSoJj+5sumFCdLqgjh8pbwRctLyh9tUH370JgeJTy5GBJkc4Bol5APu1Kyg06+EU
DdI5uox1EAsjcWxrJAba4SMyKbcf7N3jHcEzZJ0z0sM0vZ9OI82ZUkzTskkmP71wJ1CAMEMugeVM
sZyH/QPfeW7PJaIQyW2nWgtj/h5FPQfQaWOOIp6imLcZKQbQNvKINL46Oc0ffSBRnuER2UiJsHgo
4VHhZhbxkh2NXI4TXJDRixbvf4adJJSZJylKMbNQxl6wpLQObOqlefqN7A5Qu7a8+xPZA9EsxpKd
NTYEb6STHNfy0o69Dl4e0Sx/u93NxLYbYr8TV0upAEfoebcO9JDREaSNVueDdCucsTRcAauGyxUu
5BJSTTpPx8gwjzIk48WYQbUlLTIHacKtmXKrUm5tQXgNhHGHe5+G+fqchhc680w/aUluSXwqK5ri
md49zo+6x2eDemZoNubR2EbkNB2Mb6qkjXglrUz8dbdo4V1fpDZZ0+7WRxrsDhh98ct+zAyXTTNI
ht606Hqv1yIISEcE87g1lYIWkaXHAom86cfTi+NgABdMnE4puqIFvEFKzIcxKmJVOE2/V3sQPm1F
+k88YgUzlJ0b09+ZZXpIdswjnGE4DqnDXoQCbAz1GSXcb60ec/MKyGqf5e6iPGJjTVqUHpdFA3+m
Xp6qQqsuyOa46m5+Vrg8VnAtIw04vWGm0FjC10Um6eCo9bQwIK4JgwDB6Rw4uOuvlKEa44izYfLW
8cRZQAzXsxZHpMYDMaAPI39fWGM0z177Vmih9pWaxk9WH5tWtLT8+Prbms+I9+hNm82m8t4oVtVd
ABNmrceZ3meKCIH6lxfBdRK5SW+OCdrPZ0XaxDOTGS8A2VQ2Fe/hq+FrwcaipfNoWGb5ZGkFmCEt
RzRdV3n+NmCREBU8IsUuD9P7xVV11QZ4saJwErH4BoDhnYWNiooEB/4eAIQQd4XfBA9AjnHLv+Gw
2HkgGQueSNP7MhElx3RwvzrQOdFdOZgmXdn6Nkyvbi3fDl2UHVWYO36gu7r/M4ptD60yyTregg02
rMQdfd9i/05KhNVqcgmewW5K1YRA8iujd7bVKYqALONNGZ3RcUCFa9Xdxu+VkF1t83wHWcHmL+z9
Q2y04ltdEWZEpq31x07OSUzaG6Jdf/9OVXudDhtwyDMOxqxTy6mjr+UsjiHVwBAKssuYc/ghM6WX
qY5JYl1IuYHYKOqgmfPo/uGpotIVZ5FMiAgnaC0n1jbbkHCIeNhaLEM5oQBtQLbLpI1xrR3E6NLd
I6ZEYroaMRUXa5wOFkoEzCgVMx8nnWo9nG5yI/mPCXDjIRGlKYP+CNYA19M6MxG1bZAk9wXaOF2W
Phvl9udp0RLZmeS55INP3qUaBCcEQJB1JrXZCtKt56YCkCeQiFNugzNsW/vQLjbeD9UMmWFRwUIS
Pu3hTt68fCWUf4+nreSvCo7QTcVdA7ImV+I7sFwZDB/hrw18rDRXXPYwPLuheDoFsFfp41Skh0nK
0VZz+ikcZUaKlo7SQuMhQIEaC2reAdnZIAZYgVyAfM6PkgV+2iNvrQD4ybTAu8CsPdSE3FhAVgoW
LOcjFZG5xu8fyNlU2bYNyrgzRHXcnFGQ3TDe8YX1vcE6Nafhh/DkVGETjCNISTOY9CbAjFRZsdZK
JoI59con/0n8Qx2a9NI4wyMPQ6M+iuCBNgyvuRN+bQ2E8ld+fhilS7x0SBMyYWqujeYzMAbjGlxW
5Yya3MwAJNp38TsdaHNzrjeAm9EzqPio94ug5dIF83QSID6rOLAvTtXYgmt3se6S7FyBxXXixurt
7AoHewEUGfkgwAW9Yuj6BhBCT6oEVRkjPiuWKQ2XljLJ7JygImc47p9YfC3SvaMr4iEUGOPdLH7y
8UMPEN8dsRdQR8Ey6m46cjl7LUH4or6h3j6zaK6O+GfbmLynm4zCJa3h7u3h/PPREQHv9aXDD7C5
kl11pT5Gm8QfEwU0tog3AhEAKOqykN8FG5GCecDucPE09cvwc0yVWZ5/opBf7kIoHKPBl0/Xfvj0
LacKyMxrSclb7JW4oNh/vR+HjCV4+Yiz6YcJ0qAqF2EMQ3gqCuaBywcydjxlCX4HoczmfOfXlKF3
MBK0JeK1wIOtRkpzOVQ9aELwir+H6px2i8NEZSODAs0VCB1h1IWzV7wJ2qcfq3EKVxtdcPKL9ZtM
yQZgeUYSx3G8DJ8gFs6eA7XZGwt0gezenPUh4Bd/dfJz32ixJNGw2MVci9q1S0wjtLvGlG68CzRl
w02gweStVdcHe3QsnQYN6NJJzq1j+cUr0z+XgeBzPOAB2tXq6u+0iWJDexHli8uNSwBqByRGFVPp
ch4lEtqJlIE40Nv18UZ11H25hFJGgFhFkV6D5IVROM5bvs9u8T8YXtBx/wQNXaZKCvgCE72agj9i
Ow9sES05OfbZWe0XyGGLIgEQ9dxycakpOi9y7EfpCyDBffsYJOTAXcQmpBeqQ0rRynl8uvL5zUu7
q5D/HNS3OfOL1Gaw6pPD7Y1LwD00/qwgxHOgXIZjkHxGNJq4IROJ5ILeRdGIkDq113ZGnia5T+H9
GriY++U/dZgQ+7S+Bq1GL4MlrzhGlPOuowAayExbp5WFRFcNrVLSP2+C+5LctldL8R0Ov3IUxRhI
RlaTjlZhrHeRrJXHxM9Hv34m5uDrtspPZdQt9AbhcDPD1dhPBnKbN/JkLbAIPjBfsbBpQmYDoV2d
VhHCb/mqtTwNbNSTT2lPv4Mrw+Try9K0+kqZSohii+C8CBLtvUfzjEVr1jItwt32RbEcZ/gE4f8D
bP1e8NwLl4OD8fwi+YZbGyRZ97Q/5g95CpHTc4L3Ea2NtFSvs5Z3I14OUEU6HA9vJ3S9GzsjUM28
03Pbpz9FvlGot+dyrXc1zkgHy8YNmC9+q1XvMnAOBudorAHfJZPS8fuhNYS6fwM/on2x3Oc31UMv
L3YSQmHBnuFyWFfuaTvxAFihh7v0DLU75RvEY0S9n81uQXbMEu7n5BPAn4WI2evJ/bOa1X8D89hN
eJJF7GcTp2yBrqmrNl0s3TIwVf+TOQ/K2XsTCisX48osM43bHObgwqOJqJvBquNlGn8R0DPUDWeJ
gYMABbk0Ojjr5dazEzZlIU/aR4gG1fN7Pj8zLoW7PCeud63AZejaxsJjq1fI3PAT5WOY4nNKHAm4
dynXQiznuf2jng5DUy9wOqDciC2ZUu1juPvFFzd6J3LX0Fhjse0gBZ+liZ+yU04AfdvzOVV+KPkQ
FjCiE88j8539LNKLERDdI3tAuEn1t51utqvYVx7P24ld502d8Uig5B7OVX549d/1YVzqooWTuabd
waMS0UsDuks6NszkY/kzGWHDYC7miVOuQog83Dv+5ZRkTRPysyWzJ0cCdF8iEdrFmLL1IcXB/ZpW
Z0LNii7jWmIYorkQ/e6bs2241/fxdKDedmLhlAqOzz8v0WTTil4apEwdlSYgVwWtHqAzNPOsYjll
hi4svT6x/HffAYuj12lXaeao8mVqppJdrejU1zZ4fqIcwpFZnjntEuUy2f/JB5U/7YOeKZsBCrwG
g+6xFPHz6BFGamY6d8MTPvWEPWoHCV7hJg4niWKBq618rtpBLGjkbtm4F/U3r4FXGQVuawIPM6UV
J57UHd66GGCy/9HH0sV2UC2LQ4yr2OIbw7n4f1UX38gG7IU/bhsejwVuo0Kb34HP+HRPy5yNTdDR
CAh8Pt4XaU0Idl17ZJ6BeusmCfykgx/o3GlPu4nih0qGbMEqSqqzFk25rtpXEVzwZRvpkbrVM8HP
T32F/ZK3Yv0w/dtZIpKqD09/4GS2awxLufXWG0gkbP+i/dVSdYDeaGJPMk/rJh+W/xKa40PO6PxW
bCuIgomR3SVM/P4BRA59O0oaEDyzohBeJf5o4pwxSZHw0we3duE1P0uLvC6k4vQH6eSVSnhFhMmW
aWx/37ZdBMxWxhsiHX6olAcrr2M3DzWzhg8UC149tPCHW/Yx7Aywa/c5nu7ZGPEyBWgivlJkr+En
NYGA7Vq3RllcdzsaFaIheIZgpS5b+dnY251pf+Q7VPNgtdcPA/fOX8v59Zd7OIi+nIwKXd2Hu+ed
Oh1zTa6N01atX23c8ZIuyzYy4PztlCU4unFlmyM21DLnXFLzXY7h1R6zWEZLNJr6DFUMNZHqTkDC
e3kTbuMtYUNTpzYjQgbCOv6CgvTjasscUb/vvHCPUHE5cY7HZNICd0LOf6YlbVKdnd8MvlzIL0K0
R/dm+VPA1BWnCgG5PC7kirohH1mvoftFS7zfunOubj8GI2J3DHWg+habhwRJOUWd7WvOsBJfIl1e
vxpVDxUYlE/sxA5nJg8AvSNaFMifXWU0h32HowoKb/6eLDn5Q2ChdkUF4PTARbPKBgu/ogaAsP2z
PTAMNG05hcBxeK19ZZtvgC5XNcqvPchrQtAFa3//MsikB5va9tq7klCMSQPgDCRp8IS+anknAZ2T
TijyZQYGJ0vdkMjEflSSV0lVZZ8bnFZD2LK4eYUXtFWnMrUt97UT7W9bbFItKGgldI9VVgITnWWu
iq8x5nmNMOi2/VmJor9CmjezLVbnFPbO2r/CUZYOhma7FM0J7UqRZBHieQip42i3bQqI9b1haPU8
76rh/7JsTgUFZ5SR/KU7gotJ2BveRLfqRsUTQBKkN6XntiNVrZ6GoM/rZlFxrcSH1NnpZfv3Z0rI
MabxVJK6h9rkd8sq8OxmAQVMWVjiC5J9+XNI903jrIl7TvPfVH+9/SdQbX6veKOS0S4AKIunPx9A
b1A1evEtDSPC/NdmN7YFvKzLbNI/jvqJTO1Qonrf1bdkIPXwXXNFmTOAkyniEsmpEVieTHIRTZRB
JEKsBRWsP5U6PhquFsE5CmeC/0rlYj1od9uizb/IH0kl51ln+1c0ntOrJimWvaZKaWGA29gffnbJ
ypjN/dZQ+unkdvqGCSPaGMboi2hW2nsZLK7uIir2NSj+VYRx3lK4ucg3Di+N3kQn+fY44eTGh4vJ
F46DHZ4Iap/R9kpKubbef2+mz8feh9kJ1Pxj0q7YhdR75bgCmcWyl3dFnyFSzB8RF+CA3XnMLRPm
OhK7tHWfLycYbdAXT1NM9AL3kv5FSYHPaJFl60pw2H7Hq7KDzfxUD16uet4RR8SRfsRukbhpz0QA
MYgzVyReSxL5JmeyFNEFLdC5XjAXqHk2Oj6U6EOFpo+bWxXudhY/U9inAIfXxXzJ1p90A7ZfFn94
2xpA2TKSAOtfTWELQ/3RIG63pnoVN4tcMXOFHe0P2Jyo+d7SHqHAJxLwvUmAzHm0vQRqWtU6gWvA
tLlk1M+dIHuHIXZeABE4w1G/7RikjGq9c/1ql2XJbwq1xoh8113k3Du9wSJKI/sXEzTtW3DHFJJ0
T7G3B8RBg5vSuAeQwUSZ+wApWKwb1A9Sbeo209w5yUObH1bE6tr1B0amH5O15D/6qOvfMLQn0BKx
JJvSe8fAgrqjFpQgtmulQtxt1+or6PII3IST9nbWuuURNnj5PJnRJeor9OTJ6heQdbLTYx+f1zxd
pryWWa+WMMT6buykgNnmBTZ3pN/Hv6aekoiKuBfOI0i270XBVkHC4RUbWL05gVsLeloSilH/Apfd
b0S3H5ML8WxfRkZXEmcp4cAzu1SOI+m5yAJQK7k+p87uY2glfn4fHCcq5M5KMOzdpJeIkAJp4Ojy
H5pdvOBwQHgg8sxBIbklsN5lNZGwKtIFrRohZPfrLkdfVneIGzIkbGyLs7ATnxElcqGySSZGoa8d
k7BW+jt5cPiM4w9jJ84GQhb2oBrpb1XfBGwWMk2QbycZa2IS9wc0U5oWgLi6Kj0EHBcLPjYzQdaL
6dvJzBHexSKny1MR19kqJQ/8+4VMiwkO80jSbMaw4d+fuj5py71U3VqQIfOlsIyRFQ4+Was8CdWv
iLC3FK59mg1LWhNxCPOwTQNWKWp2h1fMaAuQxFMHNDwaxvIGobgdGsuSsAr7uRqLzVuDqkuAd/oT
e6yl+p72PPv2gK2hC+itcrNA35URUtId+UOEZv/I0L3WPe9Y6LN7pOKDPB7xHFTVy9ZygW7XrSMa
tv2vvsWgxhBxHx8WT1a4UcIKUFe5bw46WjqWwMiMYFhb79Hz1otJOUbJ94UGT9q2Rgsd8IFNyBO0
oe39wdOsm8rCyF/VpBjAcVYHPB1G3+RND9LLsSpSDdEdNRufBhLw+qmWfq1A4oGzhbV8A3GgZNW8
TDhagWmDgOHaxUM2qXZbO++553D9SnR3zzzhmTrOKWHMA8D2eY1LSBWKoxPH0yNQn/nn3imcuEkg
/9tFQe1UIsexQBoDYO6rurUy2uXzXy4supMj757mWRO03YbzrO39rqYR5OC3NeWKkPz751mW3sj3
B7+hpWAInV6XMmUPAFDQ7uHED0iulkfg2USA8Zgg59ljtqZ/Vvb7niwJYcxGEFziHcl0joQhszpS
IkqDjCxxQqGTudojZtqiNhH6UrGfCnhsyX/QWw8cApmw4yRdc5HrhforTFkKAxEafdK0IH5n6AR1
FDesbEMvLk1ggBYgWeUu3tSosSxP3jnbvj+0A2a0SVEsawiq7nMqu7zGioH4SVTeZYcYjQqymODK
XAUjOcCXNtDnh37enaITwMsi7emN8xYfttN4GLUjvwBYIzL8Og0ddYTdVy2591i0lKGzM5h1AXIF
b2fDbYb8U4+qZd+c7GZrvsq6YdV1qBdOnjUQJYaGINeJQGCl8wYf6CZUttsN+cjeSAf0GKJ3iU+T
qCEYlZaXXomioE0m5hxmlHB4lw5iao2ONasf/16p2pUPXMPaAKT5cCkY2wFp8ph5WocwNyUi/bRQ
yViG35NhKSc+YkJGZkZwQM0p/t28LPsrersrTuNP4fBsNFANVwuBPBPKQ2GGwiCwR/Mlf3BUaOKF
gUW3q99n76aqF1PvT3+cF0tj8+eIQ5KQyJJKqaqg/wplF0LITcjFmTxa76huHY8oWGzKzYIvMNpo
jJZHbRm6/2TwWfQGvUbW7GjrAICDN0yrtFhUPsRS7nOZbtb7fFBUId87vI9ov21IKfWqEPlWxm3F
flMNtkVviuoQHIu/QSesYrGVb51jgIrCF2qDBFF7ymCsrZE1gi2GCVlsKLD2fZ72LPSVZVs4x5tJ
xAgxBSZMGfG+MpGj7WoPdhgjg48sa+8xTAEfvDcb0E2j4x24xOqixMemddw/grQqJRw6AmQArgnR
cyHcZK7eOXiA3n6CeRso5yTYsguCxuIj6oT3MUrvkipE65KuAhxmt0q8zaA+Y94Ufn6x7f3tgYPq
8T4xraDtwT7fVBPyyqZfks5YvWIkVKvnpre3H0r2/60+jv4szJ6fywxv7fH/jCtR4lE4LEYoSWqK
4E8PSfh2ptzMJ6kEhK+c46MNZ45pPwSEn1JgbQATeMcQQXn0pDweBcV+KwePNne91GqjtXt77Enz
EeTk5/8yicfR3f0gaffo48vZoNLehQV/50/+wDMvQspxNTxwmh+tenL+wD2L5WSgtX48nDHPinCp
jBm3rBAW2gzizpiFGwTx6QnlykgkbDwC/hSyxJn86YAMJ5EQ67H7/rF9kx3yuYfkbJ/fNBvLK1uH
EF0DXy9mgUZKBn3ETO3oRCOroAtDx7m7K86hdiQcGRW68j+mDoCiiXWYK8vyp2NcibXuBY5WTu0h
CiOHV5fDwuIc9suugj6E4DYOfifWP0rIPHoqNOqhzXM/ESxUMoIpnTBZkvAr4xvMrn1fV3YRmEqQ
648zYkNmvDKG0Z81qBLDCQdRKfoAUvvoayZQFsT5rA5lviQu4ZQHu1BkNP8kteeh3O4d1v2ymtT5
r9szwuma8BkUkQ6I0UuyXxXc//UKZBaEz8WfE51IyjIyC8SBhZd7PGL5s76uryV2DCTW0D9MSj8c
Dle1ZftXwTi0Q7uZUYkyRF7+2rO3GL8ymiC+knw5DIdarayybDdw9rhqDiyq9OU2vwBslXcB5mXL
P8VT+2QjgOSzECAUHhloufYHeBwAeJe+gtDQFGs9sTrB0d3aMNns6Y+FsgVg/3FWwGrJhuvyzHv8
kyIwaSi/i2KrX7pztgLmiij7DhfAoWN7MFepOLhjW0fAHmctTWazuyAo7bdg/UKpOC24Ec59CxCD
XfUYubgcji0woQ02XppSAVzPg7BzVcaH+G7yASkjxxCj4KQ2WBVYJ47ilYLI8n7oy4FDtQvFuA/d
EbSB5iV6jenF7FbLy7e77uN9NbbTwVTozI4K/M6tjy2v8yQxCvSPEkB3UI/H14xuMSLiQNbh70LE
eoQf6sTYlL1LlNNg/tRC7smE5/Zzm6/K+U9qyoabE5NZaeDda4z9+Fy+pxzeaNs6yyaZHxggmBqf
F21efRPVZQIAjSIkivKUlRIJHKiIW7mIzs3rqE+tS4T6PyF7jnkm3VzQKPIr6cnoTp953VJecwGp
TQkG2zUS4KW9AWG8Hzve/kQd59A9MNGDDtVURIIOsZXuCKJqR5OY5e8RMMj7kdJJ9FIFIAgGFV7A
9izb2+jMFxpOD0MfR7uRY1bnJxx0PSfVAH9SUDpGRUIc6QiZd5Z4DnoqOqMPNZn5KS61Hp91nX8l
bPhX6van6EvtkSI8kg1lnByqG4eN9DlBOA+5R2zicuQuHihfp128oPmW2M8FtjFywDn3ONLJc5e3
g43QgMaz6SI4kk/jbyYUPDb9GSEqMfx/8H2nrtdntWwq3/g5XjVAnMM2Vq23m19DHJIRdmOSwNDs
TrzdnHGDjoqS0ZsMw2CIJSSn73yaL1z7x95qGLtCGBMKs8NTZzP1h0A8zXSiIv8edX5t6U0txFiK
QsXjrKkedIyf01suTnJ/g+NtNtP6QJhAt9mWsYcrTbm40RAyIJChpZkiHU6yo7QxRkX16Xi3lOrs
yQnmzT2PxbOOwEYkcWnZ3iF5bBBdQIBYRZkRp2/z+2fxPmLXCh0aFU44o+MqmuYxmj75qCuBMv1r
ZHrkyTaSBUvpyduXfuv1uOHa5/ReiWnITURjcA0z/JATc7xF6WFNFmr6NKPqe8NG1o4x8hfZ0kYC
/T8JT0ZlP8NwR2hzCfVom1djIwAsow3hsaOCpF0nTl69XThBNnOpJEaMkTGW1TY4sPzImpTz0y8G
ZZS1EkWT7IO0BtlKo+739+KGHmcMxnBvtX5/nubjpzNqzmO9uvLqs8aJIlla7F/JpunD8w3Mjq0/
38TbQ2mBsOz5iwNPY3eCGEaDaKpELZBwjIINtKtA4YgUbMXL9Mlm+q+X8Q/IjfT0Yj9qrOAaKv3z
dfXav4S7oCy5cWpqGqGjXXZUbR0TE4d+8ef625sHv9k425fAA58uMyhaXPrUhg9FtIzUuyPYSHbd
ycga5emplU85MiLgmZiZWosObLEg8GnMgcB9YZZPucYl8YHvL0etuRTub9P1cgz/EZ8P6S/w7CGm
VFdlX9NsQRS0e+Cy5R1PLnoKwkAoan6KlTmuCMFz3wVDaJPV0jat/udOnLmcpyB7NwSP2P77FSBL
eAd9o+txI1qpv9+ExMfUJPUN3OFXOTQt1/tNTw2cPSyo3+VATHAy+FSRy5myOKhNLnm9wAOtk1aO
5iKxOlgfrQMbo9mwSIm9CeQshxZXhSFybq/sCUynGtUbBeHeI0TDsae3cTkQHbe6G8Dg2GA0E43x
njjwp4SpQEI3kwAbCa2QEOWw+awnorfdW4k1PAUkLKfDiTgj83n47K69TjPgOrmNE3MqKFNgmzbr
AWxrkwsY4Ft879HGQVIbHhdP8plmQc5sBqehcRD30Hqi4PTCatGan/ycJNKOES7rqDj6icY5Hnvy
GMaW/7i1/nToRRLgZ1K8ioiF2SeFPTMiwMG8gfztvazjTY8ym1T1Xp3CwrVUUUfV5SknfpGHqOmF
reMF5sYZgqx/KRbI8BD1epil9N+n/4bfXQVBVEk3fQAQh833UP8qPooEqI639yQVMZyOmTG3z0j4
EVUTt+uIAm5/QnlCU7XSiHVFmW/YKfPBFBKs3Eu3MMYceq58i8lS9XmUOgUBHV2SQt5Bxpj7a/zH
UZjoEHZtNbQMOAb2SszUJMEXO2MF29Pp9fJy8S/DR1B58fkq20PymKih/TRZ1d36l3RRc4sNNrEU
IyfQii4lXzZ/SMKtoYshejj5X6888ghJ+odHo60aPc5BCQlw1Kbo3bJ2Qz47lypxfH92wi69hmn0
aE2PGaf9h80+PLKJfyDm9r+1fuVWhO90v7JEncBJglLSsbcShns7Hfuje4u6dNS/j/3GLtdy5sjx
mr/OB1yDT9V92sJiPFuuBoxBsRF2ABGRsRl5wVyIhG+pWRYpqaqJM31gu7xfNusBapQQbPCQ2BHp
XlWEJHNB2HDf+zMrl5PEvyZE1p6BjJD0259CjIJYrlyiGMUB+6PLgCWhDpcQlF8lv0YGwSmbX9ac
t/8E6Ri6AFZ7+y1O0ynBRLMHrZsRtPJsV5vXTXuDHCcgyvQFJSLfSPjvUshfHFKmE2r7NMA1RlDE
rRJ6GRGsbGtMZxY0Ic3kYizeFWkKLmyCSN875aC4HF70oqpZIrFcgc7EO1yNXlrga3f9uOcVPdmh
itTRLaVKg/ZEvDOIISxuEeXfCNYJ/CZOsy1lYBtdvxgYYaP28s38bYNGN8cj2gPvwA1thdPJdlsp
U9cFHWrCdGYhjGMepGr6aYj461ekvrny3HfIQIZlca5M3bdRv8XM1BbgXFqLJNS6ZcNfhoF45RW5
QwBnJFiAt7vNUULCh0q6c27d68RIxrjt05prgLqGsEA9AcoUy+GUA3bZ6HFy/H3P7z81Zekc7C8K
sdY/N4UaKotlPJY5XFS68EUx4ZNRX5RfD/fojFx092K4qTj4cVr5YOyuBnWHOdO7rkXmV3xm4VKv
MNIda1dre7LBIM++tKA1PXQIIjLJKp0LJNMehR+cIld4EMITPrntSkORjNaPBYVIXD/0Bkl+fM07
IinD9tfomMHv5MrgDiqEV9Q9A+t1wR/zkZ8SyFhBjmt9+Zb8MQDzn/o0fYxPzcmHKHy2FSqMkz4q
zFdhtm4TSWNerC1SX2IpF3vQnG4+4i65GVj+3Tvsbs6yuAyIFs0Sd46mMxfPwxFH7PkuvsRVhiMk
JBcQS9us/h67g+GPK95XeERVCaODYdNiO/U3Jl0kGt+C5lrGT4p2idJELVn+wv5OVdstWXyY8soY
16LgtboUVniE7eE8I2ZMytNHw1H3zR+Oma8fGgYEbkWDgFjvc+EOoCTpOI/nVVrUNtOWcAu8YLWq
cI8BQcvruumKrxeNgncaMPInilvWZvBZN/077uSeYrWLd4n/DhUROQOLutB3TgeD/skhs5jzazY4
Rv80hJy8cpGvaplcXY3ZBPE4e2l3+gVeyvnTPFakhcJ7r+2PHawpUO5nn6zIW/IUH2H4Rh54e7bP
2nZZ+PJV3nMgVLR9W1+ExyRaEeEUA0feOcxXywuPRQNIh/nRh01spUiEy4x5Fu5GM8hEnp8+C4Yl
C4Gqop0REo8y0PE67oxnmUin7LJZGxo3QNlyK+lhk5YODJUAawG8oOLXkIysdH+BgukbimkjC2zH
emRBj2/LYbFvkULk2O7KXxcAjgWdNKGddKQslilW8Q9A3B+M1WICF3mVAzIBLsROBvkd7v4G6Vbi
df3vLdc2tXYH4LUEph+LII3Sg4aZiH21+i0fYRxaJIgPyADx5M0oaNl3ojSjz37UZDmD6W3UlhEf
tqwwfI5WY8ld1WNetg+rhicPolt+VIHOaGjhimG6Omjhr2y5Xle4WNvDT5NwRRmecLt2bP4rfb4x
Dn9ToOBNF4DJE5kb9ZaTKOFmyf3xd3l/ROsKNxrC3pbaOT7hXUvqU4iMWlGA4CqYgd30WNfNnTeX
feavnJ45kLUCv/FLpYmn1fdhtxGRVR+sh1Nq0jboAo8Z6rQARz23bNMDgyUfSgIu0cmFAcVQSAYX
tHY7T95qaOc+MYPcUzeYmQCN981TbYho7VX6cJvjyGxS+L/KhZJKTHKZdxiD99xXyTVFjd4rCH/s
eHiT96x5nGH/ZwP2FZEEvmeeK26YQ4tGCLp6T4mSc03ePuBkLMsCTAFvYZcV02rNV3N3kVOXEhvL
o5NzReu9WU6n1lsWJyteRm3SEcoJdvqUh7H8YDrQxCcAdPxzI98zaBExV14xhdpzBGWgWzBiITt1
XQOoQW+9vFgqF4iOgYu1RPSZUyIq2xBQ0TlJDzovBfuf/f6Bs0tSMsYAPsWHs4a2UCDkN2tHgH7R
eE7mJvd6jYrIjmJkvx8FSZdSe+Zxycvz49mj6/sI3jmwc4qoj0ocJq2ahKeSskNIO9IyFBLLMgbj
RVzXnO4VuR0932FjQ4lC3MEYXYkevVingkI2EzLDL7HP3nKauJeiyVJ30jiZNsaTwLjclbSc0Dku
CvGR/ThjRiHFd+lzwJSnHN+i0Gr/igFlx0W6PXgI2nh9ChQC8rpnufzE1LPyxPBaI2JaCPGF1Ou9
DxzfP0mV9QMzZb2oz8HchMobe2Y3cjK9WygCa3aLFVs/D/KFe7oeJ1g1FxzK/xJn0UuuFxkZFHeK
uQOw+x9DQHm9uBrMWte9CBEosRZbCGal/1zgcotJmDtCz1K5S6puu2wPF2sbLM49DjOPTbM7qUD2
O7yzfJlexih2E4KSeUtcENLJSml0tOlJPR9koY2htdLq1y/+iSxRNdKvletIoqW58KoPN+dofDBP
3B4c2mb2DbtYM+TLcyquPYkEeVcySQSrqbM0Vcq1PKn8n8/lQKou+m1krQzmYKk92KaV1MkrYV8f
e5i6qJByiQWCn4hPrfNl2EbDYB1MdLDzZPx0TG7amwA6GI5FKAGRK/cP0VRAa/s6CLgzXpfJVHrd
ZYgnw5nGgjDUVIFrFnKWKQ0qKW92jWqhlaYGcmyINrarOTvjdZ5vZvYy0/RCJMQDdCr++BnKgsy3
sg/HD3plwWDfAkdNqj1CmMtCC2Aj2xngZFqNq9+5sS18JnUYbfZHaJyY4UAXgVXBxTUpTg5+YiDw
kjrcid8PFl5MYi3DRIL8fAcYX2HyfccMlTDuf9Lo7tMXeEmhF0ZHp02fILD5lPbQVsW5ki6E0z0b
om2gV25Bmukq3mdCiCUO3NR+s8n11y1fgmapcYGfeGK/fjgcUx/mCmOwNEoWuvl2EdN6SlrXIjSt
TYXTHKJgtqdmEAA3OuFVsc0xLaQJF6qQdQvI4etn+v3ckBiM+HfOnIZCsJrFTKrOtFVTo83AghBW
BNVsON61hTwcOJOmTF9Nx6fRoBm/akaAzoE/2qaD23sc8azJG68yf5+glYHSSttEy9jZ565B2Vgl
v/BrfdQZC90Tii9dDXFTJfrT1vawIbez3R1fANayUEs7TXu90nw3MgZu1Gc4Eayf0lgV1Qsj3gPq
nrYCWfif1qLoSnlucplIwx9eMIyjUQ2uftccY4CsKEFPChj8q1OKlrWx8W9CSzemXzRiVBcTzT5W
tO0Mw6wAhcSOeJqobjuGmCW9da5orPcEYRdhJC0D63A6bTnv30bxXWQK60SjlLvx2aMrWxci7s/u
9v25n0y/8082Ns2Th508ZyVjPIDySX65yGvQSCpcxo59/orrJOEIzT59kMuvokN0WA1Cggwd+n6e
O4DxdDvBNW87EijIHySRk6T80R17JAJClW0fwy6LkoOwGbykff0TKvCIZ6xzNyooTkY3W88lvIS7
lmPxBpohMZKTx17bpUl62Mp+SS0dicpzRjU9ufpaqTSO3lD5cnf2uicgoKJDObwKOaRkw91Y0+yX
XEC1XYcDY/OducpQEM565qvfrX6koHgANJIXxURvn0XT2qLutlsVIT3aFqoQPvsy5+k6tiV33y4Z
MbEPzLscmUmlr05OLhlRhbTWQwRqiDYlWqrSgI1A5fSEsEASwL/u/VxDTu67V2eE7R8Xg7nUjyot
svpGjsdPy4NWXQZMk5axbt8rriSt1gUFMbT/+S9njTOmcJ4x1pANW+l4SSnnobb2YLHLS1F7Nsch
BXQL8koc4ZUyzUADLSaTkgpSa9oqWQWokxF1GXrggVvFcPBPkqOAlHF3RnuarB0xPB+svQNVcm+D
qLnRWGvk3lo8nzo1H/HsAcibVW2MMFR1u2xbk6W87xtS8rxhxAPSWnaDjpUhv6McolEx6AAwj7N9
TdCZYvCYtKXdvowieRvNwtzEL9z0GS6cembnC6NL5xJmwu/T4FsUlQq+054PRUIkQkRAIB9no9YE
be/65N9HzO1sUmVo9lZs9KfhxxVaF00RK4G90AjifWRq+3it3g97aZIJRdp5FDzoOVUL99QX35Tk
h0Etdl+wKUb9PJa9OxSygvaLn9Vfm6PnAGXEsON8lVl1gHQ6xIwh1tgShwno3IKqa+tYIlVY5Zzn
Bj3S+myIY4JQrZkD/SEc+cafhVxRoAeSQptWQApOnJM0oMsspmHf4L7GcasKTF5/E6yhf8tquKCT
ODGMPWMCuVKbAvFioWMgMaU1CLYdxIfGFoNAiDdjdUVKSoH3yFUPQi4CIlK17uxiN1haFAjEZChj
VLXM4lxmVbdkm13U/FW6LLrvAYPLRGBQr7jrMh080Ns0AVJB1ytK0X9xYPyWSlNO4o9n9o7M8jZ8
oVnk1kI3rynrj5wk8D94sa9mIeBgiynRJ5fnR55oaEIPWmDF+oDx2hp2KWvNCl5YjT4yVw61mhmH
TuWCJqpIBIS/VVGPjL2x0qVwmLznxa+0EYtk+qDXl+FwXNBEP36KmhSeQA/7eZmmI2aNgCM8K8gW
5TRH62XRat899xWOhUu8rbvryAAmzq/QGBBXz06blwRVwWavhCMSVsMe3IPiCB+TZKwQbYudf+yX
qhY9/XmWkxpa09LcBvcF/NOX+oFaoLjmw/WTaWbZAsgY1xwfXj/ldFxz7HhMgzSoiaLgNAdUgS6i
fm4PZGt/lNqCHBGWu38dETH0LEzVhDyzH79P4rRsPvzq+fRZNLbiBPmvPlr8d4CvXcxgLazLGLqw
7bXmoohbqtFNYISyMkllhIFKS7w8/YQzp0j3sRLJLU87+vD7lnqJbKigmh0v9xLJhQZ6vclauWQL
nvYvtuuYiU9TSMA4IMHP3Ty80q9Z9rkOkKmMHlnHW2Y3ZaW9BVKlUhDyAykMZvRUg0U3H48ahg7a
oURbSdl0bmFuQ2lssKX+Dn4RMAMgZx4isqC5xb/6EzutQyfjUdew/wEVWVreRvdA3yeek3LrxbQX
zXyn/G7zB892i2ozccQBx0ZsTeaLRe3jD7RszvTn0BIgQWVrAXt44J+tM1mcatISPIvsRYDuq/py
mTv0rk38cMve7Cl7feKFurF9hl9l/TZM9SYrpCs4uycfjwxzuGdXEnq02JLZSjnNb/TBrz2xojQG
XPiAMNf1hzti9KyjDcEmuf+wsqEeYyEyBeFUKRg+HBakrpdKvBr3QV6SbqwO2yTTEEXE0WOGbBab
GRxRfCSMelnElL8yOemmjNSwz+Hl1YVQTE4EzcxqbJPGje0wGG+HX7uegVlj3Ik72Jd0EbLKNbEu
v8haJyrSyElTUJg4mVVyGtrbPJDjbsezBcYM1vAtedGID1xyffKtegNwSjWJVCTXXBv+JKDDdOuv
MoV4MuX1lpzLBSR+F2yniD5thZ/6hyMRuw2zYG0GSVdob4SWuMDDGFdmEqbh8kX/OglMFxI5uDid
lKdeiwWsPjiM7Hj/Gj4cTd1QB7IwG03qG09Oz2jGGXc8DJ3Mx5YciR5zMIuMsrAOPNCSe+C8wemz
uABbdGlIwPrcjMWaxsnV4CFukhU8v5rAPBV11jQLgy59fBE0GOYRh5A3u052xOY9KkQDxwoa1Rwy
wysckOJ6ufDCckbeIYcyfYJNqcXwJeBOfmjHiU6HokxaN9k+nqKyKfSPHp5oUeBsCqRxyKdhdsiO
p5Mh0gbHf6mn/GOu3q19xYm+f0I/5g+YMSct3HoMC8sDKo1iHAYkiQtkidRo6/CRr4UFIkJePyZc
M+K3xqrx2L7/7dj9dr/kAM4GCaPEK8zWgschb5E62BeSXqTNXqExXF2wg1UXsBSwtSq5gx+bv7V/
SDEA59f0ysFd5V5qTPr4lKcBcM2MG2Gysu90q+0OqfvPnO+IctJ7ks7nMr+rzJSGP4Fws9zHPDFF
nwivXaA3FYLZLSDuGodEgFtYZe73HLjlBmcWTqYsnGDXK9gdyZBhMqQCN/7HZgwJrS3ALosaTvg9
JHxK++KgYxys9ZzVOkkfqJrR0oR4YVLyV0ORYfxlShcW1dkzTGLROJOL0o9Enq43i1Bu5EX+nIM/
E0UtUFrseJymUGXG3EFUeGh+YnGTb5nscwdGD25BGd/lLhISW1TrOAZ7dlJ9E4zukrsPAYNpDfNB
M8X5mG+KYtwAnunst/Zl07Q5zQeKuSq0JkgBd+crOzpw0tMDFNmwx6UfZe/kLHRyNFEQk9vlIiOB
6jyQ7vvHkulAHqRBGgGqGckGZEBhVrdJK6EGgJkx6w9awg5B5hFYsmbVY+wo5QYlOWPqt3rPEjze
UxgTcqra6oGNW9JrMc1Ep7OZG9pecMYSUm7N2IQEzIwzMIWqpsIzpG18AD/XZa+1T4EIviPqNQEw
+B9hnnFReaKTUh+m6qkLe50FnDI6+2+BLGa9udp1ZjqQ9I9csgz7f6xCSwPRIz7XQcSZfI4MRPIs
AmD0iq7DY8p8edE8JJAvNtJNc7MajAMDgwmocDpX74fSjFDVcTNPNiErGHPPr90+ytDsRrVDutiq
O8gh6H3us4f7xllK6zl5Z/4R1IA/doIjSMklyDjGuxFY7HBvCzxs63uwsX64UOU+RbNVTkxkzoex
bqoDvv3BrmzCJe7Ea+Zb8QOUQKewLKpZpTJo4JAtc5wMa+tHfVCaZ/cfl0Pl+aHscWmaOJLJ1Mle
bj8RrQ7DhUFbJVeAQmEul5rJziH5OG1AtZg51v4p3YpfHP9eitZVkMMrnwBMegjBckQctThpFxgt
o/pFcYez4kyEClVxrKG4CIc2dPytlqDbU9sxHR6bhpKkieke6/kX2Ar2AuLOS12Du/O9Ue+27jXY
QtU7X97QaS/pzP7Q218j2B9XDwldn8ji22hYhOl0IRK20D/vX+8FCqPebXVIrOhurIWQ28RptTqq
jrQ1tXuLchuVy0whgy3CY9QXwXpZQRnSCfKP9QQSgtPhfoZveLbPhTOwjPstQt5nVQOzmdSbu9k7
yM6Ldn8g2GmZGN7jtybQeA1QlQPQKdar1aiTsud5isf2+m5Dshs4LE+coCcoj1xT0VyFzVnkzt8s
YjFpf/Bgdp11sfe06s1J6X6VR674H4k83619rTqDd3w6nByLd+N4JwUvDnW2G8LJHflcOr4D7C9/
2DdDHpnkgs9trqjvlQQqAbWyCZ9EOK1qkHbWB6UPvbebSnwcYKFHsP+2pc6i9cf/ohB8PzG1utpq
B/n/k0LbMgmAYtvYiPLSGzsTnMUkLfbkmPZbgRKeDFGITBgSEPzlvYGrO7yXudS+0/w6H42EmhMj
2LXRs30Zy3/Qn8Nn6LdEuVV12+cqwp7wfjjqc0xYxjxd28BEZWZrzpoYVrnbhaNZW727w5oq2iOa
dRrLnsSCR1nxv5KrQ09SpIToaulYd8x+pPc9eP50wmxbPc2NhvclsCNjFyhE9XFqTFQTh3+L/0TO
fU8dfOkzx9MHnFrUqVKeizAQ55qTZhh19/YtIQk/HzJa600sMS2DlAwcBh/85du9DWkYGBoIZG0w
wnzFCOMQShYdHgDAvjdh2kFz4b1Y2Q80gO8Jh1Pg+GAtMZ5jcsg+Jfo4q1xG/4/2PY0EP48BNq2m
++33/I9Sek+nzDv2cdCfQZ6QelNYbMZS/ZiLYk6JJ8t37cbdm4oI9VtVOpgwTS86yUeLTb7oHz4t
QYxZ8aj0eWN/e6RJBaPb5+y5AAEILqvIf3V9zCTyXLCMyc8fScxOOYZReoigIvjQF7pk5DfI6IAv
MlulmR2zdAlInTPJ9JsbcPZUbd0prCgauFeMJizGm3tbmHeRow8pobPcN/FBLvPd1kY8195INrVS
xqhbS0tICWx6kuMSPS02lHQSJR2Nfbcgqc7jaxm4hip96FD/uw7bkY9lHRogA7L/KzHpTcmf2zIW
BnJzHT9lP6gqGFTBL45Uptnfviblz55djoE7B36Jqf9SgoQPv8git/vlDqMrZbizT383YHdYj0fn
nav9muO1q0qI+nk1Goo/v4AkglbabmkOQrNq57vtH+PqBbuWH7m01yVY1/rrZ6CV1N4MGV5pfCBy
FRYvFKEzmvJxe1ohgyzPf7GQTd93C2Hg0Gb0kQgVoKoqJnF/3UGGL6oaSGB7cTpLMkwIAAHXWRLI
UKGWPV5WVJRjcACvqRxWX23i1B83C3gLIi8ySCa3/2TtArSdCCaI4QcyQSx+Y6QrOxvEs2JJbuCn
ODKxy5jw7Hr2qkiCKYhf7IKYY7oFlS0k9k3fnb08/reugTefxPGfeyXveSfIJVEivp2VxUWCLSVw
/PiJpTh22BvlQ+pElT5VgkSKl3WYuK9iTvkgIaaQh7CmLPWLw4GU+I1/2QKXF271bH7y1geNl3D/
pB5+nAKqJ6rgTaCvX5qpYVnjNT4jkQ9gQZWccWDHGQK04jkRukgycAn+XUcJuy5irT3cNIbIBvSZ
FM3jjvL4uaxMHMXNjWN8N6TnlWMYPiDLbvcg66bpo64lA/vVxzIoNRCCQLowHHyUVKmXm6azUk/m
8/QiU3UvLGd5yvEBKTJvRKuHpKGcYnAxmnuq1TIqroFnEpwKGxBpDY7lDuvdyMXNX9jxBMzIyTyU
e1LaM/O8zfltXATJV072RZuVLIIeuePKrf89yL0rZsrS+G66uUYXMKl269irapZqWlJ1VCzbSiq/
nvi6pTYHKXhXlujtsuehmQ+QB53y8bEipTKuYOjP5h+A9sguvD9HLyV3f51Ah7Dwsdr5F4rphbpS
OoUs9FXaDRSx7KC1Ku9qANHU8h4JZbR65XmN19EpGe0cOUHyDz0KXJLJZUZZpC3YvVOC5o5OM4WX
iCCBYF2gF+ey8UEPuV7nSwLSIp8m59yVJR3bxqEjotO4DldSk0oc/ihyFSWpiOtt0dxQGpGV4bNB
N/9vLMipCBWssWfDreeq0glT0/sno1iIKziV0XFVrmSO9PR0ry6RDrWALcZYK9kI+SJV2NTjlnYJ
OEBdFKIeJrN687pjicu1KhGcA6P1GPQZs83RkL86Mb1O2FBDA0B+H7vENmK+JVKIiwCLwekHivsx
hGPrNcwbGHFbtiq6TTESS/8a3Vx/96aCPabI/4PvMhFoX0sKmxCYuxw17+VoeTfUw2gdS41chM2i
h4cHjJALIibvLckwZeVS34Am18/rB1FMnT5dg4qeWL8XHCmZ1IAtf5iRjpBYmZAPn9WD/UgqkXGw
4LlxByXbJGxPOE2tMbcOKsOprnAJ4j1D2RmcnS5jg2Ydguhirf1lsYmcZFDhqXJ2WlfsbWfPdhPn
/sL4DWh09xh3+CUfeY/+tIUXjuCiCspts+8eBIdYSmgCFjTAANHzVoSudEfhEnz4IpmTyrcx2kih
4zM1gHiN87zpHFXaIHXyuU97HFoHIS5hzo9dsKYWNivm/WgB2thfjLo9F4NyWq8pSfSZRMYUXaUd
mI+0yng8zVa0rEeKIYAm5tqv468RoxAlJKJKLJwbHaVebu0Q57dHQo+hHTXn5/SZ8f7SbSIUZmtW
NLoi47tI1cwrmt/evIswISGMGx1Wrx9uGfLsLdJ1MBRS8oIO5RqoSgKYjdMdZL5GJhE4bxW6u0gO
AL6OgeZOvH52OC6jD1A8Iuxw0IA/y6R+oT+ILZA7L20MUPYt1NikT1RfjLYcn1PXv5c87zW5Pc6e
SDmJRXMeDMrUrr9RSwax15MLxlVrKJ1OBNSZgQihuvAR+HcHb6qX/RrcqIVGI3lOyeWHlf9r+SpZ
TiiSzixUomuffGlhGj/0WCBn4GdYVUyGGjQQ2aCOKpdu1CmI1fqex5zh6m7GfE5imH/mEI2Yrm0m
vbQcKIsa/9nGMf3TrsqL6iF9Yrys5kktV861sWs20xzo7Lg5rxhlRwL+bBHvm2L4FWs8Sv3oNs39
DNPddZr6dxjlYzxbiF88bZt+RnfiOCj22eAO9bGnJ9gYEN644c8U4P8CTWnKGOjqry41CWFtCdb1
O1Mu8pjTWO9abMJkKvbf1jUXFVn5xAbC+0ucyLxxLopYR6n+6ThzoTlzG4IXqbvYEfHzLsBF6kb2
3rnYom/LvaMtdQUvplPr2vfeh+CM184+yuJD1gz+TWwOg0PxfR0vzElEm8mEpVprMjFYqkvfTR29
85yiCO66HRVjM13GwWtylF6YpNuCd1Q1ZUwJ3kVriljrdtZ2k4I73WHsaQAMIjQf0A9f1g6YFzN6
pKfsoqNB1xmHzmp1P1UUJh+mKEfvCrpEsoKmEy9jPNCHmSBmSvpIx0b6VwJhEe6/p9b8QTK+lsUy
42tjd9fxz1ORopUGx/kzfjJaezxQU27TsLDyFosTJ5NjBZO/zt4Abwm+4o8Y2FnxPj3HB1zXXbev
RMXxJC4DovBy8tFShbKoQvrPzvDOcOdLsmuUfa3tD0IuVF8oDQS18ou6J6hrKBOs6xMxQvRXriZs
bI+eSgCNAt3S9U3sTAywzujN6SLZN/ZQH6bc5t54h750pS63B7x3xk2k9HAwKD5xgdVZrQpH48jD
F+bnjzhzl6bk4UuC+ktwknbszH2+2a3zj8XOvQ4Vp4Kn5MqkMCGXsbnMCh6saUdjqZ++hNyZcy6r
Y+xuVyDJ47Zo+NeYGyiHxJQNYvesEwxBBeiuyNpbM3Iy1zapolNoSTQ/8K2ILSl0J9ZuOmlNjQaL
20sQ/Low1K1qSRd6SmmaIJ7/jshqfcngyuwbLrYnWAlZNXOP+n4y339SyyEx7DrZCzXzJW4zBaup
a0FIpoWRLcknCB2dx8ZBBByHCXta0HxyDNEMIlsDgHJIyUO6JVzy4bNKbcceEi0Ae+W0SVvLwLqg
pwtokfu5kOD7Xjuasw677etf4+KqgcVgmDSR17/1QwxtYlQhJUfGPhmlNnHeyb1WWU9D2qtc93KE
K/KLy6y7ceFmvPlT1XrMZPtScofpjyhs7oZEfXCrHv44ls23NtosoGa4PEf3XANJzKoeWfiw8iWm
j2v44yyfmSpdlqXPqM+EjAgjaKPvW+ZLo1QZOhWuRgrJeqGk+Yn4Y+HCs44Eh4jCfLbcBN+wTqXo
U6RW+emAIdHDiybGnC8gNvYSdcc+RYa+A95DiIbfd2jgz/exQK5MIG8Uvj2GADUg0fJSAw0AaYkt
Bu7ySMUblc0wH9I6NE+4JdpeSDpLOz/CFZ1OcAkZHbnNpWXPepujZmVdf3uUQ4cCao7qhXaY8pbd
zfIDIe8YKdEW8m2NRaLDL56qZ4BwPXsEHKBeW2sDpthjmVY8h6odCff7Bh+dcFhy78LICvSgqiPK
AQCDY+YwjNYIykOlUX4deZ4F+sM5O732k+ipNS3iU/aG+9lbh3n2/hd504Fhr/q2ZaMaKuBEJu3/
efoMXpwdqn8f4elcTmOvTvORNO0UJM0/mqmkBy1KXHKdmmpU7/ac6CGYjy4IEzAR7vndy8hTw9n5
4Z5Yi6G4BLKOg3FrsPdZlH1xf8Udva7Llw9pMksFopbl5w1rA0KZnQHSfKwxzOprm04JclxMJK0W
+FaTPcaRG8XXMDYoZCuMWDsT5KXofXcPMGtYHiqieo5aOIrsm3kxo86d7nTf0Cq7sZZwnIScEFK/
ce6y97a28jBoCKmBZf4F4+tfpQxchWGqGN86n4vRvMf2z+tkU38E+xZiQotQl1Jaq/3MxjrpWhgj
76GaXRclSwkKtO7wc8C/fNKmyaej8vJtYPH4xgTc4+f/GUc+pKUVRg3xSRD1eVd3Y93DlTuaL1YS
JQfXx6FJMyvj8MPR8TIjFq8aIMgFq/zAVeFCh6rz/AqO5Al9BXRY1T7puf4tt2HRxBECioHYSsSJ
a6wwskftbujZTBoduoQogWwOFXoykeHz7tglB6sOIxGmp74IpCOlAPPGzQSqqtJHeJUOW2HEG5J8
r7n75l5G0cA5N4+yUTvCKcAU87MujTnOvKJxhaPc2J1972RRlFotTSqZT60B9XLhJQzgoY4UY41n
Tb7/YkLZEbdFGoXDB/b4CPK7wyeSY2GOq3ErF5QJ/JyvLUN4Ctn0ab5UwJpFh/V4mKpfHpDfPhIV
rYd4iDDZr5U078oIAmOrV+6+zGhQXv5b/NsA5HrKpMYQ6X+eTvnPMb0l90mYS4IOEnhA6+LzU3NL
U5ltXTcAXiVpTGf9Cxj05DB2HCPJ/fTyBGjW+/qY7B86+neqjctH/wekVn/qTS29iyNjOP5hEw8G
cH+/fD4+h/hxk5idKm86aJJN6ijam/KwSF9WeceZWFGuJiP/97MUpnYVqZ1MCKBuMygmxD+0VtMA
YNLCq1Kv+riHhHl4+FaMvBdYpE2FVBixifqmBB3P/vre8mslf3kvV8EUUY31iD2WuhGJskevtnFP
RCg6ej546YgDmjZ4Bo0CIYG5gzb5mJbGQNvB2YAoxPd0haeKbnPNBDCGx2xq1NT+855BoqImb8kQ
7eMfapGcQ91/cGC4O9nZ3Q0BECxsv8GpuW8+BvM5/k9Dzlk2xQe/BTzG5s/SvlLZ0uHMP1nYtTJw
/7wiaXgOtJ0WLTwdkltBh/Ei2uifT3QBXWaEFXA9vA+w97KSaRdx9Vo7aAPwLQaGZVMbzyauynCK
5v+S4ZYOSatBP5kRUXLYJWT+UAYuPKzD1Q5FVFP+iBNOy8KEYay58ydWsIAsw1AOzLKOYdfGX25I
OdhxTH/4xoF0ehJI4p7HZ+B6tNemXv0VX3R2uP9uNHZ/o3V3shZRJV2zD4M0sQuk+/t9hLwD+NYB
g1I/CgPBtJzr/w23p7EK31Id5k58/1FDxyaxWxRCpPip96CerYXbKyCBANKp0/n2N8dmNAla5bo0
5UVdUrcqWW5qRchS0uFPpwCbOKcbca1csrq+W7lGRNhj1tQfWpZOrRtq1KGCLKVG6If48XG/ibl/
tSANiP9S8zHX8JK/URVdxTxT5Rc+uHxg8jpGTi6VnMfJPiYLDTlHeDFP5kxotpKGxChAR40DoR+f
VPPUz49kgkgowKrWFmLuV8/76aDrhI/QzjMXo0isZJRnf89NbBrRyiQ8S1fbSmy7I3ijqEwadEdn
RaL0mzdT3a//ChrmaP+46SwRqgx5RkEYLNDXUhGkVMHikTRlPYBj/GWrqHxItKITPLkJgAWWPC2b
a3ElzabNbQKnVD8/VlRgm2pUDHFHDz7ZMC1cwWoaNYQIs2V/php0Hq/UXIXfAB9CzqN5LBlJn0GJ
KhBwES6VKlRxT33wOU9bCNEHAeFg/qV/cTIw4T+hNQ3NABxmb5BoXW1L7GiTNqkjkS+UcSjenzLC
0w4pC6oNU/kfMaFUjeBUoyhn4k/ULXxnkc0Sfv4DSEzJczADWJhLTlZCmXcV6TAYdAAxZxuPOU3S
VRw7q5VboU0ZySHdL95NsENGCRmVZiOoxW2zmkihwFcy2Vay820y/YF7Bjg8rDnidm6UGGGYVPNi
Snod0isLITMBzotlJKcLm2QrdyKW0+WOO+waw/WPHEabBkorYOIgV6LbavRUjDcc2U4mEbKudHB1
ODYWNgaO+vpeITYEtFkG/GtQU1VcskDxTcFYQkDeQes84el+YiB6RFP6C0R47danKY8kMIjvQxQA
/vaYFBueyfM21BN5kTxPutRFeIDDkESLx7cCwmfVqT1799WyfqIf2inygtwpT0q4ZSdaJpb5G9O2
nMLs9OLhEHeP1saFDIy0sWlUvrmjKpgLRAQpA3eBh0OKygep238OsDX58GZ3oPbtJgKXCz8zyEhx
g2npmn1XS5LIqLPig4OheHXU0imNUxyRdlqcWq8pBuKP1SAedlu+ou+ZnZYq86sq89mFQNiI32LZ
e0B1S2dx1M+2J1q3HrsNvZJ4tCRBXjP4wG75rY4ByHqUH2cQV55AkecUw6Txf/RySf49uRmtItzM
pEoDFNuwuIiIlzPkDCZHT9+nvBxKRv0EiS6V+TxYb3U7JFa3QDpad0+2hCvR0o06DZ8ChKLT0VCZ
/o9wAfeVCb6FKk3L/JcKMfzwdtCaq7wHpg6uPORpPv9A/gClSJIhPQt3drMBKE5o9Z7P2bmxVgKX
NJ4AHImvWQjC+lhSvRljufD93C6hMVVjY5+AMQYQyKDoCooHcvXVgIEK0Z1hkOUBvy0JNWWs14fe
ID+JuaY0N3y1AYe7r2RH1bCgNpG3rZIbZ17xLbkw7R8iDV7VgI8/V133nlf/lzddwerL2W9o1eUR
g7zbECGa8HDIM2NOBGR/splBSwcNllXhcWZwb8dOOzeI5cwdpDH5LGJRlymBdXCGQzOAkMeF6+iL
hd/qSMOslIhiHeWj3mL32NeOkljQ9jKUCJVcJ42KbAgwZkXWMug+LHiVc0d11jeBYU4sHLZ7YmvL
8r425oQngb4M9wD5CANy5Ihlhq6JHHnZJ/XLVoMbSSaPgpzbZ6oWvaiqCv9Id8IirpbcOJR8CnL9
i9uEW3h+7g4Onm3kOG4lGfRrW0kmLolwURSEslt8wOO5eIDkJS/A484JIV6D35SKv6TXSjDa4l6U
imbkl8xTL0E9kq49KLrxQ8ZhpoqFqjQGBlBLlEHZtuPU3bpJM1rS2gQTe89HCz11lt5kvKLEYIGr
vY4tcGmiWTeNmfNENQv7hZNBz/1JsBaRL3kVmoZjuM9VYFCwTGA2c65ky70kiAAoqCl6CGWweIKD
L/J13kWQEArBxD0Fbren/Q/5semRNlP6EJXQvOx1scuU97+A1CIzbuusaQppY3/S/wo8DkF4I5cv
ul8p+6s+G/dtKd3nlu1pgKLOjrLlpZdQgpkB3T5YZMjzq8U86tyu4EEbtuyz7egLTmdB1MH6RgCu
DGLWV+31x8Wy+Yeo4R4O2/rGLi0Qa2nqBKiWg2DfjS/xK2t+kXTFrToV1xpuRLDOgJb/Bx8Zl6rR
6YSKu5eatEHvRWnn6XcGagO/dGxfr9sMgkGYJHL5TeqNw3qtuCQj0rPYy6eLgncJ6emo7YNpotIY
/fDk+zL+HcW5AjWqNL9XDF1IYciSYJS58YRLvJPUNz4zxZipwOkTG8V4LWEo2Pmzoo+5x0EhR8BC
gwMSqzmgVu4ykDTItYQbZkD+JbPXjbrx8uu78RT8qBxO5/yZzheUl1GmdiiCZiCcS58R3m+yjluD
w1SZcnFonLF0g8AnjBKAnNV6pr4EiFyf+KvYi9r6OUn+tsgwOxPesneFCVduquqDnkwuC7eRa44g
9BCjA8zQdEf/920XpqDsh92yMGcP8V8jTfJ3LkY+H/PsiDtHnHLFSQGhin6MLxkDbtqGqRjFKFKC
IWnalQZ+7XkQ/lKPGBQIAc9zaXq4s8vkYElDA5A/OEWZrSr+e+SfBsgUZIkcxig4xvYydC7Mk8qm
nPDk13PRDbT9PXyKuOrExmOnp66AIJYgWuLLUFL/QdIrDfDCxhlQgODrA5EAuNUi80BPoaaGp8gI
3VFjrlBFVgvXsDl0tPkEmkhEGcO1Yd0z+1IgcQMEohufqv/jurYZg8O1LW2L8YlP8TfyUnhmKAjP
W4uUEyQwdgxV9mM8DMOQESPmBC48yrzGc3txAXD7MOiIeEjVgTGxkuzgESPYL/Pmqe/mwEuauuQb
6267y3hyShn0gQznLou36oSzO5vPCUJuq5b7FMs0EXajSRbSOed6aefQ3JCd6QQCxXikWlBpjXub
NA4NOLcCzpwZ2Pw5s+IRpkWZ9zzJDruDXKTEZ+jodt5BpLh9FlZBLZWrGvsLXvSNfK6DC5bVJNq7
kRb2W1DhMTH/ntdw5F1Dc/+FYuL+v5vqYhbAt2+xV9ShP+2/oROMAmq4VMS/GN+ZqzeRAMS+yYZU
UocNBcLDvKY0f01CdBuF7rccbuHHKSWP+HVkSSBdvDF5NYgJ+tJ7p+Qo1kHPNbCrVefGKdyR9dsJ
TYjGRhYIj0rmjyU8SXgwI1Fv71cKShBTyAkGWjNpmJsYjd21F9eKqko+Y3CNelVHrNy73nxbir/+
32+8ew1JulawV29N5oz2UdrTxhXXvWn+RaAvVOrrJi6qsyfDK7eEGjC1FuM6Zz/rrZeXtCI5f05t
EIVv4ysp1KShjwmVngpB4jKxQsTvlGJVMsIkL9fq4DISOG5B+G6/vb7tAxJKns/3WOkfXKxi4YkI
KUNnFQtjOd3kEGkXmLWqve/w28rkHT9XfV46It16amJzpDRDhTMq9QXe5P3zBFYJz20ix2kAtsRD
tl3jxYBZ5ohdJfOzfuA8sc3rq71KbmjBj5k+CD/8mIy4+eC00lYV68ZhybN/udBjqx47MKlds9ER
9TjrVpdP7HLEZN/IuFe5HKm+5qXOGBXFBi4mhXNombEKIh9SfqK2BKnXWenoHiDDS9iZvtkji1qO
+cpcQBO8toSJAJ+drHn/XOwV2pxEEtuRuGnTrdJtvadzpExzBZkL1MwOBwpVuyhYK4zzP5Ly7/Uu
NZhMsObZAYIEYUEdl/6ZSJQ+pzzJOocWNL7bTtipTVvAaIxbfTEjKt3WDG0A0y2VQPvh9ECkfWug
DrFWPqJw++Wcdrve7mDz/OEoZQ49NBMj53a0oKPeUOy4JGjd7pojCb5pkQgVxG3ersV17j84os33
drb7qlHjebFRlfAdyOZ+PzenEh3MQM+UKg0JOzgTw9A0inQKCS0OGTPOOmWJrcalFybAqeXfLvEy
tlLMGoAFnNFHdyE/dddiFo0XMwfzZarax1RqImcorYOTL8GbuJoj+/mt61MOGLyYU4mgZMd9jj+n
cpTLQsRm2n0ntteWZGf/PXzGSylFA1X7k1tNFVo7iVSmmHiCOmkyrABJEydQs2ZvymrvZG/g+0AU
tSHEtrP9bBY9sCi8z6SFSF/IER2MDkygwar4GUJk4W4CVyZ9piw4GVUKor/wD/N245fq1EtgDgKE
pJr0Gz9+e49vV4hsc3KoqHqbelXvmi2d7s7yw0VBP3kKD3bCwmrDJUO9lGhF15Y4ZQATP1Fwbif3
JHGxF5z+qUta0f4xMASFsW1uo/QD4RWYB9FTi45yDswTQXKwpLdjJi9OCI9aMc/xDxwl2ggo98/Z
ezMo90Nfxot1G7dx6u0XIx9hqGb99lX4lUmDyN5FgTAaoCiuRVNUyOeCA3vNMSfaK/+sUBbekF99
CdNL9ZOKV8fWM4PueUTSm+HLQLaA9KEcQo/ZGfe2QCNdohofaoRPeoTA9IHH8LaBVrAifO2+fkJd
chzZH5kV+Z346AcC+ivBHuXf1qv3pWPA6PxdN+hpPmB7X/Ubx4JBYuhHwbtdl/34HEO5bg3iNZnF
mXzuJAEUuR6WiS33WFoDgH6GQv7ikwlo+zc0CjYhtpGEVYVmCgZhW2L6lraX1Y+80J7jYJlYhI9q
ml2HN92bD4eFRREgf0/nIKSmhBK085wHv0lciwx+iJigtkrsygibmnjFFl0Bn04pi2ABXJkEN5QV
Sk02VISmlVhfIkRVzNL32hUAfAqR+k619qsLGZhSddH/SUUVWD6NHaaw00VyK1M5th62PAykqcsJ
enePBmWm8axTD8BUarBcdRA9Nn5MI6LVeunOsDaiARVSFhB1+1t0iKIr3n6ZbV1GD3kKjiWRHUL7
oIhSj8q/NMTyDaIvDXqal4hoT2UCwyZPuJk+TMAQOoVG/Yv9VmFRJ4l+RtU4kGBpwM/+3Adm8UPq
tUaDCjbd3rm5n6F44c02zAQ5LvyZTNF09hAOA0Fn1bBVoU+UlJZ6F5QdLGFd1KPAbJiRyJkGDODT
aZ0QCEWLv0z0G5rrlI0KBL6J0n1iIfb5nDtNoLw5j71e+l/r70jNQVCgP5AhAeMa76vx1Lb/xssq
rG23JukLFw+NpxqXMhsn7vdbGckLgQKRYeHmMlcVbScKfSCIDiGgPTGJbL7DKU7RqpQpvTuXgmG7
YpMIRfMMXLBtUv9Pnmz32t9iWDI48XzwOWeJ10hMuOWcU0XxLcPXJnwwCQmAxSCP0O0R6riCsQxS
0i+gi8cIgVjG3H7H8O9iPQ4rwc/7fCvmpEDjGR+fCYmiNtC8+qpGJPQMqbmJIn+WtLtZPUsPntN6
T/wkg3hYhLv57SkBW5k0DoqpKDglwTGhhCsxFAu/DfUNn7HHor38qMdyEw4xTuMONbnFvBrwz2sr
Va9/PDo6pB3h8NNHGic6BiF6JiG104W2h8rOr1ThTllitnI2so9l+U0sr31B3KJ7chLvjFCaZ5no
g6eyjTmg7WRQT+oRzRR/4n1lfpYuiTWx7+0Q+IEYBA90Ym5wwieNbxeQzv70pymKugWK29xlpx9T
gJCkGgUrkxSMb/r+5zIOXt+jPl3otUQOUeHBJkFsj8lvsSwdP5cAOQH/RRou2chOEF6NVMX3RcJW
vZUTW87XiJuVQmWYQ8OJ7k1T8eDYMzJSLT2vXHsqM7e0jeNE4iUvcDZW9x2srDV+d4Xltiv/+zOA
rd7HFjWSDQGVFW/w0lVJpC2Xx6wOZ0MNdxVKkWpXQ59fRr93rqMXZo+C1/K33omF1FrZsSQpMKQf
dIiNEJYT6ueX0b/Vavy8h68+9e7tmC7yqdljtPSFNUXAk6tKrsISaWArR2I0Jxero/IU3ArSeJ33
yiSxj9bguO9uz9Cm+a/8VgU3r1EQyYNE1Ggmkt22VUAcK6samsH5paj8DSHqmcFfgX3u4CM20Yph
++UcUBkbj0INXS6JtGGXLroYuFW2yyjA0/RgjKQhTdNj6y3qfNBUNS5u5ByhzFjYOjeOM++bQBnP
e2rB5cW3S68Cty4/2uaTAbLe+dslzccxIsaIaNj5eBrGIXnb3AzoYpHr91v6fNo1zHN+6IOjeLQm
ko0mi164JsovNA5yim/tCIJlau//Eh+4U5ahYQS/N1aMUpwYQ1QC0EMNs3NznL0xVfaNcwbL181V
vzL14VBeVmTEFoZD1SxLnpdGf3T/uy/DupWXLEYlNiBIqIDPJiQO7nCa6f/GNUYA8zqOhHf7VLZW
NACgfie1LWGIztNDGbiiggTUN7crNedQGykOzQO3g756Q0xdgPgHPGSsI2J7isuGcjS+zo2ppbHj
HDt9o+HW5T9jAR2YNks99Q2s8QcY3/gGmAohAvHk80fyQzoriEfP4GaHM1iULj7C8tEL2ntnW8CR
M24LzkffYZLnLLdcymjofiYGhwx7Wsuw1uYtlyRMnEQjakF6sUSg1Glfzw9dMpOu4c98qPO/k2hs
NOBefpdXVzDoN+PeonKBzSnlxoU0IKfcd8WgWdoRoBZ8a/3e33ISLCgeU+/q4Zw0uMpnS34HUpkv
3XDxNnOmAIcYYmjkxF/luVYrG8C2g1hQAjn9wKtLTQ08cxpa46hXC2bWVtJ0xWBS2AMPBKJDtO2Z
3z55pkWudk4aT7RkysEeGii3pqpr8EN8RYDnpnPC2GjBPMnF4rzTMUnOcfLA3MSmQnvCy19mqk1s
xclNu+GkTO9MD1c8a9Ar1c4lZky1Aj0t2O1t1F7p/92UYRnZ7Hot8snfiY7JntjTJ5GkKyvDXZIG
c1PiRw2gGEXos60VKiqCXyghh6Rhe69tJkrxXQEYLmFUZZliU+jNzvcUpDnQEcpDyKZWbxVZH4Nt
Ay/0FAloI0JHq0lMNGlSqpVEQ4Umg91CFveQ2tiBx6QnV6XuMTdZL4Xnl3WRI/HuFMbnVElrNNK6
XaXExHXGRIxW92FVHeJv64DbN5a/V36j65kkJu+eUGR9sQAYPb/qlShIluvT94DLiA8zCg/LFcMI
Pbu+Jfk6iss+trZ9UEUkpvIlRuyXp4uSqMcnzNfJ3lfRHNptoh/IG1akVE77RjBQw/l3Mbku6yc0
kNdvgiwU/vl85t95SWg9qfr9IlkTERQeQAw+eLCxiIiq+pQ7MRWuDb+5VhVrC08jczWPkqP13dkN
usMXPOhdJBH+t2LQ0QMCw8UqjdGORw1s2MzSn+Qx/Jre2REUrXJC0URi0THp0o+elpAQkUJLgUSp
teWq22AS9pZVG76EtQHlM1qvfHq/RDJisa4q2UDT0JSOmTSd+H9Dx2Jm8n63O6T3Lbk8o2zQ5HKl
kOKS/Fhqb1R+gK+WcZjVY6Yi+zPQNtCytN0FUcp9co4lWGoIkSOH+H8rP+fBF+FUTPXNebxVBT6K
NRRq3D380jPnjBxf6nEY6yp+T8DfGYeN1MYcBGNb1u2jIq5Ul1QmrvPDEhYDTe1IGWpm+ZBR6qEG
5csZSGC/crKcQ2WBQaRW25iO2u3+DGBPv3iproZg3DdEWIWIxexSAV/Hx5PkkN/ayHKkYjcItY42
6sS5/RexZbvYGl0+q27P0D6nE2dosORE2oUnAnL1V4R7gWtskpgCcaNnUkIiMeFegAt3vlrzavwE
BsP3qjk0+uAFvq+yhALLH2TXOib3v1AdF7IiLJUD2QVFzTRt8uRbLWg+54+j6VYQL0DytzVEho1T
lmKaIj2dC3xwzbWIaQXpI5M5KytbQYyozuR+OmCSQYpcuNyUNAr3ayvmzskuCSXH/vHc2aSozAkF
Sx+bv7nDvolPwM91/lcaj0zGYkH9HVK6kvSZw/a3JuJ/vFRS2t4WffBMcaWqK3IbBuNLfsc51bZs
n5l8P3Ri3M7FzWRPOl5cvj/JWS6Hxb95SnWJv/92nt0hDm8JdxbM96M+VnQ5APfE+CGAM/b1ezoR
6o5vmCz7vXeN/CwGLr+QL5E3WfgyvQd+Sg4t+sRL5RfHJksktITD5bL2J7UZLcpFahpzyIzuUZyr
Qj1SZ8DBjy6wIEUHWrMK7/6T/LbIJe/LCID1vID0slg9uJD3xX+Xb06CrJLLHCWtTN+7/WY/AHwW
GGJfoGkSVs2EtGXuJGWdbQNPmtbYAOmTvhtixUnKIlagckc5auEBlKAPqZXVGRD5fDVne2U3S11Y
s2RV9B5rX/jxJT8ehNkEftCRfuqp14445k+z+PqG3W/BkLbr8NU6tH+uzidML3L3Z9XInvbR8b9B
b85IrkoQ4NoVZCOzriE08O2LSH+tEXDdr7FUvIjH/id+PwpCaaNrsFF85whM0xNqqO+GtT8VCFHd
g/WbhrZl9VY3WdylJxrUL4QrKe8Zije7e8xeCg1+kTS3W3s2xMH0/5rnx0B/iXFHH41ouLHkTEJJ
3+U3yccYrKv1PBWuhrEvyrq3o1H5Hxey1xNw82oZ07XKRQ6vnoQi0RtgjVxNCuLhD73ryunLY9G+
cHAuAnXC2GJwuGiUzfQgaaM7k1hC5yYvnSmq1KT3LJkTcb9etyWHZduJ56z6AixIYr9i1aC/2nv+
CMOr6zeGTwnKQJ7d7jzAuRSGNf8lJH2zfnSKvXKQmcg4dyyAxBiqNFnGsodn6+eS9IeFcD2nz85s
nuNhnzSNLEPHUFligbQXQadOQ6/bcU/Swd1UzlMg227nLFlYtKq4FRGactsUxaPaxaOQr/OKtmI6
EBi8/xvU1DhMBRm90vwhX3AaCCL5uaA+aiUe/FoBUnmMPVSUdKIHRfJpNI01DLgZfZPm+eRRB088
17PrpqFiY16HsONTqHdWc9sI+/1S4DMtHRal4yC9Fwqsvx6DBMUqGF5tS5rMj1fYB0ObGgVxhyPQ
8IdLgdkrWEHX/+S5hEvkvT3UF9x2YGn3RcOHACGGY2xeAzqffGKvIorSKo1sNe70zAcorxMnjf2B
qzrUpBUq6V0XOPBISTSAhIk4bLJ2ZIyUWYr4za8h5cHOp5DI2CX3YIQVYjg3WqlH9HaopV6ldG9J
g3Kt3m+RkTDKfQl787g1/sI1F9Sn6F4cwkbHWMHbP/W011eMFaObYzXHjOQNNDY/+ftY+f2782AT
N55bvZg3lRnYJbuYRj1Lh1HfriNj5/aAnnZHV35YW0KoauRj+4mAKtYsqqUQwAIe/OEccs78bRii
YtwVwLbeqFtKxLGk0wkeOsHhO0rVdE3HDdjFDmf13RbQZt1p1pQL3seMeMzpljnEBKyka+etEkh2
GlS9MoQQT54pfpPq7tF21ZftR26KUFgS7s97gBqH/yH6JLOpgIHiHwSRZe2PDv7gM0kiZfSLMPAO
kfcH6MQ8G/QibriAD7ETsMEOY+qVrisSCUlPRhrOEw6r+321CpdDJeSiO9gj8v/M9XB6Uv+CVCpq
P7T1leWdjg+qLaepArV/bIDU6VShwK1R6hOazSw/ctAC4sCGLUVFaDwodSV6YVWRK9mneXi4Zp8B
HRqRBz0vrlY2leuWdEXCilwZmsovlr8jnFD1ix1T7i+OZ1v5SCv+wwwWCtN1idY7ASRW5k2lWFAf
ka1uJvqzU3W7BS1xWwZCcDYn4m4LlXGWQkg+VEPT7m6nYv1TSZHGCRJhbTzAAvLZrhN5AivUi1Zb
MAOpKxE8jaKqX84uOAAlOKLfn5vCkeS97QEKwU94tm5EJvUfObTbFaPErYztHGXNmMtqt34+NRk2
+bevcLoCpdAAX4tvk/LWgaNgs7eQqghT+XdmbzRQSDv67iYryKwbgRpkikkxsq+5lYdxo8DcSjR2
CYoyA5kYqF+PMtSsjghXTcn92NAY9O1uhvnX+MCyBYx8muEzXXUYf0EfuX2QRLQmb5AAvr1PQtuE
3gAbfVxC3xwhKSrk5gIWd5E5/Uk88R47VMLjcTrSpoqT5VKU2p77ABRtFDU9hTIcQuKdzOKUf5xJ
CEoNTYTjc0pO1ir2lr7gWFSLcdzRBuQV6GM2sPLKsV29J6LZDVCQcQgBOT6GQzTh1Qp2h9AQv7/8
BV2vntIlAvZhzocASsMS1XIzxwfo2DSK2gaTmp+QZ1yrQBSvnpV74mPaLJ36MYF7kF0dq4qofDE6
kdvpUwop7RmrWNQjYjCwIKyUTA8a9uIQREmpl8BQ4tkHd+wf1Z23lX5o2r6hvOWU3H70LIZSfz/G
bodGBoZlbhU94yay3Uv+SGlpDiFVoTPGaGyka7b30q90siDLYpu7K5NdsA130qW5mLc+UWpH5fAu
bPhuhcSkGUOZ1U/K/9cSKLyTd1s9RVLyd/9o/qlBed5kc0iLUFuwnN/aine/1Ydach8qooN5tIx1
3Le1sizIP2pAfHH8oOx+ysaNQKy5gNCVOJTp7cESAMkfF4s7Q9czvjVIecWnQNl3cENXi9Sk+oMh
foAUvTaeBBpl9CQTkDQIuykAlPWDQA/v8Vwgh6oAttjdPUQpwpDmYJOpVrehSMZadgKBrBPEskYU
ggXbaBtJ7KMWdH/rQTDaOLLhOyXD0FgXXs8tafUjx3ZVZ1vuDHJqWoVVGNDfLAGaRUCENqYUUdbA
UN/6WcvWKM6Q3n8O8ifvW8QPiEpPS5ejhKM6/El8/sOBjXJbCiA8AOa1FIIyy9acMlAsNvR7bCmv
UnXM9bvIaTcYHSnIUiAB+W/AsQuiCLQ3Z/w4z7njwouSAMLQUhJwIVWODcd8peDgLDgESOEWPc9N
ma16Sc+IIyCtPzkzQPARPvEim/Qb4bJcY/MwPckbgECZJHX3+I3TYwWHM84+PG8m/EVSy/bP0WSd
O77A+ufXWCvkY9q57CsPZh49xcLkNwOn+cN2IYlilb1uHZmw8/E+p8Pm2xFdWO7T+d/sOMiIwfHE
EhEN7wzoD69JD5vbWoI/RHNvkdd7vgaVyP8UGvWLQlSJ0HxF7ll36Xu2l+wlMtBexun/v0iquOIE
NDANBa7jmnZDP9N0KTPlQO5yz0b99huiXS7X58pWdA7GqpGP8bPCqEKDUydPKhXNF8/mbi4aFOwF
UkHjXWtymtVhcWTk4Ku1/fQTVHd47j9FrcWh+CBGC4oriapItXGYnd8oEgH022YUUfh2fyuwkIlq
38wA0FTNL4u/oR+P9zD3wFBX62BfG+AzERn+yqG+URzAxe27gLrQJ42eCnXlF9o9gHHjyPA0ibqN
8y0Q1ABBNV7PwOU/yM1rY59Wby6TAyb0diXPlWvXJsQ4+7kYDGAaq2jRbB+4i5zNzTk6tG2Zmldk
mZB5irJUjdtMp79ypMtDcq8zJEq2NjWawTahU1UBgvFSx4nNIM1Jk++oVjN04VLhqO133++jtrlA
srDx5RxCO/45j/fL8sbyce28mYEHiwljjeeATLEHtPFOiKEJ31edEO01MDphgDwRodEXJBKpZhMz
dqBNLyGt4kbpIo7upy3uM2dME9FddVBoLJElCzKje274ZqaaXi6NvGk4jdDPgjtVR3QVRIU18nIh
fXZ0AoKExCEF72OWhhfe6INC5eY4KWLuHIbA7eAlSlzRdFytVhgh1r1f+f0C9gzdV56ra/Z1IWMu
rH37iASIwHhbYTOBO+56vS8FMh5j/O/3VOlxkBDs1cLmfn62s2m5WpHWkj/10LnNQXOXqywk2DOm
OWDSCScuuz3gXpu0b9jmtIXbO0U4f5fk7AGoE/q680JpeMR/z6GgQjxzEHtyrlwrRkP7RZGqsLLN
xeOAjbrh6ok1fxeyhx8+maoCwHmRnIdE8yqkssvgf6od1F1NLGDmMzVodBLzszEcsrt98dScR+Ez
cBygzx0uDeeku73plHfzH7qXyzAwwB9fWgxY5IMf0waxq7ZJ7HULX35jz95Y4PydoBAmqKnPSd+I
8qYKU3iEs1nSETsFpnIlnPrBduomfO+jLwKZ+MQ/AdZegFZjypclBJrR6XEwD+4E+VCw7iDWjRnc
/UWX27cBULkHo3Yi3zvCX/VYOiz2DWeXtOGza8sVUJHn6IRUt2wRcUIPZW+hit1Zbkj4mbuEjobn
AF63Vu973/0LyGThJZ3IxWmuhJHA9QDRazs+MVKsGWMmgcd3Q0SqjVM725vMqKS1P1G9CUlrv7GF
DXhyK1K37/fIwU/2rhBw/vmxp69DHl8xsrBk0P1/wUzVMzfKHKCTZRtPwp3CppbaiM/HjJeTGTg3
erfx9oNW2sWlK1RA8xPCd/WeqQiiVAIJ1oZSwMNM6lLXfiyFGm4sWotmOKpygAotW12+4niDdZOt
T+eyzHHzKn8OF+arm1z+KQDGV+IjgphsGot84S2oAkSwpozoCvzKqOJuqS/dQxu+t1r4GHk5Rw+L
J5Ow+s7rmhIUppmR+kKhV9y/o8SaYDR4d132sM/X/6MJujiIHKwlWBaK8obR7jb8GixtonGNbWrc
NQwhOZawgwCAwwXkG9aT2Auu1JFvP7CWZTkb0eDxTNLPh7sLv6wsKm1jCHhncupdZlSOzWjHYmXM
Q8pPs6d1L94cAMkeKA+cT/i0Oo1r9WuPuSP7CY4hdDi3ovQxKdpoTeV6ygUrdXuMPO7xHZBw8x4/
ugWjopZRbuq9Lc1rOPeIBpqEsIbb1Ze6I/qzu3v6u/p5f02QXhATfJcB4LbRuzOqkWlJBvixCLak
bJKZKYWEike6kbPq5mc5SnXY1hc+G91LF2g8NjYGKUSYHXLqmuIlnvtUefZ7ZjFLa63t/KnJkq/9
YSKaRpKqES+K1wMN+h6whGh1NLzpaxdso2FcXKtgA/D7xyNcH8+aBAWe7cJsQMXO9fkyoB8eU3fy
qV9Rx30ztcxZJMCZJTo+mBQAwSXW+SH18F7TaBdGx80dMZ/Anu3G6BT4xezj91bEYCZqAPbehfPI
ybWAP9tNi9nwjvYy5651yAZmIlh+WLUfQKyenaDIz1YS0V9YYYSVl1Sv/D/dH03MpCcveSnFwUh9
jEZY2hbXWZ+dIz+rhdofhO3nsLfjT9GI+1LMICRekBiR6BihpG6YBbaEQRFfKZ7h6SPTHEkWX/KW
1TaNa1CEgIJKnCnsruY6GWfBo1Z1WIecUmfXjdSW6/bfSi1YygjD6IZGYFIMqHoT8etTkNYhL7yq
05EAxJEefkX4l8nowMdSd4wyZiN7EsGKvnPvMD4vTxHm9yUcs1+Wx3XY0gviOAMRPnOVs2T1LYY0
KRgS9TkNL7N9yjhGCWvpGZBo/8THtA8Y1/0nL7wYUx4Fn8gZHOlESwfT2N1zZXEWM4+UIYlsCmBb
B6zbXXsgflpDVOv/C/fG7RXnzDcyT3/U+jB9+b/5L0uKigxSSZqTGURNTIs20Gwp+zjKhfM9jnOA
Yk0O3x/CT1UBg/AWYPtnJXTlnwT30XA8l8O8Yu7tkFd4cpGQ4jyJGAot3g2rxuFIGFNB9nmDukxw
l+NNrdwoTq5rkKndQFcdnuk7AUVqQ3Ea9Qp1SetS7XySHjxK8eGzrv5dwCwxjL4VHunaqs0d9hNH
leo1aJ2qudqHwQC2jdrcZaOi5L4zUL5GdJUgOjLvmTNo5LQhhXErzHK+sIL2nUsjHDcc/WvANVmE
QwRBLKtgRloUNk3E8D1uUIKUW+gkrHI/HtvBlcwECQ8pRNzlpV2bY1jApMkHfq1uYg6ko0ZVsxlL
DzfeQsIjtcdusNrqmOpr+FVeaS0TfcKiLF9XeBBcCATCDSbIweMgROZHGyuptUAYSEGuvqJRbGkg
7kA+xbEVUj6uvmGAR9m8gFZ7GM0N7h920fySCLi3WncHHcouI7fbVqlckt5zyc8i8hNYynrwVA76
slgzKGKfgXKfonLgBaQDHca4Lq4SKPOp+Mwo7ix5eDORFS95gaYFDAmLAD91J64it57k20g/OLDn
tfJg6RSC2+wC7l47yNpnG7mYsHCYAF1yJmTTWg6VBexYYfCIYlxnA/bKlr5hbcpmrCK7L/4I8JSM
fOP4lp29806xkSOhUuCrvNmNpuCKHw7RWgMGofGrlTa4/+EzRvYHcm+z2825T3KdTNiKJM0H7ShB
nB1sMvMCwLDMxQbw6hVeNbNCt30J1ps7w5NbDTH+TxbKmcbPScyHk7hMuLBW8a0iJ9Zm54sHmucM
gPp43UNokEXqzYBc+NAaZo5S53uwzfOJuODtsi+8/aulYDf2MCdhykIA+cLV2K56FRtPd21il7C0
sJxgSqRbohvJrzKk91cLut4p6mUgj2u11G4+4UVlHGZGq2ESIwvxoUoYY5B1xRDEO2UPMyqeJ1Cg
v5raIT7lHMY7qGDzKZUgyvvdNBWlUm8FAM+j/eZDa2KAPC4TCJCAilZn0kcUhxjSW291rxP9rEXT
me6y+gwFUfOnR7a5QGS8Q95YYO0WZRwxXS6ELgzpNurm9dQmvM956UdigqEEFGYc9XxWNKtAF98s
uLCseTMUkt7agcXSwErCOktF2rfxKb42JiMFDI/x0lDQzWjW1WHPuC45CWoyA+CssI5jbuIS0NsM
Amre1mN46aN0XVMy7GdWO8QFx+NY7mU5t0XcISgbLlTHeuhSSV3CoVKLLypGLM7qb7sHtjACjliB
piszM9b209O/aw33W0PHZU3cbVH2gyMKYTKVjbsKE9E5To1ZfgpLxqlj3WKg+msdapl0/dvhy7QY
YIr58/6qlYAJcR87itDpulkGWutalB03lJ1uM3bxhrte+qzChwVX0w6ZLsawZJ8FkcaYyFYFyhPo
9BTWxh06YXTlYYhSpYs3u+wThkl7pCGPYCTJ6Kb+Rs0ZEULM+K5oaBYRZIAXB3VNULlcwuxNzOKc
c4u0C5vA9Zx+N7uBKeO1Z7+5nlbCtatzjE+WiKrcveeeaNH/98c9geIyBDKP0j6nkxO9tZ0cOQdq
MOewW8OEcXeNIFRNbFCIkplXCUg48npwQ8dal3mzDdiOBOo04ld1QTIilp2zUOWzfvQIBC637wIG
52XcLET3qOs5HRVCPp5h/q/MIdObM6Y5J36ToNqE6YA/s8XFlu0QkR/EFsFzlP8G1i7Up7KfPlua
t83oICmt8TQUS3Fo/HJcD4XmwMGYB1xJJOg0jgZVm8gY/16jmiPTYVePPV3r4qUF/Ja2mkGzcwKu
Dug4NwgD+LLvMQsMyYHDlRDx2az0GkdW0HF/VNgpkdtc/Dl///bEgvuLGHP0DLygeDik0aYLmYMZ
B6WdjbUDYtrYvQHMI2PRP2pSEh9P69w3ZSZIiW7TFeC5zTvWbTd9RzlNcuH8zGo99G60wSDjBrxr
cqDcAwAIsVUneuSwiXWLPl4/wuENDNSkTKJyDlS5Phul+LTC9s+gXxsC4Rn02MBZpc1ZsY7ETW+E
JRjSvRGDFQSyctLknXcJJZExY/kE9LBwYDAKHOT/phY+WMLkejDPF2PHi9kktqOGDYHqJz5Dn2rs
IE3kfWE75JVcBYarpaS++e6Ag2giwqjvTL4YHVmss8pT3gPEvG30JdVnzdqqYmYDZP3nHJXSctk3
GAajfNxJnAwpU/tM6WPx23celsaknrTUDFfmQtq6okepjTfDHx+z1DEZhOkWr6p1qOQBIurX205i
wulJb+pHpHCDFDIls7kXsUXbiRHEWKN13QoMKjQMCtOp6h1+ilitzJdTPXzHK9H1OzqEHfbkcC6Q
qYF4p41b3+tXrrwx4sNZDSRVfRJVSeGbtZTae5t1CogiqXeWqdHdhwv6PzXWOv7OWs8gK1YDNjTP
5wDGX7bt8NrXai5i1MjhBaxvG7IHETB00UBwjYP/fh5rxg1x9mAq2/5ii9XNIelAYzHIVxL0PByF
HTolshbk1P2MMR2heRCy+eJ3q7r7fodRnU9F4IXdLxoRiXs/E+2ISXHoOi4+WD7rFv+AybQ66CWz
GNgf4IPmyRIQiyl3Je/iHexnun8psZp9HYIbtW+lizF6uAAyIyfydhPOV1iTQv5cCwzLPLue1Y93
NAuqQuBgE9nBdGk+10DRdNFARFa46py0LvJw0CHl1IksvkR3HMqurYw7bplSBI4arLMQveg3UYUd
ynFa6hV9iQ6iOb7pX3FkUk29q9k9/k2J9oycjfpw63zIUFrM18OSgdjhWSK+6nQhlEYxSVWMxBbH
xfqnGjc8TYBN6snO6S+clCncOJ/l02B6O21PqoE6mPqIepXViDhKIFUbgVHQW9MRcv27tCfRBgUa
OSb/F8/gptldNsOLor1fj7KelhDNSsGYtqSO5KXq3Stb37HslzSoAQVRcrWHmsNIPrHdZ7byFcpa
9Zj3ODK9NeJ1ysMo3hMNhwk0w3NNYefuJ9BN2NaZCnzhiZFmxUvuolRXfgF3fuSOpO+fi4kxyuFJ
GWChIxpS4h2o5r1sgvt+Ul3OX80wsdRkRKzv1l8ClUUtpktazaLExesONWUo4bRRC/IyYDDdnD71
UlreSjUcYLc4k/B9F87e3BQf6foTGNCPNraamiTWSSXPczG1GF3UovNrC+UDRLwdne2iIcKfWyLz
rYavG8TKr43z8PWLoGu1tnn6urpdsr52GF0Mnp6uHoPLUEqwBeCHWMr0kIAonHmvUXi07jPRKnca
/UhqOdRVvGOk8oLz4Azzjivx1PSLr6TkSVip6xdv/DtOegL2vFTJANOj8Mx9TUEAKA4WI3o9/eeH
q0JC4PvJEvgW3GF8+gfsFNn/vs8EWVWpeiXxYnpV68OYAyDZN2Tx7Va4Jfq6lNsH6DUtm/o4VzO8
PV/cM5Z7BdXQMpU+WMMk635/HykLgvbr8aTBFLzoxxOYi1VvuXDD7LhaO4Hku2GPO38AR3Kz9DvH
qJDd+NL+M5G6TP87FFsVl4TLFnoGb/SGL7555zEysoOZgZgZ0K/mno6XAUMJnhETc0Ar9pml5gpx
OVLehilQyaxnOy6+5fzz25Aw4ds/7BvA6sXS+UHUfr6uAHOiIIJGWN4bqC1ddyKjVcy/zT4DLAsN
ZQ2DbyXmSUrCNpSmt7QcZUlKpgl/7sq81YZmGRtIAlj0S/k+m79dPMCxUdA9BRhx9vCuKbMddF4b
Iry4u4OEeee7KtAk7SDkwesQz1aaFr+1xOadWswwvQJymC8wk72cFCU5fm+8xL5Qf98lfUFBOAIA
wTePIzUWjraJFwoArNU9wRuOM0uBz84UPMVaglWg3gEDHiQFBGGa9vlCqEp8vkJfQMeThoJvB49s
uAXqm5oA0hdWRRCT1gd8SiPLzmkqcy0pehgv11q2Cqqn5hDYdHQVz9ZuRPM1Pd2lrlBqI9BM7z99
DJ+isU7BJasOhL0bnIo1e7oJ4qH+NmBBsipvWJct1FElgkwVXLhB0QItjZwrllB7+fOEKhGe2Jnd
G5Spldw3fcSzsZz8rV65PgejuozyHZY9XM3cBVNph9t9tc3ttdt0Jdl2vwUQ54OdFuSpG/0EFBhh
cwWYos+OcQSzCLTFYAVtz7EGUEnkf1hZlzOIaXMSows8Wh3lmWTGGxntslewH/rGnKDb3JhwHaVf
MLNRrX8UVtrzx0y5Ys2Fd6eOL1jSqrrh0fl0UwGjXhUp3UCC3YfzjYYxI+HVGbnlyyzN+doLaKhj
39rZlxO2ZiG7XXgWOtwwIZJmDfzUjQHNfSQijzING/BZrzwAxBLP/1NFWkPIiLvrSjtY20KJoreN
fpH7xdQFlqH3WvB4MuW6/aR+X+A5C93eDG1ZuylvuFTclcvzz0YTaXbya/scHze3nS/lwsHHZyIz
rea7566Evtt+28iRV1n29OMk80o043UCaAWpATsFKwTehV+DwumNmUiu8wISaRDmBrs1XczQoHrc
KOUHFVQWkdIQinhcUVgL4DGUSegNo4fYm+n5BTS6k3ypgZ3/LFpQukPei2XqnbFBRk3HgWqV4UVj
q+P5fZ+TInFMQKcCJgjbtlZsbRZ20wTjnnDDOdxLZUic9evaavH2wHSSKDZ5G3154bW+0VNcHDmQ
TlBoLepLAECzCs4EfCTyx2ptlx13Qwow/VIixtISCktOeE03iAuV+9h2YMMjJMdcknpBRw0uge3V
0B9P8hToL51ie6+88PWcYygSM0iaSVaEdikqDKkR4PA/sMg15LKgpOhqv+VGldoPGsWS87unrG+r
VPaZhC1/PlmRhMeP/AmC+qKoqXzDQZj66PCDZx1mUoPFRfhdy8CvmEYiv9jtVgWOWc0xFn0ajO1G
89SbVpJSJXbvi5j0NVnNjMPJ3oL5qtPkmew49gmYJjVImaN2pEntvD8Jve1PI+cwVU1R01V35BhY
dXOWqHhKJbb2mVuNDnS+262kq8byYnvFWBzbnAPYbXrrdPCNiCtgvhkfHChFGsns00sO3Vh7ERC2
DvHEPg1tisCpdkbxF+zc5aRuGnWDAKWu0aVfQMUDisr7iv6Fn83nWfbWEpxm6VXc1CYpGjwyyCff
QM13w4W4/EkWfeJfl6ryVpA5mcAwcNr2kCBH8g3t95yRLWrqpEpXpnGUaPXUED/KMHnoYTbpD1He
3OdPfzFnn7YTYpnvhbe7QdB1ZhgUDN0Sp5grTL8k1bZdu7dclYwCMIaezdcpNBAO8KY7ZhhGsY5V
y9AI2S6a1eFNuqXFOQcttphxDuxznhwLEccHVi6gmO2PuhxHoHhqg13tOuuMvymX0s7C9pdzovCr
onWvtuKkLN+O2C3K2Dt0K8t2O/CY1giRdMlM0DY6hfY3BTCSXzfEfmn4+Y4mhbAiYohjwDmc+8f0
CSGlJgF8r4qcljLzW4mcK4JBuhC3OYkRECNHKWJB68vdYvbRhzB7+k5gu0sMhLeFYFhYPxlUEIKm
eQafTLyT/ZFYvb2nF7GNP6u3kLdJzij+AYdqJs95aFKRs5ecDKFZidMG9ilM3GXDXiBGjUTcMJ7t
Of1oz8iMDfOUI/QnDbbSr9k9mYIMV699tng1h1LyVDyDpY/RMfE81VHn8ZEg2ICk2llRTxKZAVGL
wJJpXf3fkEfvun6L02+FH7YGywa4JqPRJ/iIJrma2g4LNDeH0Lu+llCvP1pV7S9QJH2DCFuOOv9+
lBIU78TCl9sZHrvAfYFrg0r4JTpr9C7fNwrtKgoGVgjanrxliF97v94bZwy6oWcvv5LUHSysoJ1k
e/x1N7TmFq2aFp6cmXUbK4M715fdvvtYdo1LJVhCNegROG9MkXhhTb+lPL0PzE7a4272XPNmEk/A
rrLpV9WQbz36BFjtEfUb4pBb8K6FBNZ5doGuwsq3ex1zvYUpCcyFKerWMXE1peVB9xGYI1pO9hjE
RzsqxvETyixjoq9cpA+U375rRRyLiqPF17Md5flvWIvHkgE9zJBqVwE8t6W4qpS8OjDp6pyHvprP
GkLBun8iWqfvgQHvtBtVme6seH7JxoT0XCVkvrFvEw2ZnYmOyCI4mhib+CbD1L/Ljr6sIjFdu622
ttJ4SuoOwflIkobnHPmLlf1h3mi04PmhUqj0WY+OFgRH5uAnpbP3aoqHj7mASkXHxcgc2PyRa76I
IuAwQqy+YpyYZE5tbArsbkoT07l5IHEdRd/VQZM/+Jmhnn5f0lt9wVOJX/+KL2hGQ1zRlLr4zTqP
IzTaDD0DiteEAl2gq5VkBd1ArTPCuhSLlQ1441HG6Wj/F2jJ8VeHyRPqkTjudu/XaUXYGpxrUU4x
RVnLC1/KejT4jz41bfpPO78gQZlMZHjASt3azmi1RicGwRh5kvqjNnCK+18QDQt23Vo7vMPiP09X
P7ZHsYyDi7P98k01yHeurG8NuDu4JN+feiVWz6dDirz+iiVcXbsVJhmgeMrkc7hby3j0C1ETATXa
xyUdNjryvPGu3ATBRz1853FVw7ZeYz+ZDowoXp0LIgvpz7UJzAET3jGQyvxb4clFSwx9cRTqgX5G
7bDDe1vWEnzYWVkHbaR52Il6byxOOsDc/ol6ug6JKkaBrD2MlGhHVWdFaRiJp2WVPOalJzA70Tte
nK3dt6EOCkpvyt6/khcP78pnYj0yuFDBvgTmsZF+/tfKHHI6fI9U+DXEJz54klhHmuW8MV0mAahf
F+cw2pOD4BBViOdlJiR8Cf+JrzSv+vFHiTrOX1KoSZFA9W3iJcMreK220ECEI6QdkNyabQuDdwDT
TZcxFdJHTtz+nRol/urMvBG+LBaSv4X+Zt/PVksqsNEfyhnCURpkKt/VvDfhhUNzzHfVPHtGlvXt
s0Q3pEqZPSkvDsjWOLskDLolyVXUNeCavl1vxdAb4jB6joaEcXvHupvvWI2N6pqnOsb7+l91dSen
oT7CBwGzOisVOrGbpP7V9tak+nJcfjG6XIF/L/rk8LJw448dKlQBCpG0yIUKdOiKORdjXaeCqvWX
aVW07ZlOqjMTIMR92FASaH2FLy1VIPhzVGwE43/LYshofzTzbuKhhEuIh+VeTd9NQDXfZIm5X67j
bbp4TMmnap2s2O9kl2Ap0UGH63zDqpC/k03y2PcVUtDlztG8m6gquTVrNihhsT7qrIP/5/NsllWW
4woC7ENCm8HCq9ToYEMaODZP+elSTE4VqpZkzoLAXL5F3ZrpADBT20OR4hIbhDH5v+YrHu7u5/KS
DMbJPlxKU7IbKEn3HSoprFKBUBcbcFQ0bwR9dt0FGRHK/tHtQIuSF+cx0+O9S2U6iyKZyx8ynkKE
U8DAApj5I7scOfWntbdTsUFEqI1YfIHF97XxOgrNxzvT2qyRBC6BND3BqtKNPcpHx/kZthCX68Kz
XTkr7Des+F2VlwyfrDpgP+EfbYcT75SDe6A3FKTR2AV74LUTnL0FjjkX9oNIc3ZVPltU9C4qgvyx
zTmp6R2UXGI5dKLBgx8juuWUSfStJI5RjIhINCEDc0b0cSZ+LYLURTff6EpWi9jMyp/6TK73gAeO
wyw0qWRa2wUFMsiqPQ40FxPXrEfRBwY3OtlW8Rx2fHj/N8eNhMVDTIiJhfPkYpsTWdAJJ1Bqc2zw
SuqqMcW25XHYuR3DhZRvcSunyKyLYyxmcXRa0ghmWHWN/+RPXiJI+WWIe/57UJdCM79dYQBzG6zN
ZZikWLGrMBAq9yGqic+XCBt5h/EgnrMbPeAE9jcDiHAsuCXqvob8ahafjY/3vmqvdP9oORK7ZSLZ
fdfOb6quMdaftW6qCa567QpakuUqMmWSs79g5qtfLF0LMeYGuUhO7Vt82CEhPWMsjGJisqKxmgeq
En7kd9UTclLgTqee+iXxHGUbwF0Q01yHmc9Rc6nlbW9wjhZcV1lfPf1UlG8gA1GTtpBFzvD0/EtG
4lpNflJEMpDzCkfrGMv0i+dbhvI93litCd2aS1gL98oBOXo8ytGhVFAeAnXkqj9Fsso2LjXQkKGj
jCH5dOCwic+8DieDWjz19wUZ3MDDJ1yWd3qkdoeZpFes9+wMYVaBAxKmKD36qlDgS2aY55GGQTg9
ShPlEfDfjr1ENK7jb4t+RVtkxxmtcMPI1IwkhkrEqRkVwphkCaHpNY+p9lywjoU48eRGtU5xKmJW
d7nzbY3SdBu+8tKfPmIbawIHLQxhvcpTdyDET3pKsOHEXaivP6ADAolZABAxDH6eSuR/4aoDOoua
WH01nzfkPF3qijpFet6DbZrAbZ4yKhzMQe0gUorUUPLCuYeIoF3PaS/NMkFZ2UvN3vW8ygIeer/d
ddy/FjNDH/zDXEEOhF+h3wb/6YA+B7fgmNLHWoKo6LeqhMz6v7Kt8pop5Vfx8u/GKY8cS3/APMrN
mRfwWqzisD4PTrxAMR0kyi2gJR46H/ZEx+U+75ASI7VZM1I7bhqAhECLhxps4MLHAWKmdqcCG4pT
6/c9YoggIj/4Qcb4+3YmVldde6zggJBhunOZKDRhBWmMRBjLUpMnEaHuV3lEyVz967WL0dfgXLlb
7nf4CyF1RddI8Wq/XONekCrNl1w5Z4owiu+FS8sCl/RapLHGC9RiNC/QG+DCwKBzGYOhfk6zs9p5
bZ6sByTpJb1areYixQ6SrdfkKR/iaA3zKXzPijMKfnzHpVt9KE06tqbQ82RqAg4HqDqT4dLyy5Ih
7d/n3o+ZY70kFvmb9/KU5tCSclpEMGD7yet5DWBWL+gvu5kC1fwjfID+FAIUn2Zw5qykrX7kg+Wz
rCqGZ8ExXF13y48Sh7OJdpoggIXKFSc7dFwX0mMe92/UURPLC8ww22BQnyxFwdzOnzXG/PqkFGl/
GhgqqKZqCKb2OTp5fVUqJnRgA1aCqqkKLG5+wbh+92YaC9wKpxLBOS1d7eQLroEscf2FHOIlUHxa
ljZHDdygSkqj+e0Nt7ht4EJrCyC+qhr18pHgJyBT8uTwpb4xKXsMMN3wlBZll0NYu090zmQ3K8Dr
RroEhmUj9COHOu8UReNEFeNdBZRWF/n1LtYUB/pHkm1C7aPC/kxXbpApQ9wZIRJT/l9/LFXRLyZp
QPs5SmdVS4rcPq305ilTJ4W8fTiD7km72BXgYHhIuXIH8Vu5d5TUQaxBUtXQ4BwU16WBbCGJIKCR
L/KxZy2YvMuyKlpLiRMIibq+GsYYWnf1l3UQnHW4zERmkLD7FyPgkL5j7xObML2fzfPCPa9bnvJA
Mrx1+IDzk0vkwDu1NwX2sQtDAj4OH7rXMdfx66ErGZ5iAm0CdctKE9ehkyVOTBlEnBqFF/Z6Wzda
FM0PmIoncJjoph7gCnHAB3APcyddbmSQtQa0iQpetDEONymc7+/U12SXlTsfltBoygrxPurfr1vj
Nf9li4bty8tzhjbe7eQGjHXC7rXHE0FEFPuKXm1ehGP4sKBqvXxhoZOxZc3a2Dwv7Xel5ZplwpBh
HvEjRdcL2Mv3vit5rc7pJgaOZL/Az66f52CAvU7FwDCh/rtkXUjCYWHoMdmzrl/VX9fzmn6myZNw
PcQxPb5gonc1M8BesKdNOo2j+1YjPT3wGN25izTTYBQ5gGbvqBk2pTVP5oNrm+drA+lrHRZ77Ln1
JdoWDh7ABP9V83y+LIQFzjdS6vuQsKicPqMa2Ds2oSqqzaU+y1oedyGXbGJZoIhV8JLpvpiqg9yB
7m5CGOYEe+1Uvf2YHPsv/MqiznX4DYDJoEc8avssWXH7xahYnnzyXFDCTgDc7Ru2a3RoAb1MBjyF
S8aE+EQyQybfvliQU9X7ZCkiKx/pr/qeZ0hXF31vhzfyDiCdFyMJAS2iRwvdqeyUV6+NTqvIuyb8
kdW3OQcKhyuODt7UNFvSQ4mPOG5z4tUKle/y+OlmO2N0ugjm4I8F65kPZRu/rtOkk4MiFNYbnEc5
Z3JS8C0ry/2oCSmTDTHi99/LOuNmY6b9XJAISd/57jeGT8qCD0iniiIp+ba6LtLYyW6YrbBEJV+l
Qa/vGE+aKKXPzLk+7cJYzI/Lzaq2LgsH4URaY6O3iuivef7Bq7WRUIKWyiaENlecQGVNQNrQmvQa
Jy9sJpGRqICnZfF+Bgot9zC94eFHbG9NByuteAZ2oZJJ01YKyqNQ6tt5WRBURCS1aQU6VhEm+Me1
vwPwURjqGzEaGF8q4yERfSasUbYqYl1yorFedD05eF6x2v8qhPhBmAXGbEBlXQZKBG5wUW/sBZGA
c8QgAw8gSanndHSjYAQP7YITJaFNpVSWIO2SDlbSEJrVFUanMMtf6lOnLsXUxlHvFQQKX7P2slzm
Yy2F0ZpBt10rxMhQTeC8peyyf79Vzn8gFM9UQyp77szDIoQbkuRgJ5a0C034mwOmViW78t/sQfdW
VjE1+/+v0YvjAUHlmI51817RxlKdwRuNr1soSwpuMwByLcYII7yW1U3RKACits4TXrJyGUB9Ql+r
2tmRNl87ezcVt9YZvpGWJR38at+0BtOikP2ooNN9SPXYqZg8+umTMWjamfWcfQ40rKDbQc+6Qh3i
E3XQaQ0OVHfAaBEsGTjcAUHjJ1UKUCcwMWaFV/LUqXVZ7Ja+RkwRY4YIC3VcmLy+Hpc2rOUm2MSK
YZDvJalwMvMth6/fP6Q3Wbwzb9HpN1pW+ZMcM0jPER9+g6OGxYrByVPKQ5aFy2KrepUERvryMfc9
WQBCk2eBbWxMR5TzD9G0SPbaG/oLshiMho7E01G5xFZZ9NIt3mMnlEu2QiTGmOdQs8kAYy3gd67l
nI2N7347Wp+RMhj+1A+LmRzE+81dW3S957XVrpF5m4X0EyTBdOJ6ry6LuuvyX6zJRbAnXEpWFvhG
FmWEoC8AVmCWrSQCQzdvXjL9P9mGLKrW9Bk1dfdATOt+0ir0e/OyVW68eYSaI71ej9z0SCi4rg0O
bl76FLswc3xiZv7ehiRZ0PgsGnDSndeBg90OW7NBAs+L9X0umdKp5UgBjfk8Gt9LGvJed+K9zD5v
EDkNKGsF2cdx3BRGsESdjXm8wGOz1HihyZrfL99YDo/A1V4ac8Baf9ABCvGOU+7ePxqahtvLcTAl
E90gSjIMvaMnLzs4kpBHIAfVM6MKnE+ydop27xUBus2Iki5/DA6eL4LEtu7UAfzhOTbUMrWAZZs5
/a3lGd+p47w7FvVOlX4D9dHv8w7mBcPt1WoFys+JHwVA5jpm4SqNu8ksA6hT+JvSMdRNTATKFAhn
LoJnL4UvTzwpkU/J8Q+sjXsKpKmmLs8n/NHWf/f6ZYjAmVRGE0c6LbXgRxcu7jPGpd2oGhXiTyN4
XGg2CsIghe3o8AnRf0DiKciqvA51DIYaVsqsjBE3/JK3bQSzngCdDWtm9GuKWECFgJrUsT01puzW
jmk3qbzu8FM41nv4z/MIki2pWJBXzXIl805wARVtmEn8c0gVf5ACmATNKSJYD5Q5zhYnbO1/o1TH
1hxRbI716IkgK2NBnDGryHhCow/9wHc51oSoHLQGXlTeEFPaZ/HbeT3WCvGgDN0QlHKPR1oj6Yy7
XqDOGC31WZLc8B/KPcjSwHMQkrFpKTPbQgJg74N0lS17nCb+7KYbczb4CltssfBIyEcxj+xzNUqg
01Y6DWqh2aE7R6dEgRHbK982Yf8fBGOChtctXc412u0ptxZ8IaKmWcqXGAtQJyHEOavwVZW2diWg
ANRpPRoLJ63ysox1O6gGKq/y6G8qO8Mg43FjBMNxZ7cpmAY0G6PPo9THBO6j7gOLMBKUM/9agXiC
B06MUrn2GhUfurHSfyAznfo9Ft2Br6btzc6JaOaXwscfi2iiq1oDegvqiWezbW5m3HFpR06db5oq
CPaRRbS0J7iVw+dy7auWk/f4zmAcGVLrSjWMEuPIn77WH0ktK0OB4cIubf+dj2dARq44RTwuigZh
m1bEdT7/K3KLgo/KBcFtIa57s4dd9CITfNerDz1/TBgLbvAliyC9RDyFdruOFzn1bfPsNFGsodcX
zXwVcGsY4AsSM3mbhz7t6V9FeK39h+jFSk6ql0n93TLWUVe+LaMamzTxtiZyzx2cJKF+YtH+ZHK3
BLGy6WGEcoXOHcUHzW2yBOJuAfa3EslqTVqNkCATbZ5+XkiOeBGMvGRnD9x1Qra/s4I0ftlkfEem
/SpADmVCq2uMTStidXwSAGw/dG3rEJ6M9+xkHdvPi8UZ+r/NDGfkv4plA/bHTKFcMpBf6FW3ikVn
bgHnv3H8m8hQ/iBXp1LhNFAqu1+4+wALTsdwmoXhI61R8ka0eVIZnZHxzvwhh/SCH9o303LRlO3u
yxoNIYVyOM0+h+JbTZzGG8T9xaPNYYqEIYuGno+r/2S2grfjhwYO/4rK2qF4ESzFowKr/s0pLdXU
7QdzpvNDv7uE7Y/za42eHQM4avJhosrWCc8XhJzPjmZJvYLtDTsP4rPKXsJA1HBSubp3836/cmVD
yNOgwWX70u6IQ4q/zURIQBQXyqO16Fzd/N58zsLuWRDH/S2qTXC155M93YASOq6NAWcZfMnEHB0O
4u/Wnl26WyLxBbFKu6h6A2ISQXrhvkOX3jJdCpc29nnEBTFN2AtrCNDyyQqs8+3lCoiMnfsGhGZZ
JaRkM5Ei2xXfeltaB+ptlet1grLTbn5jnasANlHxFi5j7xIndoSRy5RNgFmJU7jch32nPdrbJZZs
J8MK+05HAdxYOveVzmSDg6NW4yaawa1AYm7F4pmg9JV642ZZrihmk8bQ4k90HJe4sofT6LQ1CyCj
LJQSmye2+ry0yXXwHnHVSGJ/DZqLoXNd22Ny2lrwp3vhWsgVo1TOkwMfVE02c+TSF9pOzMfU3Xlp
H28C4BsVpNG3obLlQL2p7hFth3nwDurlxFNNXz+eluTdm24rdaKmx/3lXSP9Rw1LY1zkBQSIHJ7f
HuZl+hboUg71d06d7wnEJYwycOZ+ZGDnqvqovLcR+jkii1E0agzQMG/D5nvtBBWKfQe4ckSTNWbI
9ufuaoYw/q5DwEtmRIR1svKYRISxXVOKd2uA3KcQJEM7Fe7ZZcTeUf/V3G8kZpR56VEvBsjJRNPX
egtHRaiJAJbhQM1O7k521UNK4l99U6UV2g830jnFgl8HSav3BmGNTsKY5+U0w6UkKREIkw+YeO1Q
xnKW6crIiWG0Z78EPY3dDBsQoPG0psmruiDgRXDatil+9bYPyMCuoq5T4rwNf8PLleQsi+9XrqZJ
AnVAHgaQkXLWPHVQJwlGesofNKG9pjNK+ylTiSr+LvBly/4gXVUMpgF6Cz+owOk559Fb5wr1Ctfk
t1m0L3KerHGjPFnPYRhLNYWSA5keGEeoikZgkZVsmid2wVwLfy6uoicirBlgD1JyLuVTFzC+bpCc
UX8HmDRtrEjZ03N7VoZG27CbEm2bov0i3RLq8pUTIFqk7d0vDbDCPzynGjGtWSpVaDi67pQNTsIn
Ng3qd/tcziYfaO8+pA9aPAVsV0rInSA/E+F/N36tIHv8cubHfBiPt2VeFqydgcgBnHO6/hNxS6X+
Dqo8QtA4rb80ymOLJYwOxFDqcQxD23idELwxI6qcPMam3Z41NUT9xoMsXIP/TGYTL0wYyLuUNZwD
FU0dAA3cisXIQ61eByeMZrxOT3qQvNtqvMUPQbWVb9qnjUFkXMr6zTwGM9Oi10Oow8WZj7rF8hSj
ek5r56dxSFmIobRwL6WvvaRdb0eWqeNF1CPxmYe4CujkfvUZ3OX2sH1eESdQ6Daox0r9CObcSFVt
6NqOKso2/QEi6+zh7hXGr0zWOOjJHDXZU4FlKOETJiJ29zKR1Dgq5QPSwXgz+CrLpJk8bJqSBSoz
wMGghyDJRQsNOuKfZD0nvDQMatovEG/m9t+KJHS43b8eCGWN4/k7pTygtuCKwT3Q7r0jQ7RZgy/R
uGq0ZZr0vdMgnZ8GXx46wYYagPa8vYl1qgA9/8yffttO8790GjqLTWzT8ozDgsd5mXcFmm/5Zyh/
lxgQms+xCzZYGdBkMWPmijKuQtEIIH9DRJrxYGlbUpFxqt//qyXSsmGi2TFE3462VubAWa5zlno5
GMA+aK7cnrhhxGNyu8AxW6R6/Yhn1wIJ0EyDU+kBF/3keeCfV4HRsWLIDa1w0Fq8g7C0JBhZ7pO6
y+f0IStx1LyinJtTnhceowRvulHiGAcUR5tgib8MWIu0faqLu+e/JyG46EVdUA+AMzNXXCs2guLw
RnT6AZhp6ZY7ihdxAighHOCJJp/6U8nekJGg9/JuzU51Dx2tm4JkpmcIMBrEz3WWGmCBsbmj4bcX
empsBbzK13yfdr3rFpPoGJp/Q8cJN9vi7wtIPsJOSwBJ6Ppz3eZsNPqSssHUojtuE4AY227dtSAM
uGcN51g96ZVl1CEsgPBqcaxJsZ3QKP4em+9hvrKAYHZZp0KBAjYw2LCaSNUWPTi9khI2vdBLVQTP
fPTxX71i/65ZkhepDkLgFuwF2TQgkKHSkEb01LENV6QtcEPSIwVipsqWtjaR2ZqLx20pH5X1azJf
Jd/ZxGIFp63lpnfFFuwTTPxVdlFYX7Xnh6wedPA2TuBriyWyQR5urzw3BMiUO/1D4uLlKW/u46nC
PfdRmB4BACnlMndh6NLutQqbXsr+alMXJUKEzF9OXlvVcqMgA3aM8PNDSbqh+FUVXTxhJvjJA4mh
2wPzKfqu0Ivf1e4tY/HmpqZS02AcJ0jH3Y80plrJiAuvpmB6+vbT5vRaGSh6t/qHqighEaJock6y
/F7+b4ApyK1SnqRaPXULQjIqPHDtQfqncZTx8M7WoF+fHrnsCT4Ib0YTBZl+HS/r3x+4RIb0Ad/L
OEmH5LCZ3kD6szluR3PHyHdaqS4h0uDZZKd5eywK3QnIIHFSOMQ1MVzjqcFx1Er92AaEN4x3yD2b
KvIU51fEqybWYwDEHcb6gpbc8XyqDberFQAr4++t13q0xx+ewr1kuYfimghg/muKQ4VFfTwqB9Bg
FxHtqQ+FyuC8qSs5NU8FYWwHCf3vjSebX5a17Q32sGiC0zL8U2ht8B6C0QDrunp0mVE0A3OpaAqV
faa/cR/e8qFyEjQe5wIvaB4kqIjG8jo0fPXqvmLDFASvsnowys1/UAAudeleyGfRSqM5oa5ayox7
9nVwD7l1Sn++rRH1/PKUhPP0l4QdXeS4FpXPpcpN7FOhUW1GsZVWCbBm5+v6ldJZqkcbcmVFYl8j
1m7X38KQl929l3fk4/EvEBSSNEVeD6c6AZOyaj2Y9cvvfeuwtQJkCzSoGdOwMR4nKTTc7YrvAjEc
dWmBI/DRaaQrH4fxvYffdqtjAMVqUfKsDeH8zmvzR8ue1zSH3Zm+k2bRxprs45oj2Gq5rAxuEyTZ
eGB2ElH/HHodSleE1XoTsvIPH2ih0Urj5q4uNMAJsEHeTGiT7FHnLzHOfLwMPBuwfOIs8sB4yYFI
veVgdcimZF7z1SUZUo/1aR1ZL4fhMi+ygSgzfVTyvWsgdx8H6i4qKeH9K6Qrji2cBb0ztXBWukeV
qEVipC5COYyh0Z43wl9bovmutyKaZSdRpj2lz1DDa5T/LYU3dR8vgQ0PhjiGucRv1Il0EB05QrBk
ZeXbYFInjTjp1RM64YZMcZOvU1bPRm3t6EKm6FufManvZPsom8/Ow5uBLQ52RMjNWP0f8Olr/Kx/
AGoSGIt64/A4eLaU00mh8euDmOU+hH6QlyjAgLkPTTtyTw2e5ETH/7JeHhBKeXsGXWrYrmDxW3vz
GtAwrxCTtDCWNXBCVHHwfgy/Gppz+T0EOesmDbwNBPEln/Op5D8gOX8FpfA6QjWE2TmJvXo+Ci3M
Yrf2TC4p9eVKYmSCZTgFytRWFr81B55Kd1WdwJLmLBE/SUhVadonDvQKbJgnzkPHmWjVI6h0IR0c
3HrCEKQ2ZYVRMj3k0NKnqAM8bsx8PQve7L3eTcI1lZ6ZVYcx6srRaBhCJ4PctL4EvVc6noD2IcD6
c5ckIw1Q0TJsH6MglwVEe1nz5yb2CgQiwHYte81ISlA0i7O9vVqiI+ETd7k93VnBwT3Lvw6LfD7k
5pLVBOp9WXaEH0XeTMEFVqcwJh/4y30iAabtJ+PkZSZ8DoqognwLGDm5brih5ZMtoOnVhUiZgy9N
CqCw6bSzAvPJl+yhkKv0t29w3s9nZ6BQ5iV0UIcDqL698zmBxggzavKibBcy+QbUmXjhrDuZqMxe
PH1h9O7nGJBTntESREsrZyXizso1oNjtHFokEhFLW7AFOfFnYZbjMcFsOnBs4CE8Qvyuc/4BWom6
mhRI1kfb+vh410Xk1iE764VybjEmUDKUT2lXQlDP98joY8ogzXgI+DvEgDiNdiiWVIsHr1p5c4ao
FR2Pe4mSFRSjXksy+h+g2cu3qNX5WHh3apa5qlmGZN14sdT/FWbJoRXAGYCvtFZbgS3qGYQSoS5A
qnrpuzCZnhURK8fF/mj4V57+gwc7Ee9VV/DcoyPN/D611nb3xG/UPxG5Joo2OsHBtvgilL/mpEyY
vc9DaApaX2OB0VmpUOaqFStc93oFPcyH2foU7oK5CmESWHrAdbqXUTK6nRQmG6iCnt0BIXsmQxKg
Pq3Wk94qUwPQO5dWHhpgtV7xYxmaEADM7yJI1ulZ22THPZSIdEez26pm97KMYCG/uz2w49XwXm5E
e0I77xo19h+yr68bpnOiiCNukXnkNcWlzz6NxZVPEdRG18ormjMxgYNHzi8bCVuwJ/kHTSlyhW9c
AtzvInkUj6nfC2krTYD4//mC8nzlkHDDk8JNEkIAge6XacS7y5rGv/gNRQC1cKKZL6Okrb+6i4eO
XhUNS6l0ZaVjoDeWYR6DbHkxDnCVx4i33q/SudyPFVlErqFqKzNRiMdZJFKymdCjsOpBRGOaP7MM
2+pJ7bYffc6Txf8mHdv/JwQx/DXJxY3QrUjtPox/yGk+9yT1/L+Qp17l9KMN7DvdR1Y1eMCXIpY1
S8ICzJCCPl4A4mi2fH4cDqxZqWBIKTqrmMDlj79taTCle8gdXjcVjY+BtFxR4v0Pg7u4ta8Q8X54
hNJk+qEcwYu0zV5L8wkqKvpKgfibnuVWNisBvy8L6yavsHm5rrUt2sR7H8M1I6DB8CChNuZQK26f
4dLZrRCqfywUNMnI1I/v0pl/pfktp2mBBieklWqWgfFC43bVLK1vHIQNG1Fm+2y3Ec3UGKnD/pm0
2+sVKoLxMSa3KMD7giaADSiLiS6dJ1l8cfvGzsPUsZ5dzKJecIzGy0hk7vW9s4QGvtBaDsj14PhH
0armTE2cIXkv+BoGd45cqPrah9cCyoTepSwPz1WsW86EmfmbNuoMZXOpXlKI3fDJgaJysD7mCfWO
bUtF6t9XhOcRn+7yWNpZbCw3xBdz5dn33qADlEAeKLGzkDuDm//M3L1CRl/Z26pjUPH20wUJf5xX
50niu+bVb8utrAyAsseXqQHIKxmY1ZKnCtIUJ/n6WttYbu8QHY0S3CU7niubqpT1G2xfoJEUC5Ch
MIf9fLxXOp/g9feJiJ4J/DZeT/LPR7lj2fDL/HZA2+8fuB26DWARWT8+i0IlW2L1PSdVedFU/VQ7
N9kyQdfkDCL/iyUwGeXWJ16sfWVpdFJ7ToQ7rSqHHgpSr2czRu4CNudRdbNklQ+J5r0jwFtoiGyX
/c86fulET2IzNr3wNNi7DjOo97Ph/08Fa1TnlVJbcS4PW6nV1Ar5bznNQ7jYAE/6JNU/4tYdwfU3
zhIsyMX3KJRdwNg3/JHu+V827t3s7nD33TGf/Lrhp1vpgiVrO//ZeSE0ofb9Oi+B84lzBee7EqiD
drRoW6KWhHtlZe3dq2mn6ehcUMurUlXWcbN8iYpfrYb1WSrUbcuCXqdD14E8UaKIa+sY87ELTnpR
Ob5Mv+KmUa9bvnxUED1/6nVP/Zs6co/EAqSO1phfiL41BPzRAuD2bkNGknGuMBIdIZvxHX+Ig61p
HPDhnkGjciktKyy6Z4L5zRpTo0UDTmA87PUcDgHFi6Lsmo+ycbTPYx4A7p9R3MaYguq2ZJ6JT0Op
us4EH1j7yv7jit6DwAZS8Q5yNvdm517zRnOWVtRTlkc3qhbTxGLGP+cA1g3ugdoWnyxBjOJ7ioVr
C0nSAew09n5gK7/4I0gKtKekFwsHR5yu4Yk20UcGCjDiqR0BNirVEV+2ZsjZHlV17571tBY2QfNk
3nWfMyrmQLoRcXpIpsdCkWL02lzRHyTu0RdAwltbqKQAxSIzlqtIOGC8LMlzRHOn27iw8FtJ24Nm
Mc4yUZgLksdOxUVaghNK045Cn7SqoytOmd7xmQVDjzY7gQVkxhUx/nfY5Q4xbTNApeT0NF5a4SoS
aPbY8m6zQ60WKu6044LsuDtq/7TB134ToL1AjJYJHQn0Dz2WXe0dzZe16pjU1TuTtnPF9z9+zo5w
xUhYJQihBC4uZOD8GhPaEpS2N2+r3/wX4IRMmyRyzdXNu4mZEnGDrTMjbsiFoHLZx7OZzW5AMp+v
BbL0uTg1rBZXG8hV2vp5XKBVnai5GORTdaOWJXnKzdWrw5jupv3C2MFDkU20Rnnv+obfyIOf+oS2
ndygc2I3zjd8PeYE5dTzZjIONpoVqdR2Py7/sDlcOPsAREoQ1s4PlRoYfGl8FKeFqw3P/jSCWfQ7
3n589uMEKQSAiHpUpz0gFBLrbow1uOsVbCFfL5qVqFTauC6EwrGgRHxEMArVzZTEcON92Ones+KE
hyRACaaj6r8l2EXZ6K8N/NkiZspPaHD7+Bxv2JleDFGD1+B9BNuMGzKHXHyJ30IwDtDgbz/L094u
B7mOutcr67f/n+SnUmBoHBMNRzX1RwHMbad/GHm+2R8l354AXLOw0iCrAigqI/w8KL/DE+vZYFrw
ePoB2es7nQrM2DLm3x9ybcpdysM2g6jhjY9myY01SLk/9BFatXOa4x08PcVMhZYWXT85vMaLyFJI
cNgZu2h89Pkps990aP68pDvNmmoUEb84Z93Oj+6ssgieLLOSRnzW5X+UIn8hUmDaVTs5qvuYqVIL
Dz5h3xqhrKtGkGWHupwfyunejppOEO534yTjz6K2vzpAugQReUGrnGS3qVQ/cl83rPg1+YcgqqXA
eycPoL2J8oOzM+kmlLItM1WnE8j1HTLyU+GoBTEo+NgItp2zu6/C8z8U1Fn5CdEK5Al5sVl04oX8
6wgecrVhcLiUfWIzEN3BTV4Fg+cQi2xR7XtZZW7owNcRaxvzaJLWxxMsPZv9KSGrooQPL7ozG0Rc
cH9zTTJ8SIjDsOkPk4411IwnKNRifQP92gMheFYg/Cz7BaCHQwqcWcPnoBBbjRPANHRYT4lsGhrW
SypE6KPM8dIerXw9DQzMOcnb+jUc7WVeFOqBHo3OW7yLEHP0tto4xkDTnymHSeQWFsdkn4nilt6+
3ZckXErdl6iWEGdWnXufwVqdU5N0LHVKpeq2TwHajcHxqDoDnwuIDRki6eTVxrrJ1j+9UhOYIHq5
wgKiuVnkpVWJf2bDHnKEXNkfMaaLUAetYNbTi45v9R2IORHs7+bWO5XROb1a6OTIW9ZwcL/S7JFX
hcmof+g/L2cLp8moh9/dyYP+0joEZrfnroyIjSGHCL2f+mfEPLa+wHjUNj2exQm8vrHM4x+knNlL
UgFNC1WoexqBdde5hL5YXsQbyjoKkR+HlrAtCDbASouluSoCYu1mYUP/VEJcCwLdgTqLXDIvp6cy
EjjvVNM0ZfHzmRW+qzinAFmKqwotDjpBRBtvilOV/UEWDAPOGMBlaMPt2xgmXHFt9DVznMsQBZJJ
L63fK8uUvrI0jAMhn5kUMDWffXL0YwkkTnvEOZIBbu0WoVSaQ1ZWEYB6P7VsgD4vuz83NE9gMDKP
P6NBJJYfgTOTR7VMG76BSxj8Jq9/q/dmm6pcMluUPvHbF9QNn9l6RtugyODONQn022OwuQeCPgy2
IecVzi/JoWWu+AyydIKe9cFYHFnA48Qd+PeiYFNJXEy+qi0+3GD9SFFWw9/JkT3dgk7O0SbRCzQu
apbfn5Uo3Vi0cgEyoN+dFFaddEIY8JJGaQCfvs4Il5hp9PjqW3kSnYSY2+YF5ppurm1jlusUYQHQ
giZozdJWmPRlEHQMI/kHyfG6aIA07zmbxhbyNqdwE504TFxV99JUe4b46LfBFGcalAQqU48a33kF
mXsy22OkjpaOVt7S956CjV40y965kxKsEF49OEja8vKbNL4kkFSzq/yQZXRrwIBryI5sxzVrsYZ1
MHj3SYF1+I5tQlUsdJBoyKcYxFEcuVzm6xStGWU4AvY+wC4CiOIoSrouNXxImT3qfA/IkHzOeYtH
c57UjR3KHIsRNrDlWq/RHHwPH3alugT1QNrEQ+/gwcIJvJg1MoA68bq+E9CC8wQITuIzkalLAUmk
ctib4rfTLow83X38Vwig/gNIdKJd874WOE5V3avz3xzH1tqyYenIfTEJJVVk6iOeGFhTYzU9KdRE
QnIe3e5VcfX9jU+WLB2D123q8u1bKYvjj5FKn0V6+jd03aXzYIFBaDLEbbg0mPLFzRZWLKtjMj3I
c4ICetivXxn+L/KYq8VlBCEMDOcHTSO6AQT6HrPtvO3HOUqLZs+P3pKVbQ0r4mdPaYWY0chYGbF5
zvBf/S6B0VGkDQgK1kYyNO3rlifMYlClFB5uYL5eDMgMSm1YjH4mqvHUz3jqMbB5VeckVSGU4/TW
Cl2HEnZEh4vEYYLBEB0DBDt9d1OAK8dzo/t2WSU59W3Uzg1V5QxVCEsBzgPWWnaUEdI9NwGrx/SX
H494SwfvAoAcocNs0gY6Qz/JJ4iusBmOU/SfrnyI7AmObG2X2HmZArvobeM+ijww2O6ebBnAnJ29
5IsqEuDvSpwcykO1pYKhCtD9pq2SR6/uT9WsMby626KA3Zl26VpNLUFqtWzBIKbllsNnYJTLkzUg
MJ+RTYqJLe2SyHtMVFBu8hoFToRG8S30ut2DxJGP+B/sEhLBlSul+hoyP6b0eiAzNkUcqnYv6dyO
LY8N0ARRjI9sgSGZG0NNoL+DLtjIOtofS66Dh4KdF2/kM9DjCvDRNDYDF7LY/x+7uJmT3IWwLNA9
y2UgyoIeI7zuI9Tepk6PcWgcbY2n9UWc6tpOp6zC3XCeDd3C5V8I+Ygc95Kz6I4aS6IjIfuAwWRv
ibsnrvxia19sAKaZSSbMY2L3aXuNGzdEx6L0km7ZuR1OthPADOE5NSrcj8HUP/gWRSTY8UVZZB6G
kcoyMeYLwl3MeM/L98o0XgbgXYjs+dzHlIV7rWscAFrdyBFMOOHRrRCfq2BN5QbTYzs19SOrf8cl
h2Ur52qzaMp7OTF4LLbOqgJPKPz6SB4awoimnXUJkZVJSlnXeH0oL98oJqn+CcWvD95WxMUKGwzx
+kpo8uEKbP0or9K0biKYDodSYze0viGW4TujW9/CxFMGwixi+juZfxwmu6zXTDXB2RQDpzIC9Df+
GuVmhV8bjzdA1ItR3Hr3u279f9ovpMOt2StNdwXrQWnarhzYH4lxYlDi07G9LOxByC7dtHRmf1gR
FhahxqdqWvoXazIzGNnsxYx1AazBIJrHpnxN6IDKEeguQkx55jCcCH/BbLatQycYc14dEePyTGvz
geT/qG54hHl0kpAmfAicgwF2wuLxYg6N7B4rZYe8QaHp9vo/4ZA2U7Jcbui7GzM+o5D+x1S20aH+
aG+Gud3fXT6ZagCh0jKvSILaDZS98v7j/h7UTiT0syHe0RzKHX1mCazFZn2m2b1jso2/zdzspQgQ
1B12ZAlQkIbmJavrgbei1YXWpCM5tdtRTSESe7HKkH8kep9zywhYQ+TDRiZ+imcgaLAUR6VyfDUD
PXV1UtCfvTxPKbz+5Y3fA0Kar7J1Wo/HX9qqPoejY4klkc+DKhG+yQZRRiLInMns0cnt9GQv7jP8
XovKfZ2nJLYnVsg2qQIB/VxBZuo8R7xqPG0oArapmNG5Ku35W3ebll2qTR5SyQxvq/WTYf5laDpu
J09prRg2rIeif9f+Cf25cYqkTVkbhJ3ecuSFZTsjTT78/VEjJGt+stYfNVA2hMz6FPIoBVqckZVF
u4/jRslvU9SHVfNOeQK1T/t4QnULcHfxK6eEdt14pt52hi/AhrOjnxEMZnjI0EJj6lg5tNVamOzd
vJClVna/5LdKqG9JQT1B6d9cvTcgI2dVariAJT+y+LIZWuOH1io7s7HrLyYiadXm0QuRs8JWS02K
DyozkoxhUMDh5ZUEm+vzmh0qkIA4CjbdXkTZ3nLSfIa+Z4ug2Da25huqaCiTyNboFmGnBDJVA7e3
AfpXd1d0XGAzV9d78VNprope0KVxVShuMVR2i3n7SrhtBcmbn8C+AW5X4kt4hLL4lI+zhBSgUo05
B++iQf5qYeYmyuNylp5T1pO7XbUEsJK2lg2ikDhKKgJ6iZEUusFDCbEktzyswyWz6CmQTRa4IuEh
mSTMN+jx5SLjHVLxRMNLj6XytbDGf7vcg7laH27NramH0qlXNwGZ+oh21TgxzjDrp9NScWVq5C1d
lIWWYo67Nj/jyfpZHSSFqOYmzMwUE8EJYInz+PZsCIol4sIYIARwkm/l2B571WgL6rnCVDDOGu0a
6Z2OGudh70+MawhaBNXulXSqyHHAeEEsFZvzmSw0xpVgC+ZuLpu9oZ6XQXhUCDoF9ekZ8GRnLoB7
/s4niB6nKGHyF2GIuDIPLs9g3oeIrWXQH/dnoQfO1Og07L5kOWWoe7nylvbbtGEbxIwvbwOYce3I
4xbS0mqQ53khMJsnKby8Gn0Kv36DDEDaUrCkwe7qoyqg+LHCBeQScWOhCOWTd19GSspvimgTC6G2
ysm1ttEqr4pHHngi0iUZOZrhsPwqQ+EkQEFMMF4jbD/BtppHQzjo/NgXxtMUj7dGQc9JZrS7rNgv
awDozUrqN1TP8zDBnR8L30/mm3N4DUxwg0S7CHhngyF3pX+aggISbqqXcKpLu/dlupCywsSk63RX
08oFcHLQ/9LEVcw+6cTyeHEmnNGzlfuGrnqX5zuzgm/Hdq9s2hLFyzyo/SvMUNh3d7XWLxZPjsDo
SQXLeUxu33efLrLkXcMuE6NaSDn/IL6uxn2GuJMzuObCzVPim5tF2r/MFLDcrtAjcwu0MU8ask+t
thXVT48Q7i+YysOHd06WAZW02S6vZi2/v9H9bzX4cupw8skFfhn/cGUMUBlAue0ZBDS5u4pt7i4U
ead2WEqEe5musrPTgsB+KbH5sQ/YBzABGyonLAn4ME6U3YWX3p9uxCOxGhXREaW0OrD137pXndRh
tpSgxsSqLfOU1QCQ2f3fGTX4U7/2bfUbeFQiBHgEyQ4xalkzaeqZWGScn/9PtLOMtz6OqBex+rOf
cZTT9daZt0jXISERZoUXJIzJXXPi+Nn57vw45jQ756T0PlT7K7p6Oq0uwnX1aQ/GN8M1r6Yo++Eg
RflE/9BEXbKCdrrQL5iX5QJ94Yf8qju5EKVjXxhHZ5K9KKDDTE23BtGpKyjneL1u3JcL0NRk2XY3
vC6TS0ZTM20kBXc3i66DYYEiQ3oNsQ26GIlXudz2aZGw5GwQgytCgW5QMUWK7GynkE18/jJth9H0
zdap0qX0zDaadml7RmlgaueFTEV6f+3tuuilhoPl9zkzOMqpFeEgTCotyYGUskMUj48ngJ++l0KQ
uNIHXLFyC1x1XwmqlNk3cNwUHC5CuXf9K/jwQqj5PVc+ovNEjiVD5GlawQuZlmYYOR02I1k7SdCo
EhacOWazBw2j3J09kfMJ2VnMEmMNxMRXs6ZQMoZ4G+/zMtVOegUyPXkANBJT81TvXZSM65DAWRwX
YwcuQagQ/t6G0bbHgADqNbxeiJgvxRedr41etRP6y9MC2JOjNhCMmKTeEPRvWZsrSXiiM1dnm17P
pA7qJakZ1qvyjpwI8/YQ7rq0sc3iqX+SZEA0moMnm/W/ThBbWE1WKZYYxiX99eqY2uZQeVLWfN5X
lCshB8gLL3q61uirNM8Mqsx4dKg1ZLQ6xI5X4JZF/N2iAW25f3oGQN2PZwEZLXGDrrP4kZiYd48R
Sjwf+ru2c4YVkNMT3UQ6cgMNVO4iPNJnItBUynnqU6FQa2dElAoutIxopQkfirPHikxuLEaYqGw6
mlcbJngijWI8clMTgFKQe1F3kF9WCXLTynD6umERH5HJoYU3t+Mh4I+i3k7GMSCIfKkO1r5PVhDM
AKwE5Os1g2rC8TsrVfy/BoeCwcl1AtS9L4Sq0VUFUZbzHGD5RAbtQB1r/uECNe0POMM9u9JlxBvg
pf6WTkv2TlLxUBOnaFp+j7jK+GhNR5CazXup6djtJ5/suOtYv+GorBSevRmf2wdD9Gc6r8ptDNqc
EnZGyXAUFMGz6HlEUsaYcmQGhs2v1Zc6tHPDc9nwVdDEQLI81FnIQKqW2PqDg+d46HJFgEyRfGHb
zouoi4lyxy/88bcfCCOwZkZZG2z778pmQYxWyvLczNGnx1KL7ko2XMlM5kyY3fD9C67Pr4aeQfiL
p4Aa1OvfqnPJzr5OxptLc5W3uJqe/mUiCSvVGiuKqMcaXTstRZ937QctAPx5xVaGIsTcfUtaw8qm
YK6uzafaes92c2Sv/0IrPhzOTusMRmx+C6xVq6WDimSA5b3x5vBtjKEumBAdLlep3/JX8HOQzTf/
PxX/RMAPPiLw/CvIyUTny6RfZDUmnwKDm00tC0k4NnWZXY7NhZEymHP4s4Q6CB9XtD1FrMRbr6vo
aV6QXy5VW/3EB55VDIJfGVjqnnk7gAxK2VS7EtEeFITkpL3uRWIuwjqXgQqAWbnwx62TPiILV6xJ
TR8hRMXRmLv8HZyDPOyy2i096bgkpnCtp9MU2EHmdR4cTznNUgZDscQOY0bhhzjycRBrIWsoqaKS
db/gSxwWQxYbFhs1h/pkXdolft5p8KYTQNTSGKBYow1upWMRnNqQ54rW98QDMFXsJeC3AG6tatpb
Ss+vYLd8BiEw6T2gNbjRnzrwoN/O3oIJ8ipIEHzDDRo1pB5OW6FhI0BLBbR0u056hc+rMplqo33n
B0SzkZy90YiU+qXtxp31i9khTQmm4jP+emeOLKTKQyiMbaRN4vvGLxX7meEf5QhImRqWMhb/8gY/
JUaTJGIIDUgJkirvMSl/4z06/apXBExVtu6HN8BFJUtrzIpt0pSIV5KMIYLLrDLKgfiGtE3e5xdq
t773zQ4XrHUSdTlW4cg893dOAbGDizEIW0j5RYTM1cSEINywma+nMn87gWnHGi0uqSe8OmrDdcTP
ayhsM13v0eaD4m4GMk9kVyU4dpZv8FlARocqBUtmJeOgOqefv9MHfjZD+NQDrQw+DtK5eCmPql4J
cOgrQI4sI+SrZe1pESzKyU+zLe0mHjrtSgH811czLieFdjYhELawHP5dlroDgGaUKiCDYEhGP7pK
U9nGj0hCupmtQeqtQlFJZ7KYmLRhhaB1w32O36Hjfug/iLBEZvdlsRfIt7XgbAjIEKEZpGTEOrvh
tIEVbucWYZmCTLGYzEev0GyZIFa9rygF2iMHnxuClMuP5PDeyar4EFMvOG/xp/wEt3Pkd955Up5x
eNP5IZ94KE/n+HM6EALXNYAVQc1IQpTXCMeWy0Krh0v4GHfsZAPlPLXJxmVZR6HHKfYEtgRbKuTR
A0e93GYyEO8y+NF0pCrpwHOfW3pyTiiCmnxXcnZK4/UY7yVVYlRB6mBwItsgwmHPFNxproXzbmgo
ewUgPFsNGxgU45W2JIvs+9i/I8lG2+Gy2zWCFqmHPwQydpVhXvsfEvtJYjzYxJF+VUgEcW6m/of/
ip3OLZFdDCAzY1r7aGS1lJs99Kf1Tyw+oACUrFGUDZ8WYuk/BQj8PFIq4U5Txy6uSB+VsEitw3mN
r0T2NNvZdPwLxUONEqs15TzOZZsr6/6z5neAHieX9CjM8ws+cx3dRUMcq81oClywhCHTbO33pAmV
edwXWobS0OyM0cj5ofNL2zt89FqDIxuTJ0fTtFXHwFJAW0yuoNlccH+z9cvwZbEXNmYJSnPjhbVc
r6B768e/Rc3oMVf9aDys3rCtMFjr0ydU4DZ7oFlPoVDIKYGccwpCPHWQoU8MTQzmk9jvKY81gZ1x
+ebR6+SSBY5Y2FIOMDAKV7NSFYimEGrsnMoGVyQ+KvYVHe9qPffWcKg19Mc+pPCdsYWxyes+TnTg
3GGvfv+IAYNO1hINnIyGfjXJ7vGbo0lXPbs6/QbhFfAFAnCIdpHQ0W06yN5ikVhc81iDliwoXeug
ByzUFrK1M6CR01AvRm3yQBu6GEoVphd1oEVarzTM4GIcWOA7zy1cHDxgHOYIEjJPtyZWnU5tXHnq
BIQX0c0UlG5cUk70fFHZZXuadbQV6b81tRz0byEW8trto8JUf/9bBwU66iNFtA4KaCMlcvU9NV32
ZGQAKOV3Zp6lLHSO73QaN/Zmc1+XuYi6Qnp67DKWkxY27GLVT4x6FU6f+axW37rkkx+5sKKILiKC
7irQcpaGBUkYze6qcsrScKrBjwru+1qRfycs/HL/iaai5xDodue1TQVwhb1E8JfHv5u7JDx/GDJV
NyyLpeNptMuzOrIGK4hDoUO/wWBtO71QBEJ5JctdMMpbFxF4kxPKpzLxeRPDtc7gtwjb4DOVnI3P
K+HNMWsHJYTOLYCZqNyEgDroKztv1Uou/i4SuuY8VFjUJmXjQsFt6uxfb3vOCUwGxjeBjE0g1XaY
ZPiEJz5mZLq8xd+QGyYjgTcf2H983lJ3kfE5JOYy9r/lUQWbVo31Sw4oYNNSH8W0OXDi/hFBKvBQ
9J/TdMPAPnqN6RkouTQy7MkFfdsJPLiPH6SpwAZuohjB20hlTxegNStez6hXVggeu8E3AFT50DbM
Z5S7Ybjmo8c4Id8GiVH2tyGpBvNoSvkj8A6A2Nu0NVAeSq/zY4LDnF2syXVO8pTR1Ee6+8ob/0At
dZTIVcgyEJjXajyrg4DaKIgdZI6PBwY6da/mdxVq/NRZS5nQE7pz4pdONfjqD9OGBe3a0D0gNwqe
O78FhT22RueIyJ+DAqdDq4a3IceY0b0G87OR7RLgB6wVrBtXkFDKs93o3uofQzNsMWfr9mVV8Huv
HZL9mGU4YRkfHnaVU6AGO8C4lYbwJ/gUUX3vmKnsHmOXjXe4dpCwA0NULej12XHnzBconRwmAUtu
cR23e7xbFQIUJUFs7LDj4Ul9u2Fu/SrjdcxSu6BOY6nrq8Tv+MXxiA7e/UNuJcD1O7ILJcx799O8
wc7gXiiGSKcZjeWGYFPVDZR/PIeq9h9MqQtHWeXh954JlWvQWf13I0HLOEPBqhf7aorxyh2N6zBV
bwGhQ5QWemaeJHTSsLfqV2mJQXxHfmqz7Hq9Blx277O7kfmQTqljr6TMclUZ2lb+O2/3vO1EcP3l
bQ5+Qk6RdUlGvtpNw9WTQ+bugJfFPC7ShWqrbc+FPyfYQywaGQ7sTIayXChgEVdx1JWxVHqsidt3
59zKC7B0rqiTTbUrV5g5XXifAHx+zxjoINB6Z5AZ/G0QfoSs91ljKvZD/g5dKdNPvOb4aUSFng9L
Q5zDJaDei3FoRgMwx5v+Pj0DfuTSmnb83McLnvLUf87/RQKNKOXUnQadGBctL48l29QlvdXsPpnM
XsCdR9S3ddIY8ld5ODjjLe9N/8/skahLTGy6ewlJoMRbz1QuqexBtAK1ocysBYy6smpHIp//DgUU
CVoPTGv9l5cpc3+ZibI6fWKO8QphU+D8gxkBynmspk2fUqWrIJ1DMeg2HpeA87X58F+ukGk3Ajea
gOlQ9d+CBL5lTifchXKafOvLBA60ezASrgsxedUgqXddpwrt7UqCP4Foui9DxXyKV5OPJKG9sQVD
MIfBq0AiWCZK6NAi2eLDMVaaZ8EuscNt1ya8vmWBM+VOfx5dfxURdWINoOYA70fgpPqYN4LQ37aO
pG1csUx7Mh0wsdpmBsruP6Y5IKwk2u10es/M3/4x/8qQyxaKoCQQtEaqbufaIaqXYdpVZ0wAMbZj
187u00JDQKM8VqNudpGIrHRFG2KmtdFEjyhLo/OYVh8lhydvmiPeeCHU5i+5WJOJ5ptK4+eVE569
3YjmzfwU4K6KwEtXstVLd7pGnp/pSrxyksk6pi/j7gg7j21yO8xV53ln65IMrFQg0n840E3lRVsV
S6p3i/z9XPWf4ibH6BSkitGe9iDfkg7oeJmbHh7pIx00bCx+45rbdesbfKr10Tm2vmMeexzD/CnM
WZAUgtYpwLNtxFxvS06RJ8Au+pR7qtLmVhlvGI5DMqZuuTsg3cDwsmAfw5+AEvILOLqESOlYd8wY
lJykJwoAhsTUvIR/GtBEtZ7Vg+7eri4fbZP1Hy5i18n/2IBNi7keTWgZS9U+/j/kS4KAFojqetR+
SvGttyGmN13LFJcGwkFQS9KQtPkUK0OWMRTpfkSLdlXhgQxdh4k6euEnA9u6wXmU45bQXIkAKgTh
e5Cn0xXtxcyJFHbi08pGNyBKhdOruuzjAAIP4+kjskWfNB4jpvpFpTJ+Jh6hi8R/Q7FGgD3IV+8p
hmbghyWSPkz9jDn3RvZLsGI+LXkKwTd+ADI2FlJMvkgDXpNz0XA3tMv3LgtmVAedu/QxaW4wAUGf
LCBJUBW/+ISvowYunJtnMgXFTcUtcNIsmigWV4MPqfsHz5chanrgbEViLWPktdSUE9/zTM9iEjQ1
+579Gn5uSr3WEDv2EyWQZxEKbMg1n+Gus4LyHtDDJEEGnxKUxFpDZpRprzwXpzX1vVXZ0BGXsyLo
Sg+lggll/8tuAVpc63AQkrP2x2QR9iOrIM2mwoKWOtmTMD5ZbXdAr8E9thsbYYB2y+Kz3TVKSftP
/kp+UsuUA3Tewn7ctI/QbwqbYGM7GN7GkgTmOU+P1JpOqz3yVkr1KXy3ai9Q896nwEagVGH6C0J4
AJKNQB/oDBoja5/J05/rma4qBPF0vSuKSfMQhcLynnKlSm28A+xdrs52/Vij5YL57LOyfxKo9XI3
I0VGRiJm/OGyqLD2G6529vYxbusL0irXSoPapsXsEIyLdRobMEwDE9L7KSCRC58zCVKud0A8tAVr
kN/aJZOuPGaHExII7hrgKlzll/AsFnWUXSnDBiWUQbiCNEMHDINgOyRVu8GN3JQZZhDeRVSChuTW
DIO7XPJHtBA00BIyeXpIdaOSol61/3dAK4IMxQWwoHnJxtHhWaz8PkesDbH76HCmdINIPtJNWIPe
VpNBbl6CIrBUn5Naay2PIzv6jZRpyQ4RiOmqwDqnt+Wf9L4bAK+7vn4b+htY45hi5G+6t27p/pRk
rJ+KTB/RlrSRQ20rtms+N10dpqca9JqR18iEg27yy5eon8ZJKKqbOsjQ8vbAkK+n7UNax18UEaOL
K8d/hBrvSKsDhFQfC0AtPd1Lw2uPYPA8KNcawch+8ULJi2hWftWglnRdkRrD8e7QlNIn21VDFCPx
+ak549bvADAhLoT48j+FeJ5mtJe2rSEue7bxNtRivOE1pRMwbu5s4gmDxlm6DBdQpMUTw5vhyHca
kQr4ZThwsXfy9ZhfvXdUHCWUycE76itJWlbPixVjiercYCBHQZuJ5FaCC/pZTmUswjN88u2KrWi4
qjNJISMuJ+e8DWaM8CSiz5H0hNK+9b9Pj8XlipHDtWiWGcIYI9VTb/u3P1n0l+pEV9U3scumzSJs
ypXUq0M9iv2xraWmaClySZon7I4rSRdweaSaDJi4Na4W7T/CexBDbgXhFRtjKcMQ7wF+0IixqHUH
7SS6FWzc/RcgfTJxXgBX1pp2JpmZFMyJ0jP6LlDY1bgn9bySFPZewCfCnhRrOpsk9R4ouMr3GwQw
kC0zirKFpl+r2fskrkV5xBh3o9V5Il55qHLvZgWA5ISCh0FmuWdOyGxo+lQK7QOtoWE5IIW7gc1s
kJkiSIsa9telEo9m71UYTU7AMrsP+9+YoWO+LELYST9b8OWSJMxaF9E+YcLPlRuJ5MpXHVCDJvfv
3Zv8ZZcKjzYdZy0AnI9GxfXZgTWdEXeX6JIRK1QUDdBxM6FbMk2AyIVQrPSY4ffdBGRiq+En4W0+
gioxylqyDgVO+oK+HHfQKLm53+hUusfJ2QVrOMIlwFtzZh2+lvahDyPIu4mY+WKl5VrgZ2fx9PJN
ZqE4vF0miVZpsFvpq5veUXAaqV84RLM73bH4UjDxT/8EaUoh9U2HNZHDKRMrJYB8isqDgIK/8oQ7
HAiU5I9+dX1haqRCmbiXIKihYm1y6bFNO8HNsvu8XomxifDmDQH7oU5wUkkVpedWzqHO365yTiCq
WxGbTJa5z/bMDngYGOhR1sphomAZaQH9QjmCgYNjcZ38Rl+o6+6ucNlFzGhBY+FwHefJcJcH6zi2
U0/z+UUUkSrAHo341IRvXWVG7Ek3Cm37RPagevSgo7gmXOueSt2rSz+Zwp4HGBNShh/XoIbRExe4
wgcnagn87orq1zQN8oekQYi/VP2toKThM7Pdav8zkP9kiMlq/CSaLI7Pq39i08t3K40b96GrJ1UK
lMf4ft2aXwcjE7YWqogNKKhzORpPmszy6WckKrkpNZaOnMcXR3BTjgnDrJ36GEQNmBx7CxYBwsP6
9jS9a/79Jnc5Tclkjd/pu48rtRhOSXSM9thK3FwIUP1eykyPQmYiJtWSPNV/88a2uoXAy1BgXFD+
VjtexgTgrIQPGE6/h7+sKOFR9O02vo816jlswmFcgTmfR/lEczRMQ6edFLdcdGVTvxdOroTqUKbR
MfKGpl2ZJNsJF4JDkhv2OJb+Q+0eu7alDtJQNTXgo0k+WGyRxMa9aZdPO9rNVKLRmfKZ13wAZB/9
HEAZeBy1LDL4do0V+i9zSuxannpOD3mg4AeVv01QiQJjAJ0YA0z3d+drXmqIKVoOiaEgzt2nXJHC
AD07SCGso/XgcRSzVY1GtOjjOwwoGT4imtvkvZnDsebgbbFq32KhskNGI/Ai2AgM2F6m/O9Puf0K
2DJ5FgFChi4C3LlIDiHdCc3e+R7XZRoxUGOW2l14Gc0J0YTw3GZwfNm5Xxs0NembGQCtMAlCqdVZ
DRXUlDvTu+rlJF+kvOlCcdQVNRgEUabPHuBjJ35/m0Suk99SZRr9DR4IZTJWhhrTPXDE3rgu0h7f
36dxFGl52xYIIxlalN8m+FDwXfLx+UntS2ZtA5DVhVK650vW2D7Vmc7dOwAvou5Gi4cUXN0sneWk
L5xcFGAnzmPLqBw1zojFokrJQopartDqw4pPKtMwObpZWWlCqp64gb5STHUi0Ba6umJfXiGrWwkI
Ut2bidZug615vnvG1LdTyqc7FHBEZrXu6sSRPfDKZgOAhkfvmUtTYrakpUUYG9Yg2+gPKwF5KTp5
LevTKuXRp6McoXekz4Qgf6QZ3IPFvxmiKMJtsOCPD1a4RnCJ8qQuXFvwfNXwZv1U3EDuF5OjB4Gj
GDSTo+bEcIG408c5kdVDcW3Zh+TKWtokhJAdEeKXyS/eYrwDWMVh9pS2D4aLozzmVc7RiE8b/Ld6
PHzjfte7nP2PGZ3E9QUX+5bWgbZwct0gSCyLsRjiCs2Umt2/HbfckXLjr9y1AiFdQHjCmu/Tj82s
eZJswwfZLAviWurN+9K2J3KAeMJ4v2odtgrT3978JofYl0Z8GxRlfeRX0odlo1npXxtp++X5p07N
V+isWlh9N6KV065q3eZa4/5+RxVIeoSdVbGwnlaaSy/lGOsuag7zEyfmO547jfbvlkb2vBn+OW33
VKy+FdLfV5QN0c98mLwzG2+6dxpjOstNowKXKT8sYQEIRit7FZCEULGj1ohIAph5iVZIlbv/rAwo
/VJEoWAAZo+/9CuN04BcV8wFZ1y8KmFGfmnDYyA9hJ/fCRQqTTjMBnk91Y5gVjf/PZuh6G0Run81
6gzNRbTvjg23umvWEC3VvV6K+h09zrPCJ6Mgf2/UDjw1HSOwngPriwM0RezIPQ6UwTZPC65I8AFe
a0/D+f3y+vDlmAnA1fuqxddYavbnPeWOBPHwVGoradrtuSKmwqtJfztDhN3MMLx41MerBn6R/5Py
49Sz1m1j4rYsax5jAfLobQd8YeOcFdvEiB9/bojqXf/KZNMxjnh+D5rEVmG4lKuf8V9jwe3tBgQn
YI/pqLRRKW01S6uzmu/ripeiXr4UdHNf9unI3pl9EYSM9jQilUbgcC+7ZVzxa1MfvRSMzT4XdNI1
LqQm4hAC2r8wJvGSJWxmFecWHjpGDRWTDg06YlAwHL7zaHWz24LjJHmFjraDfzpwMbSehx6tVHEj
2yAlOXtgpjDQ6NruHAGjO1W0jeX+iedTBu1OdkIRB7KCbW5Ct6dBCItYP2wdogKxNPPw/35nLIle
a/d6ij5rVYMW2+8Z/pSPLquscGQHlxh/TxaYZKFH3HzjaovA6syFb+ziRu4MEgJPGkXZW884dWyf
1UWYmynVsTS7VDLUfg2rYzDUyyK2GF7VodGqcrZ+9U2V8OSu7dpGoiJLe8mcAsKmcPrHzx1u1pIs
N8ZbQv6nL4brcHE6HmphSzBfblntNyeI/2X9oK21xP1ViZj4siSUkVU0wTmbsxxSX1YM2Vptn3Xl
YLMmkxOgyijXSR4KXJU+GpwEgzsKJNq102glWwEidhcGxHpwC4hCQ8FWOSrAe7PnUcd6YLTd8OJV
zJs5Ul5HepTvee1AsSXnnRz3WYHcGqp5unUoPVUuFxafv9bAmiG1/O4sFdRSZq6EvlpeSChRFRrB
0EEoUnFJT92YOaMnk7OshfN0gBmVGgAtdKCWaVhOId2YrARXIBX88c6MA5iYkGFxc1QU9vtMJ9OX
vwlx04KJNKZCzHgNYOCKg3kI2k6XU6hOgJMaUTqWhnvJtXgODlihxUKKdZx8wXyRyZ9x1Wu12GL0
vG3r2v5IlvoJgb7CJ62R8vPqy4kwwnA3qLfEMQ8nPBBYlgMj3ljQYDLU+Y1ru8NYSeIaGNToAbar
9EXvFzBPHkXG6iXsiJV7IhcQfdXEyMM5k0mYbS8G8Mm9BHCfPMfxMKOLVc0xYDj8wyT/5bdBG+Pa
dERS+kDuLRCEZHlzRpa6cZ6Q0I8W8XnvSNBPvekFDTTOPDhu2KJ3fx5MGduYi0QETFoMKZJJufdW
jG1p1eJt7kEWkNjyIG+yZ7IiEmVkdMF9T4tEgio4+nHsFMb5f8PByjth3o4CR8ACjTVdzjyaf5Xl
18H0mJxBWITkAhryxYXIo0kwlqYSmKBbn8xKSScpDjPhExx13jljnRZaffbdsAFAgyYYKL9BnbCk
BODEqyrJPmX3hnd2R1Tk1TMlrRYDO7Doy7acrah4Zuj6NKszAjNo0tqemF/8QPs7GqpkY32y7FUo
TlHsZ7Kr6uDnfLrNsSXGLSG5SzLhuB9ovvGYvV2uvSx19KvImHq6ZeQL8lr1J8eRCGfPz+u02g49
4XCRy3i1UAPk1PNiIdE49fpDJpKKcXs5cA5wEp2grdjSETA6O8H5buMnRfK8eCO59DHXyEYAXQ/8
RGqn8zyfC3g2/QJvovWYChbfuDoertUS4PQfGyc3uuXcD7bZaMFJxDdg1Lnd4NH7xGYcFBfxpTbv
e/ArftYqK+C4BgnWdUqJujcSeEQQOwAaKvKVJU2Vxd5Yn1KuA2TKLMvLE16/ZxkTPioeX9O95GMO
eif2O0KwBEqcUc9z7/S6MkRtk9jXAuh5tbq3fm1PnFh+AcDgT6B8wmfQ9i5biCHODNavfc/qxJTv
fNr3p0lcsRv/RKIzwhhckuviKQvWZNhcD1dFa6RFEslwOa6s/4CZ0H1yQo4j3FWCvQOlB54+odjR
znEI77tssOteXOlGJ7m+iVNyTUUFLoEpm5gHF9Uo9x07oWqIVf3zSzDJflRF3SQ2hl6tahzzb4pm
gmEDNAGlFHMsez6ImHk85ztl7Jvo6NDQO3vnmgruBc8Y8/UOMgSij3k2fJt3yGHX1IeEgxnKx2eV
UNTVy/6qBSGtgTBZX51Xk55WRqJw29xogC1lIIK+Od2anOMl28pYdXXh/K21HwzJfhO0YrZRMDb+
Nljd0b3tAScb3g8ASrALa6NAbRO0cdDbo5qVoUqlOcb8/1U39OjtkmuvOGNBT9P6GvOZepQLPZ17
3NLGylWylEj7cevt/7B4PkVrD5oIybgS9PPvP3v9HDH4y3JU8/hnhk0eq44jShDZWbezSg3xHOsF
2JbevsZMtgP6IrE1ixFMTLZGazw1dCw/n656y9pH+JpersHjUkgWyamvnkH7PzT0k7XF5Bn+2LEk
Jp81qVdfLtXmu7HuNbGU1ustzbEHz4BYXSqC6s41n5+TBzP+4DRknuIdOdHpIjcglwUx5bykR4sS
dBzmLrpHBrGt6Jx45GDj5Vbl+WDcv0CCEcf0RiAGOURuBM7HqhH1G2bIEoSg08+cpFD/TcbaEI/B
LOGxYbRNbsBVALM6HWtBa8vb7mOxOxcXyFmI+PPdz/dMZ+ym6S0HmRKLjNYdVyth7TbXOIkuCBA8
9nw4KkIifQt2NfK+/cwEO9a0v18xC9oC5osHnz2UAH6VbrfW3Hf/8u7u6ujo2wGmRHmodmLjxmBU
qRgbObJe2MF8MpsITAvOOkKnFvf6k+D8F859wbMgCT62eRV6Ckx0nvuFntxAbJrKHOQuAEYzRPhu
lNZv9jSJWuXS05vcWBvtQfwIZDoe1/StaUGtpIlFw/JPGUC0o4ox5S8tw8PSnCnrQbiU5XxzYpX2
WjoJ4z04XMxUJt90EvSMZe3SexCncnztYkXPrvjwhafZKigeZddz/8zGpX0Ldx/iViEpKsLINilq
96rxKS18H8IfXkK+3FGh6j+pcUW9mo6aUg99iKOdanyT+/wogxfL+re+Wkc4B3+Bzyl8G3gjof36
flinRjxcDi4cevzDqbQnOok3oi1EG/KB4sWOruaWuMhqJcJ6qu2QPjH00sbuvQISBriONDP8WQN7
8md2mI17KhGNnFzsI+3t3kwOL8QzOXy2t/2NmVVabZ80fn+9DbjcAh6WvRygAHgfyEH3noPK6kg7
PLIatIoYVpNskYwWMgykFNeB/rjVUVEl7cIcCNiCLxTTCDv4TfsTVHuMElyDj/47dbIQBHK3/DLe
wVKpgX5pycEKPnX9PuhouQNyBTpva2yOTSFiNQANm73WSlbITkR0DIOgkwSnvMUyllyQptSY21uF
4tWjCfT7FgL4Uu9wiBMNkQDgR0QJtiSqrvfjM8pfSBGU+JZc6gxh5SB+RwtzlSxZAlzOBbPTYMvY
oP+93ErQfn4Vxj8CJN1AZrrFea0gI/dhg79jbfnfY5JWuED5TRE63ZzpljuEgbxYxWNBb4vjoIhS
c2uNRMHxnxUxwMD/N2JSsE5xjVzhiDzwSGW5ecZDmQxAouDY5UPfmnCkdBeQFvVSIa/I2NvN/G8D
4NwvD27Aq06mprBBp5sUNs7PsO3icFYjzRM6ATodlI41rlDxRMsFU2P8e4spDKh4V7BmTarFemz0
TCa0IkdKdKG2g8b6Q4E7NoWWg7XIUj3I6GWDCjbbmkyXuCmh3ntzGfYvmIfrbo8ymUBtxUxwdAwb
IHZskn0khGX9WxJUPHKGXwIjoa534upOWP+zwNx6CH4kXZPV9X5yZY04mwjTio49jLB+eVDYFhst
OgduapzIdJN0c0yOcWUVSewBqCZebRGnrEOuuPW1Okf70HPKi1h9udyLJddhy/Q43zzcaW977oT9
EPxf6zRLvcfXuWym/AtrjBIClolxGKJusP4WcmKBveNzwd3p1Tl7k5UkcpC/JUJLs3ECSe40r0FE
9m9V3/9xGrNnRkvLQSMQcGdZ7t2z/sxz2YXUesX/+1wieVLpSWrUW6fyueywgK8JsiZ65oFKu2sk
GhRyyjObTaDo9CFJksqn1czpPM4qSIw50I9gobfWQFiUiQ7Ch1y15uJUeYz3QWLf4JKC+Z+RjrBM
i43inNDyZoY0FhU84scEmBhxyViFv5245dLadoER/FNvqWlgrTkR9uD0ZjrV/cgcAHPO5ZXf+Xaz
eHKHfFh8ppoV2dBtsNuYCUuoCeq9giIzc5MUWqCLUCD6DerMQpTqtbfzRh55kjXgpTSYgi0V4mxX
nntHkUlZPjxd13UJjBIJSAPgs91BDBhtz1LTgMSdhWcT4bGpzwVxGIE73JvmmV21+gH7lFvNrgay
bgTcB8z2J5PpsjDh9U3D284ItVspU2bE2DTOnoIHIrMVpltw+FvS9slwEmE1MvgCf8BLr+BHD+O0
cIK4uhc/tKe64HK1lgXzgvWHJl7Gizc0wN8RcVcrhanCGRiYM8tV8uqi1YeAVyWLSyzOWZBII+N8
oAU5KZL6R/bdJRshqb42Vh8y+WWBXlbh55vB/DE7/5tNl6I0n3C8JE34hQik3OZ2J07FkgOX0L6T
gQKj3euzRXrsfp2iWCpf9d8G152CYZeDe4mmDcskhZVtr70rC+HeQPBUi0lp2FazuwylsE719y62
yZ6X31XDs4rxh8Mg/C4ONDmTAcQ3NQDFUu3vl0lOqGIi3bish25iPmcTXUKcjFxrHLlRMsQIzhRT
h09LtZOR6prwsicCn1B14U5K79Gmo3wR+4qHbtGvqo2hq0Y0P5Cb5WQ4qFWHGUTLPvOOYD3g8/02
ZXSPfG/g1UNXS8q2NEc7qtraYngBi0iyGbuzjSnCm/rZebCWqDKgTxTA/vajkLIuLfor0nPPWhSz
3aT5ZReoubQUsHdIZ2HP8brf6E0X1T3KJUMCXN8bP0z+Pfd/nefI3HAwoUnSMnRG/K2Nfqk/9Hny
HGvl/984kNw73S6sJVWfkN/6HULPgqEA1YSgBSAe1qt5UGvd/kJDd9XiOd3V4zEQn1TaMoHz/t8U
g9wc0EHMuct7JhcFx9mL8x8z/H7DQYZMwJxO3cAu+7EqT6w+gTlGz77a1985E3DZ6DKiwKk64p+i
mH8WHEZKi8mBzAaVPu++ufEXRTEPKN1UsSv8nDr7hl84z665CSdIIxjzN1f5MR58vISdXT2A2nCw
SGRj6Hood7OZ5tA/UEbMjB5nfYMmAZtruj1R5LcSnIKDLSCKupfOG7BJ0n6/Qx507GBd10OP4eOk
NkieACJjLfdXdth863VPis9goiUBEZrinxhwThKKdKH5dP7O3xquTC1ZWOQ7aikwcqrDoGX0vDXs
k7XertHfqWlSYg0Z+rp0BFSbCWGaMjgOAah1ZsA+Vd4+5zrOoMM9/HokIkmPbgIPmvxK07OffKoZ
aakxMrPquyiLQdjEWUHD8KwJUvua3Ef8HLhPZGJ3riY5J9pk5ypSYfPKEOJcT0H1Hcu9n885fI5s
jnXduh9m/QfSlgVa1jF03WMxEePeez/0Gt0kY8B2i/lTICga6qdMhwHiP4IMSgnPmTkYOKsU55ZI
qUhfCopjbIdejSJ0lQaqeMkiBizlZ1sAfxoAcxJW9cer7sYG7W/l2HMDbKPPDu7yZg6JCK4NyQs9
ZIP+BY4yGzW0IqPhSx7cOEPXMV6sMCzNrx5gRI4tAv4XRsdVLsupOkedWQGyh+QlBjbdVOYvCyiZ
0fLZ+GuuTQY3JbNCkbxQHMXsuWgpwUVSQvxSXn18OZlvPcFFfSy5Hynjkq2hp5Z+t16Caa2a5RL2
BT8E+WymfDUUCdn9cwHvt3UCmsgS/+awY39TL5bwhUeFiHgZAFjjQrSYirTVriHMDLDiccPmfMyu
x/Q4+tKr+JXxh2fflrfhEtjv/T3d8WArzy1KlP1z9+ZXkSzmEdsBh4+7u7z1/CSy3EKRciQL1HkY
35K/lx3o2KgJFkLf3JQAxMqC77G4xSf3T7/Tgcp+jgkCaxVYKyIZCixoqWpTUhoIkG4J3pY7Yw2k
oNLHkuiXY+xJ/wDT8EEJF9ftoerypn02mbHrCfTVSMDQD/pWrdQp5B81bBsjD89Ul1vxT669qoqp
VzxwtjP2fgYM33vvQMe+/TbtUv9+UIVF/kWz+s26dksiH4RjQmqQ9LwtsMojb5NNMMzDN21rk1fy
qoNNf/gA5hMTblUAIPkmAl1GDXFkctPDVCUdH8snC+91W2RYw9sLUr04m4uhSyR5YslhGXYMLsN5
3n70BinJQJ7cZC+fZdNE/P8onGYL9YP0l6sdjfhQsVokvtcqAvRgFQjIXNz/hIGzNGwZbLCTUWz8
93uK8nnLC/oyRWagoGRe9cU4mTeMMicu+rEyY0ha3sHR1PJoPiEd9HzM6+tMoX93LHHjE9H3Hy9o
E00XmMUsGXOybW7eUX+B88aWeW8UbpI5/VJgTaseibZCaEhcyaQFT3I0q5TXZEBvL/9OvQg/LI4R
1uhnchHtllzo0lw0ygA7+s5gkL/M331mLKPpR9d1XgiOKYdO9WjLN4PIsIhlL/AFxZeDLkUUtVFt
8ZAnGx6hETzEYnIHUbwH6+7HhQZssjmxNKI6dRVRtYkBIznRzgUVSu3AJNUHP2v8jJFsayhjXG9g
bhsFDBWjJbFb3vQlyhC8sLjfe7RidU+ISs22ZPnOkcNd6l9L4caTmQnJ6s0uqsekks5+3cMSOYfU
bcXanPU6cIqPIYZECgogf9ycK9nuU4eVmQjVfbJiYPboAglVSVwV+tHUTB/OWS8QmmzAyGNirfJe
CYtX+p/b2fAor3AHbBuKNU7Pbxc7Onn4g77fnvjIc0UNUp/uF/hrIpO86Og78+XLE44X33dzviEz
gE+LpCXB6P+7hHd1F21ZaJdEnxgQUXMVfpIZv2kW7yPLwkJRTz2PcLgaa23VFsvK90Db3L6dygW8
2K+abHME4KjYsEXd9lfsH/xwKZ2ctpzdZR2cUjTe0qHwqS4BFSLAnSMr8ld3W1AvHR506V+KqkJ/
TdQK2tv0Y0LAJQaRZZlhbEH8FpJBjxj4boWxzB0IVJfB+OB2i6XG6XZmof/i+z6K2nSlCBJAL2XV
a8EvNs5DMltGhJJG35Y0+U21MCBpNqtKXIrf78ApVp7aknCSeiOowz2/h9GRBnsnP/NzCgKfJ+A6
uvj5l57I0mXcYC4XnYvqubS41/m7LzuPZcJisdqdNSUU6qEqYsZT0edTzJu02G0u3kUF6O0Su+Ei
nauT6aCddFx5rJnrADZ9JpH+5ut+BItTsISLiIVRgmHduuUKduj/uyPq5avGyNeR3tFBt0dnRUb+
mW+oWPWN54TVU9l6O4n/PiUteeO1r7lxnsWGLTEDj99qtc4CLjQ+qS3wY/B3fhuZfMLuUebUnLTV
GOm0qfIvTc6g6nJx/bLgg+H1zxmEDeoIlF8oMY0YGc1tkzmdD5PXNIKq8QgvJrV4ps8rlZg0ao8V
YkfOytKTsRPFMP1NZaYWni67bX61/wn/CK8dc3IS8uKuaVa57S7txTbz/Bo7lhzaNn+JqxIh10+d
ODJKKByYyuZDJSUBNQrZAiGgWbtKP5n0uY0aYhfaF4kg5kCBjpKEPsIN47xaz/nLtN9qGj9lmGAP
dxA+YK7z8b4cLaNopxTmd+6B9yqNegAJ64cZCiMYcoM7RUvKyA4JTo0L79GwLQy1OMhiCSkae4QR
wX9507rqwXs1uoznz0pWlJZKrc2eWGo63bmXSft5iEyiNVPfItU5NUjESxoI3AwKaoLeu6aKwNix
H+aa+o1gyAkg0moN8/sqINdDHzLdJSli5ljRDjyF7JCF5H5pIxpEihki8KfjVt5vcoKRZryipAOw
e1tdeI1WEJ1tJCPmskkaBW7BZcclHaOPLdF4a5jj/D3ietgo47jXTSSD7o7vd2gpNapmvKdwCmX7
VqY5kH+/B0eRX9BZw8pJu/DojchQ1gtp2rXyZkecZodhD372Nej+v3Znlo2rTbZ4kE6xZhnmro6u
ADxYmg2l/hVLOfcM6bAoJxEetamzCDz8CnQ0jsrkNRojb1fKp56lM7cwS3nhSYFrSUROAyrT84NJ
nEFUyC6GVLLJXjAl+Z2gO9tUjsVUg+reJ2UCv65czpaU5rru6giDSK0XxO+GEFOj3Z6Rf7A4TGb7
nOL9W1/kGdAkxl0STQmkybnmuO9vf6jO+BifVOvFMYk7JfOZTcLDT9dkPAW7CjGSER/K5dPLwZRI
NGFArd6UeD4p4BldqatY+LMgw/eYL4JPHyxPhUBFS7gFToRy4oYKqNpKpNQSThg0g16QaqQ1E0L+
o30cs3P2S4+PsmSeOgEn/5WjrzGt2LOEiGc7brswhnsZEl3zcwITBxLqYgNo8NJg+2rz6GHC9GDk
QeCKwwBEy9+j2sGK7jiiK4IaJ5R6OJkA4sHR0rm1jV/n29zSbatFz5PnHkRTLnWFIJwGW4BdgV5Z
bla1KbzEXe4fVGuYxZUF7RFS5NKu367vnMrIeX+loRyW2yAS4EA2/FxYmraTdl5p2BB09EEZ0ldR
ecvK3jD8vF309wpbvJrjUiugd6NYHg6rm/IEspTdLwWx5Yph1soSBRUzv/5UetPewj4fGI3u4Uyx
YKprEpHMxgAW6dYVE5uqiTfuULwP5Opz75KDu6niJ85NoAsO2nOIp1BYraRyrrCVjIcDJJ8lDaeD
U+4X0Z7PYqYqTGdoSczeKo5IIUVJ6/9RODSW3ev3lg/K0aOKl82VH5Mpr5ZX+UXyCI8EEXgWINGG
NSwYHllTwLm81CAiJHyBxo+UIrxeBWgVeVI5AHINlT0jfwdbrWjpo+wyo2mC7eJ+Bpaqyi90UY7F
JcrQvZBuxGXy5ntthYRxzCN5h/Hinq9L8l90jqMfQ3DpRHMPwV/GzViA4W/fYaXWQJa8jwMXLS7K
wt/J++VbsfwnEkOtsLWtAlPa5ntIIjm4TvoukRVczRULSsgJdy4ubo+AG3jjFO1qXluGAZichkY1
0G6W0eEmxtz1rs7MfupEbYe4lYGNWwIbjjL7CtPq1YQj5e/OTJKrFtPYpmf8gW1L2pNo1C7ukmnf
mXKmm2rGFHVSmGHJtOZK7H+uwSWY7wZRlzeVP8lPfja00gOMKOHZZQy3DLSPpA3ypnjpcs2UVJ4F
Ip3AXhIydesmPIll00LoNJ0C6iwG1htdJPhB1JmvYi0e1xV2m7g9OUmyBd1Hcr7xlCcYHbKPE0BF
N3qLJiGjy9mI2kRLaTbZb13HhcYlJ3dxMxiwKW793lPkQA50puloJYiosby1Qg8xxBpVlUbb3Baj
Bc0uPU5iV8GuHssOZIcfIZAggbuDzItRuok5sADdzQqVneAgwwWJPgE6o4z0PZYWdOD9sMCakqcG
x1mE61xUN8JLMhEfBE/WsazSCuAbbeog7SI/h4IcPFR96f4PqruiabRHkYf1+Y4ApsAPPEVM8BX3
IgKQVE95pqAXzj2WFWSgtofNmhiwzG4DCYiQxL9lWtfX3yDDxXu/dPbVnv1yaj2xs2/Gq27vodXN
KSmgWN+bewzPcflloWWnPA55XGe7VTNNfPWEQgdLlfVg+wN2eOIZ9AWzszetrtDzj7QRZlboayp9
z9Oyya3qqVZlGhNqHUNrt/bDs8riOWqPJp0wvnniupecx8XP8hjuD3yHY63nXeZyNksKfKzNOtcx
K1oJbIAOSd0rFR0m7Ki7kJAsI+LDGG5/5TDEX0MfWdxYs7f6XbRU5BQITxiBfXqLy0SWb681B0cG
i8mFr1FLnx7HsulXN5R/TvYPL/zaDjmCNAfXOfxmrLiAX3qceCU09yRbyAUBpNzTaNJ+mRE3HALi
iVhWS6LvS2Ab66Xzw3pWFSzXRM+SXATF+BfgXnmc7yryExeBYcItDuwG8AVvK+y62sAgxmQWoGyb
YbfSJ41JP/yzLlFOYxHkEQvfRkZz4fTdOzWPj2HFv376puumYy9QEtoUJWA898qWoF3I1ujf4IbD
BmPy5GqAcKzIFq4F7aroVreT0qhgD30RBF6PgcNBohVJF+2htOfxQMjsN4d1j35W1lMW3W1mflLh
tWd6CgowdkrUGWPZsk9/ywpsSUx3ir8HJHQWkMGniJ4zxcxuU7hd6FNx7CeWE8zCgFUnaYEnL08/
Tn1D13G65mt+lOLyYtbcDG5Gh+AuG4GNMZlQmThvU/nxaAjknR7/5TYIVsrId3eDUSSbKSWTs3Kx
PJqZxi8ny9mTWX/1kHqC8wgcQwWJPKVyJo21YGRAmFO5ANWVcH9EKkeUyyejyzAZ2AXcAp133zhe
mGkVmujEgZtgrkkKpROhpGSHauxd46GcFdG4O0xWymAfFiEoF1Qm53WQo6BI9CyzzW4PEdzQYk2y
/dpKggcgcOHOY2me3gfWKyuPuk2apG+jPP5S5D7go8JtmbuOtXf0sXO1n7sSJSBYD9Z+5OnDGgTy
g0VI4oVc3eDO5iMZ+rV5dBnbtWzLMZyH5/EW46ab94/E3myg+DqRQFcPJ/6pU6kp6xWcMRp2rJFi
fCod8WEcPyt1CXqZi9fBl7nAdWG2ZAU63Cw1ULSBkunmTexs+3WbvaKANYZ9WekICBIWZQivFHv6
DJkyWL5b2qhMQAlAvbv+vgSdzFWyGPlUFrtpONH3wYoIraaEOQ1XBkZROBBBQuy+aHyuBtZ+qnZU
yKTxEUCuF+lE2TBLmFG0z5SWL7YPrtvFkiHXiCBNUmAmsI2pHloQ5RCL5tulFqoaO/gKWbSORmDY
PVnqQIGZmSdqSHncAA/spu7fmA5C22ImxG9qfE6kdRdfRduHVmTN+i9oCQxS87oHaf7IsTfS1UXN
IYx4h8nef3t/8ELKPy9HlHSz5E3ShbWb1X7c3/jD8/XQ8tb2GQlOKxX1ZH/lGpQqOdYfP+n9ZMQx
k1MFotWiThif5pBeMG6pa3u6IeV2T2iRPQqk4MafSr7KDYHCqza6yEQxchsz7rTCESF1nglvjn+D
R1WADV91R2uz3KTqzL+438WvCddVdLvUfFL3dKH0mqo6DfUv6rE7EDaeElkEvuRSG2gdb5tQZyeF
Fa0o5d2ruyB5Vg0XMb6eDB5BceMS8kyhb87iJl2KkGoLqFB5Sia4eq7+rCE9QrPf++yCIp/BfLrv
xAqjN53j6e5PZoo58bgmj6oQb6DhIXZQ7RFmFqHvBxO7JagDZSdEpOY6D2njn6brRrldmBEujXtK
Wzs9CU2y7e02UZvhLONVC0Pz6ZL6Ym+l2ipTQPLxTImg8PXCE+Kajcq0SAi4LOeUaJkYWmwP5cNB
k4hyaLpIhvmi5NfDfLbQ2GKaXXW17548WzpnKRUmLKB/qxP9pGJ0KC5TgQ3/Zy0A631bDeFEtSmQ
jknhZdeSSCCdZK20QYD3QwrCnigHnQiLO+qqYIPCgKdp9o1MlQ2xCfWk8auUKL7qadKodxD4ujfe
+5bLcvjSWeUJoZZ688udSt4ge3rB+YU2vWtf4hm/CdcjyINT9UxG/60TmSGsG7wdawURIGC/PoUM
2k5y1/4Flmta7BGyn/l24GWiSTejlBl31nXYUkkVg5dprbt7LvqUpZtzfr4zW+qqzhKAkuORmoOx
4mEksK/61WfcXQgI9ZRHJcnN8krbNS6w+mRr6qsOLu6bb74FVA/w+mjb6On8NKKx1rmeA3SaXYTm
R+s/u2OR2opJDpDCPOf3/VkqEhL/2yuD5iUCviG5Qei8TroGytwfqlXC6KYIpvscwxVggmHZhoxy
Ah7Tz6S4+f5MmUkKTFWoHlaTqZKxsdIGWLnaGPQdbSObaunvNv4xOtMahSLQU35QuD2VI8gwKX2e
78skO8amEzvNg+UtF070bkO3Zo+utC7qaYxp1MbO5xwchYLw7vqCxz4F0VbI2bD26lHSQUZUgC+d
/RAKqL5H+R7hdjxabnXpwp5e1HINpl6JDgr5I2l6jTEtpbQzR1H11mpS1zNC08x09t6W3nNHYuQ8
a3DkYxNgocu0Ytp6h2ka3lEzVaWpBf4enaatZCHHdwIGGctrKEJPVZi/nXBTYm656ite0U53kj24
iclMa/hDJXOmjug7MZ9Qvp/ojl7FoO6pT+HXzE4uJ/Cpnn9gXDlFsgBMXAj0VTvsM2yyMC0Wx9cW
1lgpT5Tw/9ykZYTGH4NazM58B8p+K95O2C/e7MDOm9u6oNaoUMkIkZDoTnKMRMqyrnwVpxIJV2AU
KOqQFDyplFHCuI6eeFI/izqeQRL3081kYTODhP68Fl12Z/GJXcV5c+2GUik+PlKOiQ2l5r4lBEdZ
oLcy6izGmTthNOB6NTYWcVjG/cxIGETGJj80ju8D8+zgQtn5iSUG3pnDSBKUbJ4VUVEtExow9GbB
BjFFfee4HUhI3Aq0sLTIFR21BpJ2XukMs0abdgOVWl5JLMIhAGGpgZHjI+RWtpjnwW8m07mhIe3U
mEGP64F0bACkEMBy6oPDINKpHriz9gHdNGiVdZnZiCDSXFwOtRZwRhrPRuXc4zkcFF4NqiXau/kk
KlB4UbooCxBtXQj0MIIi0+U/hrHpRtXKddgKsJkGoX3i4JjB4I9cFd8SxqFa1jw3Uxm9l8Gva6lD
dvnqa2WR1LxkFDwBjGnSZaDhIyFxpXkJzzUX11yULhIE2//0HbfdaFS/KHoO8qoTJjQWNzPUroSs
Q4gqI4jRvs1eSJUEjGjRxZ25NXyXOQnNDqme4Z9ptqiKz8zbSY2IGJtQaLwJxe6S0ImLT6DKmeMU
luimqmhgxOd499454rdOtTgo8ZDVM/iucNkQFjMTbdmMHG4bLen9kZoDL57IyrzLLnfmeWUGa16x
WKOIogJvS6PLvV7RXu3TzLaAO27U0eL97H4cldLaXXmFwc4PUUjQS2D88AYQV6u22ozEpEq5TYih
hTlyc3vUD4XGOiI8uAYlrrMhIyrYEIrF4xMJu2x67aySkJ1GRnGY8Swm4Nc+KyCTFjAyROo6BQsb
SB0e/eILFqinMtcKRRc9jKgxz5sQwIvabooVfBK5MHOEBhcJyz4VBdWPU3xQ3LlA+7tYPjyZrF1Q
pGm0zE6XkNX/Pb//VMrOfZjfPogvx1w2WH8FpDGek8z1GdFFp4EKVa7IgR8OU15ImUVzsOoqkW2j
VJslxKaRi2GbrQYBMX/zfaDdwxzhwr8h+qlH+gVGMTxezAtMpIuEFl2LZEMhdD/gLplS+au6osqF
Gdd6A7/lHEmt9iFNu+b/rPHTwPJkAzBatbZKRQZ3WZBj9bcx2XRIUAlPFgrc1JtlzfaMllAZwN++
pKdL2RF5CTl1QhwypEPOMHOWU1lqQb9lc/F6zmiBvMizaekARGz8C5dYxwDMgDzhhKY4jbfukPXu
/kuvrRxFTFKaYMO7er57IkgFyWxpsOc/YUBztToZOijcD5cJFRiBB9sCS6phqPrMAW9B3wrLmREA
V2R6wnPL/NmSmsZLiPcYdyYK7hbU/9+mb924vQkYVaUWaMHm6CnXQMoGTmopllt5ITGdAnLmqIzQ
NZbEUi0IQdIuSod/8c7g1Hue2tX5RAbzR7MUGm4NuJhB9EmqbDN0WeC22hL6qciEB8/ee3VC/IZz
BVUBpyGxK22jXfLMg7OIJBUyvEyURRdB7D5WvVW4ePfveyDJz1zjBQ3oFIeEpEHhdAwqE80xrB4X
IEoKFFJ4DaC+WZcwrXCr2Rbw2Ft7O1W2jsQ0yzT2DBxt46pTVjqvMf/RfnH9rBLNsFv9Iq8WrGv1
vxYeYeYoGpxFFObEmERdyJWvKAZt/Czam5q29YqBXaDm5hFkMfFy8BFHB6vRRRkBIyngIT0PIccm
aYSJ4rljefIliGH7VgFNXnt9G1jzgWrqtciCt12Xj3jAdFkRlWuMU0wx1h9vmZttk6UxvtOxREen
h4AxK7MniDkPK5U44j68GTOBhiymidp6iltXij/KNDUgEB/erV0vl79+zcXGVR6CcJUmCMaAuAT5
rr2OXwDHsy5GwN4AUxNsMW9EdrO/rhpfQB8jFI1jn6XRLxPvR8FLk89R3kPnTv9TIKTbqYLN85KJ
HpYzzIBOBlXcJMA+eoBo1CBZ17dRkZxYcJzQy9lMqV1s7ozi9cSyeECn1PdP6LPCTS+eB0G9G1uZ
RPlgd05mz8/IOkOEZvU5gPtx1AZGh48UBeLndbch7yZNtNbJBfx1gtbLGFZRfskOlM7hbv0BC7P2
7LfaOnbhmH9/L+jNEfjU4xg0PtQUz4pQc54vLcnhy3OuC42WNbbZvnKBygfSLbS0sGqi5DYldT2O
shXUwNfMRjmAsQU2K1o+qiWO4YIZlEoZnEcj2hm/zJ5VVktW/Rg5XpNVNGKX89dXt1ZP04lVaOHV
hUBSJnaTQ51XFoRQPCrxOzB/dlAddf37XIKJuFXHJmepa3YK5ajK7gL/tG7ecFeZ8IdDbabw06+r
NwEvY5mNdBgQnWXHDpVAACh4wsJCH42bIRX1jTS4qg2K6nxlXiM4n08GPd2Y4WZTJWWYulKrUUJ9
CJyMteAnLEqcZmFuTFkdQJjd8QHmijiPs0xsa3u3NjpWx7LxLMgn+Ec24uGSDX7r+/oBzqpup0RT
Td7Mixh4lDPLl0kPGTNZ6pZZI2Buccumm3jstjB4j/0uJeSvQhWpIQtiHAnvBmVojA+aDKQ6cktp
OA09Do1IV6bLw9DQOv5rVww+nNJn2Tu54mveMG6MLo/sEGbWpcmRlyjDRsr88YvdhEGxczAVuvU2
W2peQHcXI+XJtO9/f1Tsn0GGCl/bvF7xfuVakxYP2dvI6sm/egDsctVqQhNTwxng1gUG5guiiMXv
0c+asQLcgu6FJ+mQkjmP+s2dPiOl1Nr0X3cQbY5cnKiARcYADCeRtcCYRMefArFyht464uP5JyEr
Pz++8Vo007lAV3VhkHdsf05p0Qx5yKvz5/A19AwGGQlbnB5BJreraRAOIzVH2fK8Rvv/eTX/71dJ
veOlU16zxKqDfBBQHViLoGosNryAfp7wEAWtf8dePNNKUzx2yKIKyFmrNf/XOVTcrFxPq9qFYn/Y
PS71/stdy6zYaupbr5l4cK5uNZ15LFdscYOPkXZb2wsvIRRMa1JqN8U+cQPsiufzMGbjcZLLpu3T
BwErOG5Vyawmxlj/D961bDBpY2jbDaZ1+TcgoQDpW9k6WN5YOJKAALEAKWnZvltx4JZHsnuL3jSj
nYw4pXAOP6TOROn7giNQTUF6JFWUV6UB7hFzYatB+VlcchqagF2ZprNC/vUC+5KVq5BZU4vCMrSQ
UYS0WDhOv+ZENPzEXMQDsw9KxrRvekiQEI8+P0rO7bqs/630wlyl8eeEIpU4lbKz8TVHy0CwEtnO
Zx26KmeInO8P7ZxlB/eSSdXhe30+nnoF3mE0t/khx5px7BES0CkeYRl1/fTuppIZNefaVEvQ4qci
KuCnXAV20fvWA+wMrtFsh0ngX04vZqHlDbBQwas4y4I0oukXRef645aoc9KtWzq/olipj7uCWt95
YALLFbkT8y69DX/kL3l9XmQJ6WOHLhzeD04O/q8kuVSYUZK6Os5I2CvkMznAIg9P7U258rMX+sUa
k4HMwQXB/nncF1Wc3J+88IiCKb430Q+5Hdk2yOzDwHU/t137hnE6PVEngpGRXgnRhjgAJIvEgBdr
U/6fsWXDNl8aNGXcWBOYiU6mgtxYXAifZTfKVyHfD8L64leCrrohTSOnUnaAIH7ylHj1CnlR2psj
XqZ0p6fyhXmbVVVjrDxYdFqW+pJoMDFkHvvjYohAz+c5hiJ36zxIenT2+dX6TCfWsuJIFqsLcbkT
r0Hl1kiOon+9pRs+UYSFbJPr8b1ctC6zKb8b3hlOkJ2Gcl2tLNGspR+Wtc0vgnRMFlF6wth7me49
W+qRKflQsYDBLeVlghESZ44Uv4tX7+8OM0DcLGXsD63VMoH1Yc0NWuiNqM77d45DUGBnbT2HrFqA
oaECcgW8PodbyqbJ6cx3GIKx3/4R+bDKzNpJ8COPfpRJ9dovk7nsylkVbVPqf39deGp+fGph9bJf
ezpOI3fadkcXeMHKTZ939fFITWBCHxgxWhpgwlLpGqCmIvm6kYXHbHAdc7yJUFJnjRH9Bqr0m0Hf
z6yW1IERPpfrLWcMHaYiQRuKgg5NxPjovTY4ZYt9G8u8dY6iymX4sk/m2AXjjbzuWKJGgS0gBFXw
WmDHAvAdGW7pIuHc7Uc+QXUg/V/XfmOXvs3pCw/3pNbU/CGVZni0JQF3jl22xdvN/BIsxVaozcAE
kbiFQmD7RzbmxHHnBeFnN+N1mU6nyAtkR/UWeD8OznqiJUiCaP+XKcumOi49e9+fTLNRpxF60oAE
0nDu5xVAW3YphrB4gCWJbgUZ0DmlRxk05dBcPOAojcBSOxEtM4gw0lRBMW1vMb2QjuDoY+JnZQKu
fZngbqtzNx7fSH5FRKmVX2VH9lg082hkUUKoaADOXGj3AW20C+KDTRbXx2dpXsER9eI0f/LtpVry
WG0NpZ2V+kB2GfbafCZUynq2KKML2qMvffHFqiZtL+H4ZifcsVUHi+Ic1UPeZFVp/EPPyDf8QpJ7
2beACb9FZJQL4ublCyI9jSarFOTeuQnY9pEyvlI7WYo4kRnquNuG5DRonQulaNIF/T532+GOelf5
SoxnK7M4/rvCjantxcXOGueBt7VLH5D9cTA6DEp3MsPy0ThtUdJfSgDuLHshyLAUs6WGxyIVXv5k
eY6xUhFqJD12WT8ktnzM0gP1uToJYbHKVAN7xUIYJ2NsqSbY6KmX1bt/Y0OtYvTh20Kl57oQ2W3v
AW7FALgJiQemBuWzvokla6BBwmCs9Sgjk58OhOSrkYOgzu7gCI7qAPu4Kww93/aRJ3m0cZGi+Nhp
qyqbgvP4+xbakH5AJTqxtrjizIImR+VdJ00JzZJ4RaNHT/6GLS0APIa5kL5H1TgfPFpKQQ1q3M8P
/GmdoTGIakWFnV4RZLBXoBCozagyiSBpQgMrJkmL5KMUOOrnG7otbnNDp9GH2R5BNhmLWYhKlyd8
ShODbYs07KYOQkdzN0Z9sgwzrh6tM0b4fR4Edi/WSqNgLGXq5/c4ytZtEnHRxzwwwu+VnISnG+UA
jXK6lKOJu0GuoXxSzeLCC10tIE2lSKq12uov70RPjYRUDNNkQBLawIc9fRJ8HGNjKLwksVRBnkCy
AjkLKStUJZL0qpfp6esBH1PXsQLy2IdX8e3IFi8S2VVwCFegdAF7nIkDAPjdD0vlXp20juK5JC3n
od0zpEh7cJvDUa00Nin/E5PninxdgaiFoiyLay7M0pneqxZGfxhffnhWghQCpF5BQoyOo8SH3a9X
19aX8Q0aFPlt4bcnh8nbqSrKc0HSPZ0nKvw7mCmCVlx8dnO/ZOIXZkvHNrl9Od7OVhE5mfezHYY9
TFuUGS2VO6sHccJPsb3FEwb/iNYilsFUSrm8sFlv8PBxeG9WW33pMCjT97EPXq1m3FmbekXABiRv
1GA9tdxZzjcnHE1WEFPTUUIX0bkNvRtYBUbEabyzee4QfRbO5cTr20TvwHXyV5+bg35IU0kJLJTz
JyxFTT2r5RSLqRhFcIZmE6GtI6JyJpYyT+zJ0cuNei4gB7O8pzl2yvf8l1OgPpmTAVdRwbJgiifN
+B8CPxI6GbIyZcC/NoAUmQmwKvxFvq7CVjV7qXKHsqSrsIwwZoFP/Kq+wObBo6ruYX8oT1+lDWxb
akgTvt8cROoc8oQrfkO+Lk00AdnvKqpq1svPx5PsueOiiluTtcqMmbrKyp08ZDey35XINZkaedKw
ylZQf6spBPJgFIVfljadF/fknVqJjnWC/Q/v0PR1+jvJQYJ+oLZU73BLw/BEKgnsuseBiXD+S9Ov
5whUZE+Ou6oeJAnIVcHFtiXCNn5bzEziZc3FHPwkpsHo1wg5A3sesv48/C+QbWHGg7r8vkp0fqqH
JaCLipc1rC2YJda3FQM5D15rtiHPZsEs0xUPt14z3RzwFUDa8XboWx8FRMlrnULmlVfZ0rj1J9kT
SzddUovr+CSY6O27UwKE2ko1kp35Fq75S5QCr4NoUh/CCQe368bhoXUxRuy1zaUMQNQ06hvu941Y
HByaL3+rt1An67QxFgWVBhgmXl37gVaE+P7UKdgoKyrDXGxxAiODn3mR6KTZopkqTI36gwAWCycc
8MlyOANyRv62Kglw/C7wRCs0FBHJsP+QGVEfDyTnNqt6dWAGtxkdc4tKOv3+4tSXAvP/0WhB0vtX
9dKm2FHuB7GujeRXgq9WWgWMh+BX4VXzYI6JhzoocJr8iWfeOTkmbNwX3KO6W71Kcu6MsKG+N9sz
E8R0uyLwelIfzCLknfghF25KcRFM099YVsBw3Zzp1uJh8IXlanptJUAUFiA8Qu4MiQvXA3f3ljPT
gbf1+pseH92C+ncKGmzv6DaVQXPcU8V/TYa9vlQq2+KZGL06s2sF1ovJIVYP7ipvO1PDt0OkaABg
SYJtD+vyNu0zqs+l5Q7q8CPOjNTGZCGJAbxJ/SbLAkJ+ZnxovUZMJ+Y+uwkQe5UZBvW8bVCaGMmw
o356RL33OACSVo7o4k6O4nDiWwI4oiPETgHdBbR0n7befpiYvHEAnUdQ1mNgH3MCJknYz0nrJVYI
SoErCZ3LyrGQgJv7dLzAcRxYtgF1N09ks3Svsz8yKulRCf4kIELsnL63dSfTbEYNWKvScYn4zeD/
6hOHsWxXvhQaOeuM/SZhi19EmZdtsKOx+RDQryAQKp/EtFlWEv8HbCfh9eduXtUlRdlVkpzkIzaF
B4eehycaTg87s5YrO2lmVVldIq5I6qSJsQd9WJ/qHgpriacAZ4iAweQewWsf2wFSqCq0EwdBUpS7
bHD5BxILQY7kyaZYrqugsoiMKLg6Ml0PHs4E8tacpqbzRz+c9bRGCQJb3J2P1OIm8BwHawJ50icR
SHlGlYh1IA1ApMKbuLQs2YRxbRhwF411d7ndEiMwU0IGfLAnx7s5v4rOh1Dwlk+PBaJ7AcXuPgeC
x5c+oN+MZdnpd+76K25kunTlSbqbQBhZZmBOtx6UDRn4GDVFkaxM1md4wnTO5C6zt56EJvfKr1Nn
XS6iRY5uHQu3KdlampwWshsETaKVaqnDUtkqBYLemb+QNiybMJ8QytURe+0ZQiPlC+wWncfnE2IA
W2g2crEzPYkfBzBBeNYDVn6UJFxV9WoF4JcIUwlad1XxFhhg/NViqFbVuicDQGzxoxmAX5IGkefK
2xXoga5eUweV/1LN3UAz1lopSvW1pgvpPTlfN+z4RhVVdp88+lQ6OjATaw1D6qdurdYePqKpOV6F
WRDOVqMgZYBL0pnah3a5kTR4w8l0K958jdI1qNJvV9zy3H7LGTal5izyDb+L8O4Q2mltLJ+0umMO
LBV090NMCEEnArcGHVdIsbRvo+cnZj/WISUKpoULeydMjkICACT4hRotkigikXMlnRb+arPlqqiR
5vMYncBh//Lcsvb4XdonVIL58qK9oC+FONtx/Wk3TL5JNySksFu1i0kpVNZh1PAXz603+pdzUybI
YHT+TyLaUo4f5BLTF4bossAl/EWcYYxYUtVi1yEP10DtfPU6V6ssvRHJw5quxyExExorRRO0hENv
nIgzFGVt1EpSbnbcEfyPs9jRcHs1aM4pgiumWAuqYEAs+8NmgJPHCtlssNyh0EWL+chQbt7oN+DG
NJS/BmjMErkiPAXGRgxH0bWoK4vWpD2LFoae9Hbuw6UiiDRAHviASGO2jAi0LAIQ784JaXl+lRG8
kU7KJ9XBJHQPHwMUhIIHGesioM7qwiO2fG4L4EndVpsBlK3YIftHYlTXU8ZL3KH3Jbd+dFrUaYkF
KpmNa15t951NUKQL45RJbjZ4wS9kxMQzRy3t6isuCu2FFoyoFD1wBzU/fpoCo8MnZPOEjz1D+WHI
kSMzOxkatQJh7MsP/7iopR9a3M0taPqeB9nHwyWHuB8fflyKb5Kt3WTXbMHgrGIV5a5IFv6HknwD
S9mE+v4Jhca6FKKhGGV9MXtusDYMs21IqH0v3M+pi85HzmmFSPNIcnuWer0OZf/2VjjVxu1F/eCJ
3uBxq8LlPuUe3brlE5nNvqQ69vHFleSQ3WTpg+7Z8fwtziQGdUzSwBrYKqBdFh5qoUtoyYnJIeBB
Xe3BVKDlEvw/bw2elgVl62hVZeBq2Lqku01F1u73cb2tCyu1JIRsL5UcvTaaqgBPqqPiRMYABZQb
sadDaDp2FiKnPTJ4JHawspNkuTr5nwpMAxBNZ/GtS91KhYVq226TG5/v6S9UplWVgg0hdAt41O0u
8RjpUHzQvj3H67uOXFUAEyT5a8SuudYX+vmlsU40vgXnfmobBJzqF1DHVyzQYwcLTMUbg2ARJGwb
xRfymFzNUs/zII2M/uEOnikswj6OpIk4m2hp33P59RVMFMNlNF0sK51XBUJ6PCxbzMLWzR46gtZo
7gcKnhdF4QltIKJ6T+Zpl/b/m8+VDLEbx8vXqY4xNvU98VQfoDR693AohT1+yNlPdquCn0nFWceK
dM5TSy59ik8C7uCj+M6IzH38GLidE782CoGfe3iQRJEoUdROD2iyKveU/Cu6K+Zt16hDH4NW0oBC
FCFR2oJSeRmenpDYDD3bRbo4KYM2QaZLhoufMIbDiHdCzZ+wuGmxW2TJMPzJcjdcFFQTMEEfRsph
HNiJqIV8irAg6TE2lqYtAw/71zfll1/7NeD004XasHjKyHsQpXONzKF0ViGBqyS4evmedPwQRitg
r2FkGDoSxdbvs7e/9ruzxsz9rRbVFDttK/P7JuezCQRYwKkyDsNpz1wQ0KIlPyuK4BANSS1YWfXC
9Vn/Vd45aMVOaPKVcxE0knkuJlGcZoZxk+bswLdQBcKCygQ8nwSwuL1ooa4Y/Ue2p+bThr89XdY8
ydIL+HluhVn6gm0it/3YWWzOce3gBegBPNwY+9rlRZfnHl+e/MF+egYATGhbaaKoQHg5qN8+Avh7
w5WyC6TJudrUrzgSAT/5D8m8pocn0WSMclR4/0EKE8ylkaWNGTeGutoTjtOQaKJw+TA0TIVaxBcw
R6KXW8+ZLrpam3dXLbC8Ph06jEzt3eSmE9M0c/ulMq/i4bbrJJ/w0DQG45u1ONtsO7YNHVv0gjDu
ih/nU4Z42pgxO9cxH4NW3rprHxINoiSimgu4yTO+MidDH+Se5Wa1GxnZ0gqneOfa7ruZVrtwg/uZ
wRYvTiLQHnY1apRiNKoSUynZ//XBj9l36t5bgEV6hD199Q1ZNAyQq/i31GxAOIStX9qew5+r8yXM
C7N+T4vXOLyEE9JLZ0y5V/2AVl2MOIID0D9btFesL9b1dBiF42J3YUDu+xTEsbAkHr8oe9FyWfzR
8nNziLRY5gfbNkiw3s9EinYOEW173zzHORGvU3b3ajF2rL289SKWSOfcZeWRJ6shRisnBsywmouJ
2BfrDnfEoxxFdmV4Zv8wQpSJ8SNgaWLfe+KPIemPeiyCnezgnM9O3EYYxWMtVllooRbio43AxsFL
d4Y257LnRuVS8AVDEnsL2QqXkm2mforGLg0O/gvN0iK4QbZwVMOk4yWtgi2ml4C+D9QU7BcKMoK4
932wlCXfWm3o6u0KjhgyB9xyU922+e5VL3e+5AoKWEgqgtrEOWMDTLKEnXpNmIsc98+d+CsnL/Tr
GChL2S71wiDUGlNNwcozy3JDqLizr3EopP3obwUDHzh9M+7epO6Uy0fz/oULTrCOI+YiOXXkJ/y4
gafCHYCm5J8xkV7NFxK3OMny7q4sdcJLSsxNxlDHGw47wS2AOQhGblf9bU2MR0FkBMZVQjgzh2cG
8h3a5oEK/2etTFmp1Ff1EneL4pqVwe3wAMq0PcDEaYd35e2nurSyVeRdhQjTw0cYbRP6Xpobx8I/
UL0RU+awbMeFMl9SNICACY6pP4g87eebY0/YOjvaVdP7adVmNkvaDMqwFFy4vhEBhSV9WyrDac3X
Nezx8ypQQggxxrEXf+aaUkDvdlhE76YYwkmwCRu995aYhQizGkblzYvQtSx2CBKRJ6uAkfScSNVp
1cMQhBsBPPkO3swvfiDpXaldJffxy9gObaJseVzCnGVwOzHsWIojh3nrh1My5IFhQGcd8jc87bxX
TTxgrBLZAWanUoH696FEACgVXPVGe86kM5dno9AzozqNN5LeZ70aG6tSuj50WTbjwYCgR2UqgAbx
Fgo1Dlm/UufjvEmjj0hHqfTm7IYsPXbp7nJNGJD3BowGt5Pgd8mQjtiPdJI+vgVvBrFmhgnSfceu
MlPPrfuYlC5/pR5ZEqvCIIsfKo3/xvnPNDADfGaWOx/0sPWpiuViEq0/9wiJhWpPwcNNNtrWFn1n
xQrqKhXjk6XhuWdp3KiieI/hacDPzksk/DmMtTkTeVqfoRSHMvjE4pDFXrj0zEeJ3iZQ/TYI6MA/
KooBu6vo4QBU87440O4GKcAkWTiDDO4qSOCV76djqrG7EbhSiFZMerYgyQdK0CXqmIdRham+Bmln
9Qx7hyMhbn4DPlVAWhBJ9mGeyXVsO5ZtSyaSrgIDk93ErJtNXS33tq8KsX3fMVV/4nDYEHX2mCRQ
xnfCpYF9sEAy+aFafeyR4RvdDwvVLgRtHdPPawuaMYrZPTe+lsZsmw7gFZws7CUg1BDhUoOQNqwL
8Y95+gpO/SL/0itktZ+YYN5nZkCk9gEwb8M4XSQVSozD71shX5YCDi4qtNzOQAUifFeU7P6GUd3Y
Y4Rq2yYehfECNhVZV2ubzVaalVfbUr8vKipy24ce1ho3ethV/AiEmWh9mrBC2r5a5hwlBkiq3P2+
Rd3GuLvlXCDI8ysbnWPvj5H612cppXUM0t0DJFHCWNDuLgTUm+46KxuzuhX8hAYA1R9/F+rPiDuQ
d5W2AdoM7bsSlVR9MSSdZIRiP2/7/81hNyi58+tIv4bgNZo+wZxUv2Pb7rzBJgg9nV7lknXRdbgy
8Uw07gA2S5ZG6Wfm+EcyX5oUBERx4JwIAs3LqYQSXvuwIjDaeTy2yto+03s4hkmKHtyvK2OLRtd4
zhXDUEtTnHABbk8UtJQLy6AlXtTRsZMdDNRNcis/mmZwqNQfZ670PZR+NSTO/oBa8IL7SUzCQLAV
zR3Rvrc2pkLnyWuYt9oDaeNma0vTjPgAez9cqqVWDdUGLDIr8tiYQOLqC9+73oS2Ei3a26H7zWK3
0Xckdm5ArHsIhG/yE5ERW0Ja5Zm4ynoomClYgSb6NTz7dx9nUUFg/8qQg42+/TBZul8pmeeoT6fr
Znb8pUM1h74AI5Ulw/PkINNJ32RRS9pDttO4nFLELYZkHQeu1mliO/J/NsqUbnAVFLYsK92SDVof
PyrbkQC7s1rOXGC8N1ylopGWdyZRGyaQahSTglPCLjSlzNjfDxq+SkFFuGnFfAAnG5rxONjXW1sy
h+tDn3eRKn5x9/bflKkKG+coljwbo8AA5qBSbg0Zo0OytorJMTkMsL32DazXRkdov29LVJKuM4kB
+KXm1vN2eRCnm9ybyygOkMTeyw9mg7ywrw6sgqhAN9yyxpE5FEMydVl3da4ZfQ7r846emB4UVRIU
W7bN7+SHWqTojOoJ/x3RmUsch3Fui/yKQH3rQJomM0w6m1N0mg9rYeQk1CFxeUe57WhcVVMfJrUk
OttJHxQGeENTLdcwYUnPRKpxUmhOBULdqtC+GNstMAMNufF3rQsRJZYjszTmZgg1YMZ7ffgV3V/o
VBcUT2nMV9QqcBF4E7nthZ4fPqGLpFaZIQIQaWrSoxJN1sbcAFHbX585r7kITufrns1sdo1MNYQ2
s53gPOVh+963saXaVLAd1i6ITTw6WQAWQ7QW//TwLPbPeNSwyKRrXIIHNI6YnaZY9pbk32RxE75I
4/10gRrow3uFzGgugKKpOgGQQwvjBXYM1PZHssuzWKazoJM8DM5BABHcdKFxXpFY9G+MOAGDHllS
PGNNeQP6T4NDhRu/Z0aB2QEhtjjr41v4rlFsOjdno7rzXxFc6tE6kejISLomq0A6ALpIZhC3UZtR
7DH8jW2OYF3UzYY/HPWFEzWaSy3gs28y3z3YreowBMOMOB8RmRw0t9pDabmxgDnIfYdoxWO9VK11
SxJkLDSK8EWH+IWrzgUmHCaBDzPKv7T/mhV0ESyVGigK5ts1D02HK7chhIFINWSytX4zn/apIInL
vreqWKJjQU7ZPT5BwpL4WWzvZFud/Vx8fbCOX4Pkt0jgeEjslj3csZzoQyp8gVM3ftqO0IYV18p0
dFkzIIXywunBEyepbFgLneP92ebi0SK/6lI/1gX+Je3S1XwtAG2BIO5cPvugocg+HrRorK1cfOED
HFCpzjeR09b04APRa622uDxIPQMJh9BtJ5oxVE3L0dBUknf1TUrhxXr7w7WUtVoD0PeT6USMAPHh
WpbhHvoaTGRTQvnLwFIv8d17ZCKhrn2H3m/k5MicwYal9lGXqMpI2d9pFwZdbqty5PAsaOnBQ1YF
ytncBDp+kq3GBeo4FNRvtDnlWwfSpqJ4cI7/anGRUL0rQVcYHlIfqo+KKDjr1AfATykj8y2mLAL1
1h6YkRRXvqJ41DQa3hxB2tkpxSilC+iYVKj2P3C9YZKBeyHxNcM/dwbiqF1heZIY8kvODySjO+FW
NHHpKi2EM6w9NzJGgmgPQ6goBUaAzaGymRSrQCeSqkNWtUrCDv3eO1rTcuZH/zwqi9kpitNypLFs
+gpnUq2K+dHzAIW1HAP/JGxRHqFhoSVhI0O4UpV5Kyrxy18IN/0Yw4JL48jZBK+wKjElnpwqufGD
5GjPhMRtgxs5/b+mKX75i7rmsvAf1/7SSOllJfPNSsXeRNH4TAny2Ll2uZvR+GS3aeE9Am8PuYf7
1vlKY4i+nweDrKxRMUPPIU7+1miry7JIO2cjkWGJggvb2oporpm6S12ZuCemlwXz0BOE4ta4DKDX
mEQQE8nYUkRcmtROKZJOV5cz/soIjYPzDnUW9p4bzbGD4fBCqEtH2gOjjgWpJ6BBZTPXcCMjCQM9
sOFmbnqyTqY1PdHGrEiFYFlCOnBWPAFcB0EUi0K5nJke+KYx7i/rjxMkFjOX8I+aLmc0bSk+UAOm
KczeCN5AKRcUKjzt0zgi1xfSiAk9LF66SSrXWNUq2AxCKNyBVr+KNXB+m9DFnQUzEVDjy1ZqKKqK
UA/Eko8hw3QWha+QsSZRvRUu/ZoSzZcVbC3+ZGNuZg/NXw5W6kwCxFI/bPccID/hIJaqSJItECGI
VsJM3k3TdgxFRyJxOpyeyV4HNotXiFz8qhIb0RIL4RlPiQ9xJ14koz9qa2XGcI/nhh1E17rs7bLh
3lCmQalUKij6rxK7QAwSo6qjupxcr3KavNhYZOm2juTJsKto86ffWNfFAXbqedFwjGsb7WXuAtOa
a8YbvF30yvPpVwtPPDWK9jDbmbfW1XJ7Y5bNGpPkrlMK6nf8HHvpfYLWvjSXrXddPz6FtLENndMQ
Da8wYS6nzJ8WFDPXW5+76iovdA2q3WFofX2rJRsV2o06M/XKzkYSGPlzB9IT2zg4mBZ9bFU0yQv6
iL5ezQ2lyNRSxCIEcYRoJc9e01TROBfwBwc5+cDjDsZ+Iq75XIcBjqCoLY7YWAmvwfyYTw97eZvy
wtdNZWCzH4fhBoiobH9jTA/3uhumat4llK/kuxcJxfqXMiog+4RBffjtkrRHb2/iscpWQAmBqeCD
lfwyyZUCjx6v+M9+DTmqlgmqwi1rFp9n4KJnRO7ESwoK74z2Gp2oM5zX6sMVcK7RKzErJn3YaIfu
Y/fKV4sr7U6b9rgakhMpWJo0jPlaGbor8pHnDMJ34UVkupHO78R6x5IZt643oxQrLAc4Z2RQWkIh
wzWdztbm4191l6p2J/Yvg8Y90YISmbSv8Hg+iPF2KpbX7z3AWw7WyWZN1NhPSvsJsFiGdSkx0hws
88U1nHgwGLVupx365dC0yOqsinB22p4W+uDnSc0m/6DENiyazRQUKIpYt39m+hvbRoG9dy6fUWuU
7FUsi022ParVoq+YqZnvEfB1ZWGauAlIHz/mzGia0vnupnxTLDDEstR0GmTj5JIE5VhfWPRbJHmr
Aw7FXGfcEstYO3T0PICQd8Hh+l8NUSy7fuOAW0e2AilpbMjfLAkHv2YTC3dlmIQe4bNsp7gKJPFy
iOYN+Ip3WF1doL6zwmw0d1Qsys0Q3GT++yR71zmbPp0zCUCemNh712sDgi3TglCl1oMq+KxXAQdS
YBlPESizCC63UnVQALeBvRySGDG3UyztkWeAmdJzHyO1pcd43mCtwyQX9OhLG8nz1PD8wgmd62dG
57nIaih+d3hRSivW1lliPi/YIRrGIV9JutLUgSoV5zHFubzaYdJNTNOmqohNti9hLgFgwhspwjvl
KzOxSOYNi6s0C5pwtdGEk4F7l3XHDorEyaswBBtUaTnGXLyUZowyxZPqZq0nX8+27zIWkJ6AGOnW
z0PosqHQ14DAMWFrb0goS48m1nyn7lJVlViu0UujnoP5etKFOTTh+sGo4x4fwwu0lwBD/9hc+rX5
nFdXV6t8+voG86il9K4ILIEjxsRtS1XjPXGdzBJ4dDl6bh6S4IWlKOTeYOKFj9emQnP3FLrOQdXN
bxpn+TqKnkK0aUX22rKFEQvR1Fanh484pF/GOwySLPBervnlyCPrmHRDKTXpTp7i+nzJeOMLvGmk
v6VScSq8vR5re/WnvJvW3N5qMZENvIXWdXGNoPo9LXG2GZHNXJugdq80Cny5szKo/3C8hAo0cJh3
uFVVi8OuUXIg+BKJ3AKJ/4BjH5dSb8m6XK7svilTewrWEuSXB/MScPvUDeVUcWGr0/l298UEceL4
VtWxw0JErJZ761vAnXoLIyRU0vIh6ZeS+b2ej1Sr8yUBXiqRdfAuW/I8+f8hnBinHhHmpZ08HbZL
CBZLIyA/NH8a+ddJ59g7y3Udz367rHZSU5aOpVgLpjl4hx7BoIcHIxO3q6KHzhLKs1aLKCCNp4nK
paV8TjOPLQw7uc83fOmVKZ4JbC1Yk4qUYs48UWn3zK3v39I0Ed2E0tX5GsMsBdVFwpe6g9wI9HPq
HGJigk+gBqUHBoA73NzZPMWhJaDdyg/nhfb0Sos6KUqTb9pWljBwkJ/D63FFnbJ3bvLJTRMJwaw2
uUAGH5OKZrpPZyvG5bNAsCj0unxCFUXeUhazSWPhDKLzlA126OqNUx3oSLzr2DGnBt8keNWg5fpm
522clj6DZdoh8p77194C9nIYBMvZ7OiV47924c2fXgSmcF2en+rchTfVo2XSTOHefSJBKRTKb3VR
REPIb3FFka2zIqT13qU24gJvOtl30OmWWn0mrjSmJkeANloCXfpLl9FjUtahbwqIIQpvnxbXKE4M
8Qzcdgb14kwHJztgEVk0G+DcclxVokCsLebHWBuS7xHyaPQY7YnNjN4S7CZe6yLFO+gW1iA8O9SA
NaHI9XYeUfuAWhOgg0g08dCBnUhlopYUMQShL7CQIY3m1F4jgf//vXd1bp/f21mels/H+kF39RRQ
L0hZ6kaZj9jwW9G047bbX65GWOiZm3sNAovtnASKhE6guzZKHdB8v2zPjthRFg44PkId+/uW9TdC
hbojEnKDiKXlhzoHVVX1v6gU7iUyWB8v+0GZjACqSi//e7cOCjAyxxHY5VBchec+uC7r8WgjNhes
PBrC4HGr/eP2NR0FT1DuOAejkey6IAlqagaS/jNlmvPgNDciyuJWEphIi6/HpglC8Q4W5moWHYmj
5caGYx7SUW4PFhRhejKp4V7Ff9Z8nWiXJ/ljFwPJijr+JgYi0epv/INLGdRzOHDMLw7TuDonff3O
k7UkGmiDUPRk46w/56HSARtM4P1fKZ7NKNtv/TPMgn01jyBItXFqC70bYG85vOAYlT2iEx7yX2uP
yf8ioAFka4EDC7+6R81PVQ1DYsyI7NgHvCREpfu8S++TIuC0ELnUJHtQbM6aIerk0mou99VmEG1f
OIadG1Osm2oT0jkjmeKaC684u1tdnG3htefGL8JaqMsaZsSx6UKXCFuIeoJ86I4SdKx5u60w+P+H
9CC7WXm1enghMcnAtgsD8zCGgjHvRiM0K09a9JfRTjDn6iSZ802bPMoUrEoP8qBslAaVRSrB7+1d
iERGdyalOuQJJaQz4jUbMpU+LjuK1sAx6oBrlLPHL8tUuQyaoaCZEdanxXwEY0h549WhYr7TYL38
FBgrjskpVg0D78FZgVUqp27oNsaCq3shxYFVxX3ZfytCOTU0Qi80d+xjwryDjM8VbFS5UAs/qruu
oSjNrz0FbHenotcHpQi2qVCO0VOiCQnnNYODF1LK8mqUzlcpAMMeUhcNkASQK2O1cRC3a9UlXBwM
RGkWmFZawawhn9K2g3ymrbjoK3CgI9m1io/EknBSTNTrliocWGTEdazbXkhZkR/pgDH/LQOnkywv
jf/XdMkllwV+5GqTXBM5LHKhzjJ8zP8tBMgpPX3A2MWmt2fTlGSDwAMw4bv8NrH6hxJVwUEReg2u
k3YQ9dO6XklLDWyPdL1C9B3c7K1nxIOe76kCHrb+3Tc5k/3PZtv5uVpojtegh8xb+JdMRslPIgly
DkfvrVMjvQTB9/Y84DkP9/Hh9ARQoPsacNTuLlc0vBBRGHyWsIWVzhJgJmvqyJIVRcrmq/7iqop1
gJoORF4baW/jES3/2VT3Y7seIdsKwansvnq+T+wQIYu6SvaByVFrbUU0qMFic6rB1hYYyxsO9CTO
eugeKZtQgWAH9GqRUF0vgoUuXw/kZyI7rp/4P7+o6KXB5uhDkidheovi7NAG0r5c5KCXTB60AVNG
U9UWExRm7uEddw1zSXH6lzXOXUFwZS6mB9mGuxnyUY2lD7T0C5CkNtlxKJD6X549u+fpQ4vLic2A
xDOKzeCdrOWbW5kNDmZtcyz4+A/uzifo8MK0zEd5NtNu49LQ/gx+cnK/S9n/MQkUR25nsNtqy3J/
Vy2RMkXVupfovbLLGYjhbYGGSrqYnRH1uGbQNZidbFE6UEA+7qdpK2okeZ+8D23XnpHngMnuTJ16
eWMcy8kcmZaOHLSXIhuqiabEvVHDYuY50Tl4CGwGdjyRWPkAiaK/b2z/h8uIfFL7KRodYP8ZMwYp
jSPa+rL2oh2144tktNVhFIs1tI15Gc7qBcd28pxL8fagEZmPiK5wUdSVg+TjnigRrGrwHR7z2iKO
FZNrgLq4qPYeXuwfkRzKNReTIMvHQIGj7jzP9a4ekQ3WPW9o5qsmhp5RXkZIVamKBRnM2M4rJeJt
Dy9UFmRoVwouXAFmSaWkQOD77UxV2PtOJtL3NIKQG3gtgfMHexcYeEmCzL26ZrHOcI5ZNQi+RmGw
72AUrt7vrDBGZBHIfNY1DS4vrNrKj1V0ai38Ih8Qw+nLCqT2hDUPbz3zYsRZ/7HYNjkF/k8g3Mjh
58aCc/SS1e1P1Ze2juBDq4BGPhi/WhIo2eMblqYHz5OG5qKxr/p8XRvSXCwoqOWHSfbnapwioCQ9
ytHaRAGwtF9d/rtYWzYJ0QQLx663D3ksfgx5FeU0KF2fBqqfb0To5+4mKttmBYMZnBuP6F8SLB2u
jZRz+HDuNAjW0Z/T62bfVv5W/q1Lh1tHxl5WVFP38J501aE7LGLu8SNKsjIf6BX+jBZ1bLWyq0Q1
0Z7wVlzaGM62B5dXXWL3O3teYcdk/tlGkN0MOvOdyh3jLEnDw4waCcCaoJSqdpuLA8nHqDxoTwl0
mEld5tyqAYgZSjaLc7+FsZn496D5XLBT2HwjrwpN6zONtvTdbOtSM7ZmQKZEKd39LgLc1lUW1q5N
LWrSE0CWVPsESYD3EaEPGxVu6LsnM65P2uzD0QXziskNsrAtMtR49qejFdZrLILRZKb9Uy4n90uW
gunWVnBIo9OziaM0QTrlgrWpbWFIGnwdZZ4SZhmBfPDVLNvs1WPd6UDwVU75dl0KOKV7bA4kEnNr
oVRsaEJjqqwIRQXRLI/pndbzZIccIaj9TailzSH0OQmuZTCWy93tFoZlZQTengpypSoqQrzjwQrb
Po2sjtj35DJo0EQP6FOQaQQ8KJ80epcy5JPiTqG/tme2cr8tJ1YGE92B9xwgcm7hlA0Pfr5SDCz4
M0QYc6yYAH+folOBUfmjokaiRcFtTNMCXx0St5UtlCRg6HhuWn8nisyjuNJQu/EYRiVebw7Iygqw
kBlEYGo+t28En0+aQvy/hjqxuxz0JdDp2sLIpQkBVfdlT6AsnQ8WkVvb43bcHahHdeTNrGOF3JkK
1gLM+JEoEg7qFS337ph8pBrb68jVO84rj8AcLFDlPVPO96aIHA5TI2mn2+4lZ0+3f8FZnL3e9Ooy
r/HUU4msFPUmw85yU9F7P3i2aef2Ak6n6OeD7vyYt1GJh6IswVt9+45eM0VwDNdUQHw6kdw/483N
1LKrNn4qvPQtuzVRj0egEctT737KBCtxJJ5ttgEFdIeCSZ0vKXiUPyMBWgEUukX+CR1kGMI2t5k3
I9ITzNai1LL4N8qVB/N6sw6+CP0UfefMqHYbTBaJJtG8nOLSwDy9gA/QiqgKjebsq/4ne6aamJFV
vkv445kWykrzmXHx5XTIAykNXrRGJtGnCovljF0uu2d3Ur0D1kMuDuw6qrWKV2gRT3k9+obFAqk3
KvqpMgFw8CFJRjPmUMe/W5NAj6R2jtJbTS+vshFN+X2kAvIqx7Gs6Qys3r3pbMx3CX6IFULRsqBo
7WrXq3N5tTa2HZLm1gyOl9Z6lTUywpsEPq+UtS6Wilxs0/FmLeVCsSc0kMVbMZysmYRUF2hSrUdn
HSinObjGXWbInY/jP1zcPkVEFQVnBJS0NP5l7TDNvLshkayJEp174kJ9AfYAPGX9y941mSphrxrO
d60umENcRws72Pl5Mp1u2gHO5dAKydkhPMv5qZd9MeEQUk+nlTwvusX/IdKf6Cu1mIoJSyYLtzYA
7S6bsd55w0fa6Ingd6OkOsIazDiiy26Hc1yav9GSMuuYu+uV70Y6reSme/JtzREv+Ar6K2fpRAU9
tIBL+7wFvP1hPddfBQfH+ia0yg05FWmez5AqJ8bUG0yTPGNc7ZEa/hkvveAS9t4QTy6t/db1ngk0
3wLvtJCnWYgIP4/1DaJlr3WQD7436QfGcJT0Pvnspc5BYDonh1PLxgJev/1Ek8PBPGdVFwUUltQm
sLoHczlL+SgBMDJQMjLOgqjCADv412ApMIYZ2pAfgWPDnWLMBiO/m+qlW7YQfHUNhQ4G7nzz9i1A
y9Z84WvLAT7JaUxm76GkCEmW1vpGiAJaBupZhtSyI12F06guPFdNpixX3DzW8GtIRYa+kmQceV3+
GWomJKHZynaJCJr4AYpnmKUOdGQcytMTu9mzA7VyjTUJFaWLVPuXCui4DRWAr8TEXfr9ksOKyKqe
3qejpPGzzPfSeSmtToBsGBzI+Ga9FJeqObtcqsQ/qfvW96JXDb2IHZbmaH66oF6BEPamNMz4lZPW
vMvb2WjAghevQJzFA/gJqguNptfaK1RuheLcsFOMc/GrDqBVDQG072fPk7J0mGvbRvMSjLjGX1MM
1QeDEZzxTXk+bDHlSh1CcGbNN9rJBjp53/AGgT/a8XOr4nFcLEgrVtQjBcA6GGhuLYBbcXzvB0rs
d4TjB5NUEnqUgOLI0jZZ2PdUi3nbVsz9AgQydmvKHpC1+h13Qrz9k7nUUNFwllkLbqq2CDQzWaEn
dS4N1wnFtgM0leXFnkTfEC10Gg4J3q5hYmbbihRjtX+SfQVCthknEXyVlkEenpCvezE6Au2ncXSm
6Dn2P3m7tVDH3fynTH9vS1c94jUgEQYSyWee31A3Qds9n7YuOe2CdLv8FuN9FK5zqezK05jmgzOj
yo4PMSFfyVJyypcaUqt0FZka/06Nfs+WHYnA3MMv8s+NBlKNnxD2s5PP3wO4ONu7kZi2plsQ/GlK
1xiU9TJEwOf2ApfAdMiv1453lSzV2q6boRpVMGvTxx8lCmltc/boF+dOYvgldyVw8GeJASGrLT6/
TXwyyhugnZ8niIB71q3uz5QMXOu64mUC8Rw8fK6xvUq8asRm8UnxVoRSEy+226gtMnR7Kt9iQCSt
BgMZUhEyrdougMjJZq13rE40c46/CvE5C1Xwm5M0yTu6Mqk1UxIFVAEN8xJOz+2l3mRPoyj3OE1p
ZVRZtL2qD1cPJgaCAeWZe35h8Gb+8aV9+XpB4dz7f+g6aYjEGBPrinzxC/s93KJSCh32cXKe38BG
wMhkC6suMo9DKg22ovjNkFK1oXlMyqgIVXmo+jdp//YK4CQA9lLbUwB4/tZgaXxNAP96ZGdI75xR
4u3ybmDfVL99wCTfAeVDYaV9Nzt/iU4OTjITnFmJkMS2Re+BrMD1YeeLCBhZTsHoaGjltIr6GzoY
/Rsgl5RzR0p1lZFVBD25z2r/D3z18hEX3ZkvE6bbC+rumTnza+qZ21MWmPs3uhNvr2S94h9KT9MD
t69LkNWqPpOFuEJDOq8ZThFbQ2y/rTAfiOXLOcgW0GZ/nAQblhOfeGOk7COEOCn21hq5EJOTSZ0c
MSuHS1WADRrSkZ3+H+G7X3hHvTnM+Ya5WNS35mwt1rHxoUi611W5cbxI1+FBOa18QcSPw35ONxDg
9bJoYe+TWs9g6T+6dpTUnoKUdNi7eMjNV3mjIgPOSZRumDXqjmPp2CuRsUkUgpPHNk1G5DRRDyWx
0Pte6nogHCtJzGtQmHbl9D83EU+k7nysh7dUZFebSMrOoHUEcgdPHd5EQ8I43VUwJJL86VjVY/9g
9LQOuh/ll3Oipm1fajOtpFWZ3ao6bzT6FxT9rCmlcBuGNzYdkUcEptlK31cH5LLyT3+/cFKG5ZVB
PXphSwMZZz15OyT8u5/TYL1LbhI6bVLpdYee9x8UKSoqMue2fp0jz56kOnKbtwDjZAZT8bzfxFZq
7IGI5adK7mCXAPbloCimx6ZFjwDeP1sUZqyLXLPmRMjMX7m35PFYIRtfIIjOcxk1d++lL9Aa8Aps
vO1QBSOAvsY3sGZs3rbie7gzJhxCH7s+rRnGM/zEohHbiudGnwXIL2fkmxhFVs6QejKijK/mlagZ
JIhSrHI+XgVVrv+0W+ixKlW+WdUjdPhwlFkYS/5opl9RLq+Xk/RShbI+4t7vueGslltsSCyDi9oA
BAAEePOTGiwpX4M4X8vY6vgPrdkJBg3Y+zHGzh/KZ+p733YCYtzjVvBQU9Ki+YPhnULuk2Pat0ZV
k8CsN//F4ot8oLVGjkilTiF4cJRplnqttw2OONUy45Td6Occ4W8zDp0O92Fh7Yn+U+VfoRlT0fWv
2j9Yjar9B2O3cZXMJ3wzGwCXvl2vgBFdXF5af2G+H1hMnzhld660xcIEHtFLcu7ef/0hXU8dJNH/
kug3miIdXtK7rYVhjyLcLdsBmkWJv4IKKOfTNWHoC6GkfSUkVItdqRuYZxfdE5lqhkxdGJwem5Ry
PNqxZByEOY0XKG/y3Ija1Pn45UoPwPlLf+HXtPuP+iTqv+B5Qzo/diSJl2iDpbd1VTiUOGdnbyd8
OUDQ4xKWLfbJacErxo0jnlSoKz2wElpQDICUVpDTuugoXvBE0BjZk+QHgC5Fvnu81elpcVWw1X+q
iNdMLCH3kveXd89QbghzbqWNDi+bL7Q7WzCGO66iLilO08c1KeB4PscglxJRH3rUz/HQE1GmUx1N
QHGAzuxF/G9GplBu7/shbKg6aK+HzSECth9PfEqdAsWiAZvhKfuaxhAD1tkKvP9cbL5Tf0vZkRHX
/iwJyGTXzDV3YvxamkfwzFWMaNZznUb4EyzVJ60K/FUmEY+RdzKEzd2wcsdEewDRQfpqS/w2nWv7
2hTwbfZkG4hMWCj0zAR0uQlcCbAKspZlIBkEjBjj2HqRE/81rbt1uWdGE82la+kK15CMoUnKsorQ
mQmrkJBt4VbhaOUnBkxZazrRT16Qgnr0HQ4mYu2sEjwvODpRDa2hFCKfwbLELA9w12et30feGFvk
Z0xJnu5TrQN6PNTlkOAuM9kSIGPwsu8eYZw0h0f1DOuWoQ+lIz4tdYAeG946wx2o3UN1n4sdDOi7
QWZDYd1gIDn07Tl9cvGEs0p20VwgYSNf0LQKxqET/NowILDj2eMhuvsRbzQstLkw2rbB7E26I1i1
TYFT2s4F4DzQOznzTgdXCmRktCeJSAjpmdCJDo1KgqKXhBpVC+VgViFq/I2eEh9KnJWDrpMSp57e
da8r/n5fLnutfkGhOGEmTPttbSTnZutp871JuR17K3SkABdgkqhu+B1SurdNt4pdpF8BqBnjPNvC
xeJl/NbwcYkyTFZhkFFS7fkkvu6JEcZSuWnJJvIyea0A5WIKokyJR2G2DqcgwbCXN9RySFsBF3Qb
k67vN5MB2yyFg5gkOYMsPKVIbYh4aE0eHU9PBmLVnpzCuC34v9i/t7GIq3ZJUo1P0rAoleh8Qugj
9h/muH7cpmouDpNkg4hhtccctVgUhzrcKYfkcUJhFRUZm3iZX7scFI0tj2QH+x4Acm/98Oyozzr9
wMmHCSpasjH8iDe2j3RJsCGQHYb//qTbLjypTjncQOtTF9xlbMCzT65kFY/XbyM12Zbcfm4LhzB0
y/pOnYr/+HSWGI6tufnyJaa5KvXyb3gq2zRHWNs9HNjm8T+EW5gRwc/OibbfE3mP1EqwfqkG6LtM
2JvwgzSZ3PAbdMmrDKKLBS3DHZO2AuDJ9pgb80uawhZ3OPAYtSubjdTGCzVhrtETg1ao+r6InRrg
0hZkVXoP5LVYdN7u8qE786TB8BxX1+Z10qGa/mwxYPgB4QFWp+ruDMMfrTqrJfQhRcmB2YvDpjGZ
Dcd2j0sLFSPQ9s6eYymIU/J9M/k01R6wdympxQMl3ngdTfe/MePQlnS5yG3pzRrRIDiPiVkd2Q+C
YJB8wFr4VbdxLdMkadYNr76wnBz7FGNmdHhzSIBL8Yn401riyFH1HYFkroIdPlSlHkqkRf3U4bhP
S1s7I3aTymXsN4c8wBy6LNN45KBmkfGkS66JNxQG8HMaWX7uGT/ud+Xalc7FguDt31DidXeoewEa
OawH7r0ozf7TtKQhiIl3hwn8OmzTpWUjFb4rgm++PaVmvJa3yo98Xs7YNxmjK0XD/cIBCqAxBI6h
1Un+zgsFaW//KSTRuA01PRb1erfddsWH9Ml4PBgkZmF2NTxkyT8uWn0gyxRRXW9qKB9LdfeNAwmv
4YIQ/8XQtjXj5qcJ4eLkWcn/Z3TYNtji4V56Ds9Wp/jdkKBqyprEzWpdKzREXYgumuu3jlJfrEyl
3lzgYjMvNgXEJVZweXlq2dGgZEZOo+E5GmIWAgBajpN6tApY7Nc5tC/cPj5YohE74iL50I4Ds+vC
eArPAkQRSw5unsUSINUTS1KUln1lTc+mhaQtflIVY1XSPNJYNriJLF7p6qF1zbKTOxB5HwawPpqC
iVx0uncfKCokg7CDOWBiWH6tY6Nb2r5F8BKjSc8lD7fr8FLOo4L3768vdKrDFhM6CXoavPZ9fVhI
hPfrQrexJzTGFj7h9CeiKILDp/2Fce/laXf9u0ap7BFs+MXPraSfbosRHNhnrTMV6+y0XW8DjUJw
50+rAf7K4fr7R2rSaLgMHmv6nXtBPJUR+u6+EPZCgWAzzotwxGajH06BEFHzoiYitJrJAfbSebnH
Fw6ZcSkWWJNvmRG7xxWJBJDVXtVcGr3w7ayCg/dmE2570RKIgeAYqnw9O3ei2Ky1Gvnl8MzOuOsJ
6tj8eL5iqAz8miYlExOZcf7ouGyyhq9t2D0DT68utMtXyVNS7A7qhwUQTXnK7gIwQmBZM3AMxtr8
+UAbp/kC00yelQT7eOfwULZKUZUOgBi7CAhKFfF+jqMzj89SBH/swG9zjMI6E53zko6ymRP2GUFe
cGUE/jSU5+UhLfo4SEs4F4YWiNsPN5Nku1BGE9SXowQuWGy5FSVnQHeZISwyJk8xJzXfOijg/IIE
+gsQTGSK3swQSlcZKQIZOJAXu41CWaLupjJSg7GRsTj8QAD8hDRB4BFqctusewNcoP/qXY+afeCt
pQBzyNgFJZO6IU9W+TQMLBGgMKClCAeeBIBsF4v77R8IajUP61/DusD0sx/tYQ9A94MTRbDGGuI3
yo9Jm4ffxOTeVd3ySQbj7xawlwB03JfSFWPfqsLtU4SW0GJYosYFbYSB0RGiozbYrpktrya6VE7Z
fA+moT24ItTJnqNWUQWCwYbTo+2kob+VyUXIM7ZtJT0BAjZ68JdaGKJ/mdxuMfrCsQlcjw4bq7EW
a4Ee1DLP4v2x6nz8kFKsCpwJXoJNoNLXdV5NbEyX2PqwUe0ZMIDxzp0s4IOAMOJV8kETShM7ZQ9y
HPDCHRL+BCaoJjk8+Peb0gTpgbFAWXItscFKkMIvEqS5vruscc4G7G5+fDeSKmQgUKErNeJS0p85
XzXSN8iiip5m/Rt1tnOnLFBdtWMZaUFMraU3FSVjfk7YgaUQL6j8eE615QcUP9roNO4OXDl/rt3n
HWIENd7rVwMaRV0lpo5JjIcMXXkMBJN14fUcoPgrUbILhinGEDfJZj9tqOCtuYAcXjFNug48VWMs
Un5lftfYuJdUsNGD1M+JfZ7mGLNUD7immnwYYCWZlm8vZfOh0meamwioyK7NdoNfXdcfWbf7lPaR
QgZkO9ZdFE+U0zCtmyM6JLlF5S/sOcj0jl17g6yDJJz6De+gLUUR0ivmgEn8y+GCJvvFnrfZJO5c
Bdz5JLxXh+BF4KVPU2qYqk8BnssQ5slRKbtdjZ+46q53jihY9RVenT2wgF2DkGiyIVDM3yhMzVgw
B/+rkoctZuhrQZmFPBjMr+3nvYauLPSTc2MzXgiPXjooe1b46Zin6OVfI+owP/ngiY0eQJf30//t
ChtyagpvN0flIHBI6gRSWdz5iYRAJOS3WwezYuBEXTJz/5M15hYz2ptnBEGs3auSfQPLzdAv8NWd
AljskVypPRiYHtb3YxkAC9APMuENqpeFK7C+sIYJMpr6DPTOqGRs19/DiGQzK521LZWBWlcgghaX
nyTMBIBwU5xWHC5SKb6h24Mt+vR9zkdWc4/rO8eOiAH/Q2XlFBTwSxIdeJVVR9QobttVLt5lKHs0
nZ1rEJq5RBHw0Ck75hAuuzwZZwNjhw8pa10GkdNDkTm9TgEWl+kPFlnfZajUpjVFk3KijeE0du3U
7N7UW5iquqbt87xuBFl/kT1P8jVtQjFL4SoDTV0uZH6Ib9lRAdnEbrWYbkuxTEqB1XGMgarqDG1E
pcVMaTef3ZXNLh0ssD2shqRnYfwNKEYkm7xjnu4/f5pHPdFqdZdRzN7hCcB1dCsg2EP/8Pzzy4Sd
mGOV2FlHr4U280pE9n/IAZMYDwkaSqM2sOs+bIBh9ICjbvw0UAXmybpaTpNhHEaSzcTV7hSbHvIn
il1/vxGNARrtUgk3SGgfi1bMh/QJNk59+KbzKJZmDc60MjN1odEeoDz6udiOf7FRg8DV+uxg65d9
yhzbPF1qkpOmVgF1W2Cq7mcsgMhTZuqWd1FB/kVAk50UTMcf35nQP5T8q/9pBMRbUpjwA4naBEdA
GoSxpFvMEB99YVuzNyPZT0wjDyWH6K+eZOYSt3kqyS/4R3pIlB6HXwVnGkxud4RYN5iSwj9ijm1x
w1h6LssA8snkjCnnnTG8fgVvGq5o15EK0SLnXllQbLUPnVyU0MF2PEtTIRbS+qGYJhLzfXIcIMxj
7zjlI5r1iHf7XM/HG5N1/+0Sshrz6t6LkXbPi+B6sqb4GKnKpz9zcgnwvJ8QXA7pnUvXw7P/1F01
tWjTMDfDY+1Cx8HhQkPYQEQ2CzdUX3MWWAObLxQbzkReigyXt8BXQqmzofO7JIhIEu92RFepHiR9
YIkdgo1yk2FcPFtgvjpxsgCJBxmREYZhmIxrzP2Tx7FQ3ncF0+A+23JIrcqfMjf1saNfVkHepmBN
Kwv4U/SkdfZcECpp5UN4pdcMHb3QnBXG7QAtFZe0GJSKRdKJpVvJrPiZA6suDCYcZJxfHCO9p65i
RtcsZGK8FdVV9X3pma5B4lbySVEUhF2IkN2ydAvLxdL6idXuGT3VtOXCie0gtdyDGSqH7wVu2alY
HFO0J5t/vh67/mRmO3xV39obvv5uiMZi9FTA6Ot8zVZUVoWYqPdF0HCaIb3837LtbEXfTBJDT83i
RCltZjk0X2pg/qaV4B+U2zTjIIECitgWfmflBVmOGbrnAS9eEweonIccvoQ7Gf2bDm2vleLhTpv3
Ww2rqaYpZ/bEw3zMgnV8W2vwc0cHGT35jrrWr3W6kn+YzfIW12FGPqPYNF/yaF4P3xQoiWvmkWWd
231UfMAq7BIsZyIkekeMShe8PpSLMJJxla+BPWs7rYgOoK+/aTeb+158r+oZDoAoxqhSobsqFof8
uZ/tuNEpzFzsAsc9P4xvf513XAvH9nMz7r5RX5M0JfX7Bv/cThG3Ax1kkK67xsQL93KKrHRAkH61
l4XeeoLLnNzigZZlNb8pJ8+bPqbspAH3bIUhGFNrfBDLaUzKLeMRsCjvlR40JcDX7JUE32SoUYVe
VljvYexJ7BHD5tE7tsfJ8Gjjv1Ja25P7Ln8b16aee76e/9yd0qqxsaHTBfJX7VMEDBTH1Ll8+GAA
1prw9zJDg5HqnOt3DqSnCazskXNZyS0aP0EDdSBeJAQyogow2ifaTWZbKMseXuQo5sIn8g506Mqo
IU9BWk4zwS1a5C1lQDPNKS5rx3qxe3urAEAlW4jMDQxHQWJO7rjX2cPGj92PXLm9kPvQFAmvBUvY
IypY/S8HcnekI1Q4nqGpbaHGjFVgRETCsadCvudmZqrG3xcURoGB2CulDeaSi2yY9+u+hi10g8zQ
6PvU+OfnZQu/2eCcSH4UJxdGCBkSTpmI0Rr6dpMFhYYlh+0vEGGScJAiXKVtV4JtGg3I9wFPtIdH
vl7TQBnpnLIAmjtY4N3mkUgT+6xxM2+zRCJ197nlbZtpukcrx+wGOLtjmRhhsg2m6kq9jdbJYEO3
e9bsJUL73s40Yrthp/6YF7NG3HyEG04mLmPmdf5YK8L1Nob1A8fJGL/YREu74pDPOZIXH5To+L9Y
2c8C96wUbrLXYlnC7TSSHZaBYrMpLvLZ5fe+BefsnvkKkbBczLSTggahAayy480FbW8+TsE6iB86
yhWSEXDQ7gFjgSvInPpNM8Kt4poiMQGAFbU7YcEjui4PIAxK2zWWDOQAD1icZ/VQvsVj/7IGuBwo
bWenZzD28o4RWVWS+Tq1rK9GBlv68FROL8uZVfZ/bsFQuorv7jzduFiyTefggizalM7dps5OqQvd
ILIBAYxSLtqPqFdsUP+7ftZAvbb1gTsxwZbg/6e/VWU4n7kXEtbbiNwDVDB8q26nV9WzkJWUXY9+
eK6q/aL9iZJ+nDFlP5Ayt/4BU2MneVeFVcV+oOcnU+7UjzEK0BS97UmSReYWLtuw6hHxrFXdj2fI
k5EJSU03A81IP3C4S7tkmAupJ1OgOQN9DVjT11ojfKfRjbpnmQ1NJJsT/Th9KoY2kR0+Hh5hV2HS
ECUMQrEv2VxeCfh0SIxkxWN3nmy5xF4CuB9i1Z/mpyVqxyORd72/0cUc56iO39wK+XhJUtGs22Ll
6U69IKxA7XDap+a0kImF/q/sqoFksAJqhRzXBwjFj2zYkwBUmvItQ+OcCnXyC1VR0iDxz2Njl+Cu
fMFFnJm9rm7fiBUk8Pv+q1R/5M8oJxTw/QIb8FZWnHAs4KAF24K8o8j02Hq9NXkY1n1pOTeRfmOg
2ZGGIq20J675A0GIcaoNyEfQ9Ro46wpnBypFZs8P99NE8NDd2XjjE0S6eHSyLV+y42NOWcpNVMxB
j7/qRHGEqwfq4G788FXGAnHqh05JFCY5kFziypXhbtY3epcFjrbtcKFApzT19Mic/9DD0O3CUzsk
oPQXTzKqnX67P7SH2eUnk83s5jwyxoh/XRBhiBuSE1Qutxo+VQ6ChlrZeLI9tbQNg9Tc56dXYOnS
Wuv6chbyFqLOE0EseBjJoWk6RBlvutcxJaorSUF1Xx6s+gR7NaVWAnuFfyEAfeN1ACWPoP81Ulqx
iA77HzIm1rh75LgAnhJJmcs1EzMT3kmZXugGot0chJzkMSJz0jv4jTgWiJQZBzvkls7rdRxdxdmQ
8opRCH99kHnGWBRw9B7QYzElsN/vnuqWlzG5pL0sqgmVKOsq1A5fdqSC+xGrijP7WpIckA2OyQdS
XL1xd1aLjzkIACSUnc0MfXk8VqVihNMbq0A5m7bwdFPsH5nKUBC0gY7TdiG+6OlTZD6CAqGcxhzq
QIkPJsjVEGIqKteNUuPoHTEPU6CG56hlSSuAUZMi/z4GQmSHsGePogWToLHejF+78cKV2Cnff/O7
BRWbsizS738fFncsaYZdBIjgDDcdqo0e3CmGZK60kEIzwC9k4MGqe93c+1UJU7bnhCeXnmGxk54O
6u9KExxOnn6qMHuDenTA4ksJqHLHeOeBqN2nyr656z4377YWVk27mbm/BMv8qNVf24t5mfLo1hA2
lST28KJ8gBf3uilwJ2yuP1+quKWMudmLbM81vmc38M2KOuT9UryT/v6nb6u9DnMs8NkYoJSiAHX6
+OcQ66WsMhc8t6EyYkupF6c0xbIAij2r+Y+jMtFYcDKTL0Krk9rvP5xKmV0ZzeI99O7+h6pKK+7A
7wVPJ4znRdCb5ZejowLk8JBsjryNbEMyoqnkPrj27vht0GYG3EPEyNPIOyWjeeDMcVPUlU0fREbs
EwMCF2PMcdfKlkczfgNpf9bstnndjv3S67X10zzpKpvLRQq0efjqUmqY1trXWRgMoMl4ToFgvSTf
1S2kXhCAy568jhi9YoeF88gI30A7MQUVTB8Ywt/wvwiMgHLUIHtshQGI6gM+EL/oOIarbtw5mDWJ
9IPCxT3jtAVjHfgxGudleFWEr4+ItMpgVPacT5MKllUaePJD4km+Qz3bm6E0DqVOJY3RmQl8vX7Y
kSK4aoVOgcOL724ZK6atgM4zWNMkZLIOOgRvsvn1e3rMz4uOhnrRgWStC6EAQIM65YZpvAPTJgdc
xjBPEwBmbYDXV5rcJifXT2g7CJvydORlrTq0lldnk9aYX9ZTyY7jJokMSbQrUWaq/wLd3IVoSjOs
anmKCdVDQmZRHg8sEXCE9y0eivj2d9Z32XXn4gj3C9YjQp0q3zrdZTLppmuDyXjNDShddA1Og5JD
hRqTWN9sPNxl1nMAU94pHGLIuQNPj+zs/epjNyS8rgkzP3XiMpCvzPdxYSr3YQ71YnkVtQPU+WlM
WP45CzHfCv8Z+KPnzN251CIBYQf1bAqIMwAS7gPgShgv9aNEfX1m4odO/WbWncpkHm7a51KViCvS
yhsKeOymMJw8Kr/D1/EjORl26VdfTHGRg1ZBUOvTkAH40wPURGUEOQkbHkeQht10/HIYjdZHlB3V
qFDy7JCo3/pZuT24ZZhVS9V3DBWPjzy6OL9f6G4f3m6LQuJDw6wsRlLSdCldpz/P5XXkXt58V2tb
F+gHNjjtq4VVYSAt1zXtuI63Kf3P5LQ4Anu45SsMJsNpfNhrZWRiSs6XX3bXWABFGeAfDTs26PKx
/AoQRQ/3i7Gt6seh8/TRlz8iidVN8hgWuwtUhIQnLlZlPUnZlh7m4IJQob9itdnDlt3IkPHNzrtw
qMOxOHFiKTvTF113DSe++s4++DGBk8lWbj6yXZJEj7a0Lg5b9qvxGNw1Gim3Ivs7l9RhplVj0wf6
ZRJAMZ+KzRcVh/PuFRjiEUXR4/UBbcCPvSAGbDynBd/8qGWFGpck5L5buKbNZoU8aT+7KIYAY4qo
JvwQpT7AYaxfsMXidE7ty1ebOJAEMpjMEKWDuHduawpDFzE8Oc9MnkdluaQ/oDzTGrYHaIBRTxq0
dIWUjkEx6coc1binEHz/88p4wbnCGsYwahqf1D8YRkkguW4cOV1xe2h1PQwMAIv7K60JLeASzga2
o9ggnTYRmIW1PpQwHTutu0uCvLxc/ePVV24igPCIMXhLgpyaAspOzAHRfpQIFgYO+PoOeVxLDL6t
KuoRMyg4MmAC3c/g6fKyJoOc8GIXtAmpn1gKSI8MnVaEzBN4gt+sFXyYCT72r2I51AVQGStmeib7
ySyKk5nwnGoFkTSMXycuCOq4pO4g3MD0bHV4W7Hiz7HtW8Obe0J3bRmp1HR6WaOpDFTh0thH4CQS
Y+FLZNFF5ieKyLwc2yuFJ9Q3IPKXr5ScC6g/Y1aRsOew0iTWU+dKuaCwU/sfhm8YUF4vEitQW4qQ
QCia7pBu0gTx2RE7DcKOsboUAzccLvxEHDqRJEz2cXekaGHXFUaK0NiGoLFI6Am+VgI3mIfvdJwL
6N5pIFOK86K+6eTQra419tQ1JdXFg08zc2IfCQpArY+4/6Nm2nrpFJfTgGbhg5GGXgY2jAyAY+Yn
ukC42nAydd4Wi5v0TmEg/+wAO9EsWI6s/rFl+9r9lKdO/0YTpY5uARPXmjWtRvM+iChhuRCAOWXy
F+PmtbhQxpXoGU9/0E3of1QMpJPKAgBOk9accfvzUT4ZsNDD5OzbZRNgekg2NEpULp4oRUHuXMRj
BMeRTD/+ZTtkm2atfZgWkHZiBx2YJlgHsBDD7t/EzHMA00k+8GbDagz90AAbWOOtMnd/yKCMGlmM
/1qkMibhcMDFbCTY24W20aFmPFPp5cnk5nXLV2H43z+Vo5RHNdlmb16yWJGYoOLy55zjghJjFoi9
mfc4LGvY0mP5sF2+oVeak93vs1+tJz23khVm4epQAvBsSKVlM0RE6DgnTg28vb8nPNKK7FVJY/Iy
lP+GM6ciWERHMIQZ8J+BkoDq5PJpvY1N08cjUPWP0JOZdYHCuMb4ff3lwCq88blPYeg5DPyr/8Ul
Q7SNPqodCVzTg7pG9cALRwWJnkwS2Za6jTc9r/y6zOZo834rCV20N3OVcajhXuT65Gntg9sVViHI
IuHFXvGEAo/q986akcC98fAxdYRGkUr2T5Ep8IP/1BFAhKm5xOASiqZ63V1sTIDz/EoSrRcuSpwD
Jz1aE2ZBH50Soe30bWxuQtWIiCTs1W4gcaUKtyxlvKqX+SBuin0IB1D1zD+W4Y08DE/PKZnFXd8O
qv1nGKm02DjHD7wtL4EW6eKm64ZL9RUULnESW1mK2O4btCidPK8eZkfblmotnJ9ZUh9A1OqqO5C9
Ijs9f9vJQQXUFBKAQVwPKZ+nTTS+TxFxAMknL1GGWIeDi+nYXyOB6V3ScbTYWCPKakqrnZTYG06F
VUaZ/iewOUx88IfTyk4NhZcC/eRrguEGjKegUq52ULqP19Zs1WBUzA+DEtX/O4ovkb+ZNAX0UJvd
S4OENZXCOohB4N/MQWj9T6ViRi6ThkhG7ApETEHk4A1W/2otX12J0xkuy2YXuEbezVROUnp7WRTT
RU045P6RHnJy/xrWAFYiG/zsm1x757f37O5ZPqiJuNCkrCUOrmysBl7XsCSlsZJTD3Aqo/jJ9x/x
cADFMoUa9+QZ29Yi6hpu2xm4j0jN/QTi5Bpy/FJLGGmQ0x4O83jMPnALy8mYF6qiWk3N5sEgddME
64/p4qFID7OmNHAlv7q8EcmnsNJLP27L63D0rLQcJvjwUmyVxj1SWdp1LJ+XtTzS/HvgrWKjmvIa
CujIo6unQwjLWlgiJKQ/TntW7G6SUlI5+LiwW9EvO28KLI7vy/5gMD/pKXOt+oFOM0abEjju4Ikl
6r2SrOvG/Tr1Jv1b2fwLGJDC01QKM17OguoRJKsAD4pQnrwHfIxrCbWm+VmnB6HeOueWfA3of9Tt
jAOixcMb8exfre1akoTT+jAMlFRsmmuMauwz4fP+s4JsAg/o9g/Bcvo/ghyl8tsmXIQVk54dE64U
8QewPKqEHli7XjMXeIpoS9G/bLQ69GKhRtbmrRFD2WtJBe/sAY0LQ1RiG0E1+Bdr6H5qTvuUWqEi
FPTAfkdsVRIJHEWSVuUm1SpX86S476BENoNM8VwvLf9qxq550hu8BshzzZDK3UtAtzCwbibIhRaD
4RCxvTmxbjfJJQk7VGmVcQzKVw/GY7KhyEw/mYB5Jyfz8nbFX4XDbe71uztkj42ZD8XL7qTCxurp
X0CYUuFao+sL21eXpMTW0tok/zgf+/jfH8epW68wLp2KODgpgshyZc+9tUtdqTzX4+XQWBZj7KG8
jc4TRj9wR7hmrTGKnTp7UnLPV9Ty95jfxnQ94jtUvPW0vmWaAzb1b2W7eAO3e8LmRRUWRmnDC6mH
EWNmZ/CtcLyhEcXVwUjMVEX+Ome2HMoIkUk7r1QgajjZEuHh3xKqpTA2173cehIyEcBnSyVg+FNf
aBdLgxCcfMNJ1f+rFUnkP0a09HanyefbSJ0sBTMwaYQOicBBHRzGlzvbg/5YoCD1db2ZUG/TN36X
sWYXUGtPGZmn1VkiCZEhOBf0HhfWqX9U+5Ae14esIYOrsxl0Qv+pPLHtPEGHq87/tqzMK7/toK/z
Z903ZuQOD4InvKZQtqz+USeXJa3cSua3/cc6nV5DXDQZf+QzFOyMMF2NzAx9OrehCl+g2fo/4Mtt
mCRlgMGWMegICmnpT/NrisYQOvwQHIrGpnMOL6Zcip/lLQ1DQiIQHYPaCxpb2cbPwrx4zaRC+Vj3
WmQ5eHUZlm3V0/qVDaQzL/KxlzbY8JgpDt+UZI7mtNVzQOBdGotskP7JZLqngBfTLuH674OdGG4O
Tk4OYF6tIxZu5vL4bQZuZG9yAmdL0XTSD0MGI8mlbH2bthVUUpOBUneJUe3ClzdJUcU/0oG1QTmw
N4esNpSaNUo53rFmYt/pCga6MUQ9unDcsJzRFHnsrM3+z0/jfYLXyGmiGUkbklBqFZQnGzRSP1c2
4S3YR73y8CK/87jAfZ8wRA8ki/tqWNb4kd/j3NHtX+N0OzRapriAqDIIFyX+PQW66TZ9imFAR8kM
e1GCIekOWsYgFgbDVdRer8IDY+3D1qMbYDC8XHv+xYsrWG5X4SjQgJ9OsvnkgJ2Fo/rHLqhEzRvd
ztcK3UNd1LWoNLZJqDWBIeYwOJ99WeTWXPDAx1RAeRYj4lt+WjWJs0fKyTpwb/jGnzCnWxdxk8zq
M2S0doSm7krPBT1IckZ3RX6oT5W/M6feXzPwPpAn5MsgS48rH5CQnCTwwFLirVrnKyd2FVF0FPGv
eVHHh3yfhWUGNNFid63aHHpaoxGgEdTNwQGS8b4h4L9io2TDesNoteWhVeq7NfT+MdC2VJnQ++y6
met//HLXXVNTOoTXFMEkaqXZO6C9BNCYsl1OYc1I0tOB17eIWbw07bkI+OWMH+69+Y0urx3aObVg
VC70JZHtNeAsCVuTlVnLzI87ywx3qky6zDLQTumm3+78qfzP/5he3csAXbz8vvCbXQXFfCTqX4Us
7/j4klIeOj4ExUNX3ta1egRVB6BYh49FrrqgqSGhakylgjOBwiCHkBVaH0h/7WHS1dC5ConBTVGT
JtcXCwxtnjVVwX6L94Tcpq2LsgeoNuzbZxqyg9JDIqQT3BmrXL3dDsYi2pgiSGseIo5pOYuH8z+G
vVuzLGDkj7VWn2n0dP9Ou/vRIVdZdJ+dNQlcp5riF+/b31lqdrP9kBa1zhm5WhmRKoCDK6uPxSL1
TSPcdzhz+jhzLyNmNWKfzPHLccYeyNkLAqOgzT/k3IlCHCo9eG+Zowuf6x1u/BMKLVDvyPgsd0u0
VSrG4zQmmGMxdI1OJIxq5pSvEHyQL7XHRS8t9NLx9Hpz6XkfrMWsw1HY8xRnSqt+bMp55Q+NNLii
Du8x2iGCIpkYW/heyb+2wiqIZ7jw5w6u4m1H0/UBRhgOwCftFakU0NluykdtrxaQLz+YMIQQraKt
Nu2CRcLqdQGGdoyxdVdraPt1P0cXwqu3G+wnFEYn+ff0hANjZTU0VmTDLF8Miimm2QwujJuwIzJR
GNUrELGNNk+ppIyGaDggyecFyeCIqXb5K/r5dYm650kPb7zZ9MDcYGWbgpqqWQXYcO1U6IdrHBRO
um+d0rZGsEBxgWSHT63d5MOoINH6Axdk4bUtKVa/LS5Ep7YFbn8k8mXenB5XuIWHq+X5ccrSQQbJ
4X96ABsLDPMq0mGpsOXbpHoTwxUc7Vby39vbYWfn25P3rm3xuBLpp75mNU/HXGlk+dDWAXO8T65d
31jyCNUCR5/zE1io+EdzomWoqn7MzN23I6Qwsx+QfvMVUMH76FSpGbaqQJ5obKZnQCUWUx+eTRJ2
OgcArYQ5vgYX92L1Lnpy7myVbLmYRnccVlFd37RDAJKi0bcPoS/G9m4ChVvZpNEtyg2wLgt6SJwD
yzKA+Vc6EH7wuFVd2ya9v5EYAZlIWSeVydMJiBJ3EJ3BOdtEDymphbHUwfVDeX7tjeDlA4W8oQPZ
vYn0RRFZ2FXtUlh4JKf958Sa3oDFhDHVeeDni205CkJfC5Gsif8lPMLDnjl8iotoyM/JHxRZq0NP
5Zbjez0N0g/ZBwsvHteW/UJiwf8arvtOYtf5zjqJiZM+A3Vg3WTCXjzkQ7YqC+YalDvRJxN6mxPJ
L4QfKH2oaFGEJkPhH6+OzIakI46Gw8ZCIxEyqE6jYeNIOAGhy+qgpssfBUJHvQEQGjTaNSjYuepg
UfDrNJ9jCemgjReiBZcYLoO2mLMjxMI/zATHEeNKzEE/YuVZuIu801E72PEkfgAyEpDNM2Q7Zdoa
mMoiP+V6ZZznIDSQQ6sVfCgtUsSeYOtDrCFvuWhu/wC3puwRQjaOTjtc7Tuwrcp+4v5lvLZjITBL
7aUSHTphztQdXsBbp53j4Yfy45cFNOdHU3t6EeC1/Cx6IfXwRqI1t5bDbW/4NPk4HwTNaf5jGTB5
ZLpyqZByQecNBZPFIwGgzJG/cB9+xGr2qu4yGnH9iFwAxfBHpvWD5xf8naTbBfiz8NGsA9RStAUT
5VFHwcTMr/9IdTMuD5iscHdcqvSdTEEGsCCOmFeeP8c7FZc+MbAdWYZkmTiLPsQo9mjZnCIiNStI
jBVMOvC+16x63KFym+uCftV0Bx0DtFw1D8vm2VL+kobYZQXHLeSk1faspWp8bAcjnqNit+H2HYX1
5+ofQp2XN3AilAh6sfW6OlBzk/LOh893b85t9B3APAMGZz7BBxEPF9DIZP5UqHBg7LTVrx/EGtOW
ufwPN2wYE/QL4bjO3U0w7T0UPlKGSCWt0unfWpLguAhyPVnI4Xg8hXxIXHLkE5KtDNUmdUK0aTBj
mSuTsdT4yBmuwp6s9fsh0P5kC8oO1l3+HJcu4woG0vqw17SO1U5LTe6uN7KOVoF7TV5Ya3wU8dtI
3EKAgDPJPjYL0Vu4mh6kXb90pchWGxVvEApy0c2Plgktm+XiwovA9/VhuCSS2AEhwNOF2sKzUutr
c5MZKOANWWpz6ZaCH7OOLH5B/l885KPAEjXfqEBKD1B8irBe0flc6kiE2BN2PsessFhHQAW+a1Lw
ZbGYlksPf9hwYFY/StJjUh4ZyiH9m5MENSGiRL3rNFGGMMCgCYfB/pPI/EAaGcMl12M4oFwbBIZF
3IpnKqD91Vlks23UM4/pHKD9Hk+cicIT0FaPHTk1rp/DjuZYKxBHrMzHgB5lbw3bLqrLjhjYAFUp
PHGc8ur9GpxFT+Q7+MFLweIMhhFFQP6leYcR/9OOWypiISSy1CLVcL9JVn/mua82c0vGhHc0PhfI
u4Kfzg/Ug1vGRXWyQOD0dBKLeYlq0Wp8nuFUgBvsau4DHIqHbn9GjXcUI+hr6xsFtnJfsTA/EIa5
1c52P31KvwNFolnQk/Jruto26j0KxE5ZMDiW4JdI4rHMm7hqZlIz+yeuBVNv38lKojhqaDTwJXkv
/CtECHf26HwtZgG9h4Daq0iyyj/OAarCUbqq59EPbM/9ULru9u4wcKIUAJFSldwJF+CyyIuq3RJ7
nsW93v/K0UHdP1cpTJOroHrfMrIoEPahGz+/SKRxcpgzKp/Y+wG2ByGIO9zxPILrzxPAoExQ0HjJ
4LN1dc53tnAahQCzlFQywSw+NmyeutOfqg/GV40Gi3Bgv941AMhgAgGiV1qpeva8lGk/MnUg4kKF
bRPBf+ByxxoqzWNu+dgA5PMOGXFOmkL1bOGIk8kmEm2UHFVy/M0AtYGo/35Qy2Ll3uBPtETiFX5v
hUbAXEXvQjyCpK5bVecSY4ozSpb2vORsEnJNS7ChE44n6+HzMozhI+Eu4ldB1upY5RIToOwPQAtq
Prw1B5ox6jW1eSbQ/4lg/9Ru+i4PknY6yjeLXzHjTgx0KP9sTRNsy0AQ/QUKU2g90kxvAvtyb12g
OEbYmPd1dBXJBbA9bDNyWHw/vYBgKvythOr9t+C4bBSpaCVyLPtLvuZXE4k4ypYFV9k/qdRB1DUs
MnOAR2sFclt4f8XHXbYRYnOlhgOuvB8E48Q/4buJjaILkyOmgfqU6Ao/T9xWtsrkqni/L4+Dk1tJ
cWNqksYrbZN9QzCZkSRnjDOA11F8zh9LtIu90GjWTUt2X3WwcYj/JDgiqNZzVx3PbCotS0iaUSWQ
BUbJWKFSK1bTqeW+TL17uVtiu1LeXs3y0WlmOx/b7W2j6NlMNw/EhdpS7FqB7q5yd+C137njMh00
jI4s6IAn2MbRsnKElTS41b9hatsPjTYzaGoapp8kd2CTBmmGoZ8c2Nq7tOnRZA0goKLCBGLYixbu
FU2wCs6/YWfnV86l2n+CR5pw05L1//+YKtj2WICzaTGlNUuYHG9UeJj70CD3E6dCTqhbA4M+TMsx
1w/lQ2QEmJxfWrMHvaO9ZkJMJPkLCEye4QECGfecDpIQcjbS/2MfQVifoQZvCDYZ5hIG01tAU2eQ
haE7SK2hU3YVBKHHYtluMn8VLP0oUPGEe6mDEDC81rqrvUrJsO5EI0C4JipPmjhF5mNn/9PAPvNa
Mxt1mJuiKBmp4b4XvmfbVdVMUdjcz2qDnqqI1Af7pvCwqAvhDwk9jfEYlYt46MYZtQCnnOZmuGKW
Rr5SKahU0CTxd9AoC3JGYQFqNVI9b3s3Lb1fyZxZBkFlrRFhXDGH4d4ycG7QoasKZbasm3hbbcfX
TsqYpmT2csUUtPWUYkGh8gOJ1VeKJHKeWU0ZKM1LzU9CV/aQFuBnW+5wrxq1FQUDGAQsQYPIRTQa
0iP55fp6wWVkjhSQaT4CpfmiO+Gf2ygrJUqqweyQ7Y8GCoJIsjzYKuq7DM9lnSAdYvRs8+73nP+H
B7RirMqzqCXppNNKbthE/RFHtOUqml0Cn8J7yU+u5Uw/+4wx+katyBy0arbtl9mgwRRAct59ghsd
LpJgP3Dj6UW6WCx2VwG/9IBj4vhqvd2cCQZKReIahBS4AGFOEKQ586bh0KDeK2BgWEEvU2UKSC5g
3WD1f3Opu9689nz3oluTmdomXKmex0nXBHbayT7NXNkFF3sWxZtavIYhJwpbwrpyabm8/nZfZqP1
J8cpViYCZREFymxTqSO/RYSDeUz/+CI0alhzOL1EcDa9CFYHvWBHXYFMlNYNiQcw61X00rCevYUL
ivqS+exsziK+SKD4WFXbt9+6YbwAWJYIFSfysEliwbeQOplM0UNaR5upViTuAGG5s2Wf260TeW+V
s6eQr0TCa7LtVYqhUvtIBOfDI+ooKCkkf7c9hBCyTLmkovr4eAj0dL/wZwGe5txR2e/pqMINpJ6G
1oNB6yqpk9NI9CgU57XBZ9TJ/m+e5BB6qgDpWVPOE1g51cAPBBZsnjgQZfpw7wxXB2AWC6gRBef4
uR+NBwdtAB6Ris1riVFASey9juBjikuipWdz56nhyzw+mlAWkyxacIPjcN1iMXgopX+tAvaztkEA
Z8owy/wpSKbxsDWBzwg2iRWsshyLk9530VqtPYe3Kq6D6h8FgxkaXsCBzv+LJ46QyMXP65xVpo5Y
MJO0Olcc0IPGXeKi6wbVwCwc1c4ZEdcENiDIYEfX1YiInU6EW1y7RbUSWMdSoLE3XVeuc0M+qu0y
5rsJlQR20nd5KTMEAYHul1lTLE2PDauBbZJWFuLErAHRaeCZWXFGfag3t/gpaZBy6u783gTGbLbY
tBamjth3mePkbMjPIsLDdnu2oMVKgVTfJSXOy73dBpTwd755+ZbUPEnDxSD3lgZEU4KvaFEmRlmU
sKeV29id2gZZ2dRJpXSjViQPg41jYa2z4YJmVonO78Q8PKd3OCeIKjODl5CsfqdRVmhyLJQMZQKv
mLSlybGyM6Tpmukp3HdHmd5z8xeUpZJIA/MiXgRepOebkULKksDQxKPU20pvML9th0jp6FKCOWBG
I8gVzC2+YxzqlNFOxX1VgoHRflBcyYG6UeVr6jL9PttN0/hjmsV7RD3MN5j1g84IqAKNUtG9nTJb
OV3DVjOnuHaSCjBbV3L9tgI1XE/BYwzAdNVb9omYWbd8sB5JjytNVpwidFPVGWh/7+Uw1+/Gspj8
eWveEnhc+gsaR5Haf30xrlNj+/Dr0b3wQm4ER+jNgVWcYIOFHYgA39U3Sp1Vp9tUwWNNcHr42mRq
JDW6BqOHkmZNG19J3IM5FOK9bvDDrpsv/qEOpkYXxUBdM7J7mlFZ44i/s9ZuqlAelrzOQVx7DKGA
tNGRS+ES2bt7WM5BwWgDKH3WMhumY9N2otgy/wKROegQZYaFHrf60oKcUuOCaqlpiSri2p8t57Nr
lbKRlB6EfHizL1QDWzAEZ0gqf7p3XekGRVUv66QZ+70Myoqc46POwRFmxZRi+H+YuLktngiB13OT
axNWOVnTcytMYV8/22bXtB81HxYk963/Ll+fNQu7vlJOfixoq9EGO/OQALaIMjERabazramvJyoZ
Z9EnioEJ4R320uG3hfJeDTbHJb05HLkVUAQViixFlDWG1K0xLMurQ9bmUNedpu1gbO24vMhsNf9B
0vb0dh7stJ1rpZFCN2X2lHrUhQeXx8xdZHQvCilmNAxPa8whtjehbYYRhWL4jMJD5l6WFQWsoVnF
odnnYq+EjDbTXnZgXzWfop7PnahnhSqqOautssIw3I1JMQ3rxwPsNtKJqufNKhFQ+LVqJbYLMT/W
KL3kBhjIO0bw/l8atGHc1pYDJ3f9Oen8kb83TQj4wCSPxpR3iKAUCsBi1awyaVDEG7wlpoA29APt
Y3oEG0UdEeQCml5rQpgPVxU0dlIaL9XgzhYhlvikx74bIN6RU5ZVB2Mc/rIF9TMxM9ZZhpg8D969
Ne4p/zrutdyKBJU+ffGker9d955BZMyTWzw8iyb40rLtRRSlMzZoWEl6CDN0qQOfSy7DUYLkxuhz
2uEc2pDslltjv9lKCmQe+Y9wbrpzDelC2z1drwr8XZbmBYcAfcsFW9SC5tn4Y3P3hrX4PZ8mMhnZ
DdNSJgicm+maSkJkcIHXmxTV67ckN+Ndfxlegyb8cEhzit2xtMQ+15WSBBAqMXCtqY4dHqEv1R/M
AYXKAZNKGoEFWs+Z9YoA3FH36MqBXrhhQzdVf6dfWGa8bd+L7AAPr9leQAynWruHLag5kAzbDZT/
Q19hK1qL/QDbTIcYd0qS+I//3RaMCWNPYAJZjx8lJnYM1ysw2pdagH4iLtHDAittSjksMHZaFSyY
IxRlEp5pZTFrhFmIZsPPlji6+4YF2Hl6hWjDOubwKujtl3coHBA5EzvuUdMimkj0a5RQ11fD6BVp
rtxNooGzHMkKkFT0h7/9yhU/2erFL2cgRkx82KNv7ZGk/mW9f2Q7ogGHvxVFJ5W/jeBiiHmBBgc+
Gw54U63AjMmAYfyaFQ+I11O8Z1RYQhpIZWjcr6TfGbTb7EZst0DPii4oFtmrjRThF55NFiC4UBB9
Na7vhrGVcS1y/JSXqPEr/FjSlX2EwwEhjNnLeSYE49IUoCSCBi/dRseM0TCKp6JRQEHdpOL75mjZ
g8iUe2jipF4DLU66yWBCZ+LpKmcEZKrfjbTW7pHcihaODrsjuF7/zTe6AOSIHfYTgcSfsUXWQD45
pbM3508QfCbczScLSOLsIY9OB8y1UZRqT14ULqRRNbyHvIbVmBJIzQiEf50c+6/0ELkMgYr3aoNl
/EcVYK4NgXcZVtOAGq3POWEnmL6iuqQeROA5o39IJPCjuvKup2ZSptmS/lgsBBCr8z5A5m/Fn+2X
IfjgAX/rCc0H+vdgf0fCoCLMF7D5gRkNV1UxAC827czKII60kEtOyUDVpwWWYQ70fLVJw+JJKQTD
insZutOmcqM8q115wZ+0UfTDxpoAlJygrtcMjpiwaAZ7fiqbjIttG2sxpGaSBF3b9gHej8goZZdA
5zEJgnDhYDOgqvNAHdOjTApKAo0N7/hdsg5/+OSSgSGQRA5hXMUuSHLs5OWc/PsADzfohliEaORG
XxdK8WjTTzz+nWgGmIljxlQM7v6fPcYwqYm4871rqFk6/ug7c7kIgR0FDDcpG3OcTOREpXEL/ucE
vgc7hDHIWp7gc73FP+PpWqiZrvKJ5LSmkVKkV5T/PtVDXpj7dPygRgO3fI1vrfKF7rgcDiAZnbbA
8/bf3z0tNAD54zzILzUPH0Dhv6EIMNVpBIwOxw/E7jojh1E2Tbb1UbgsOfY4+P7rFoRqDp72z2ZE
XTR7hZ3SpO7bZE0B03jSqksvN0e3DprKrHxVwznOABWD9cXgm4rnzG3ago0QsGoEnaAnhDYO081n
6K0fVnWPI++IlhN9CQMX5QdkDRjt3yHKrTUKZPDMJhxlibfT+L82NDSIKgXGBA+SdSx6NAz4nxUy
4klx/0soEOtdNqu8tGOytPp1n8FfNBX9AMg2Ro9Mxp/MpzCX5PF0FiyKHcHWuuqxUHjgXaOTGG4y
bgEGzdHs2SlHdrK+/GE/ZnTmlfgkJwGlZzbWER4wPyQ3yp0UJpDWLtSAYOQI8T+6d7MHZDnTFrZP
GmXJSGw/WOhcR3sRJYV5aIz3D4ylivtg2VVAAxveLfRu/1grn7KTcPMf2grnub22M4qu163WewlM
qkZOG0+MWfSJFn/3K3WUfBRpaMJKGWiPqXvPAhugOrPQPdDg1cW2qe4wjUnie0VoLF0MZTvNRbGF
DINebkGQxvanMXxaiw8dt3ay7onqsEwxhbpRxYDex31mvgGYLeb1020Rguo/mD6xASXm0ytX5ijU
oKCZYPtrqsEh7NhRqhj+GQJle5A0yF+JueL2RPxlKx7pBtS5YzSveYMxuzUZFB1aiHHtyWANQW77
ex/W2N3gIbOWpLVZb3DRucsQ4+LBe3Vgz4h5+uuoZmh8CE7VzgDrNtMS7TTFyzNAEMKryoT6z/B1
qHyM30sxIxE4Hxj071DAzDT0HR2GFqURtGvyhp8jVS13NqNB569+Y5/JGqM77BJXHj/LtauDH7CB
gIaiVNXx++R8EoyGCZOP6cUC9CxGEG+ns1+7ImBQC5uN6koyWxsuCj0Hp83ewoSQ0aZrHCh4K0xm
I8ZqtvhiwMGXcgy07lrmDo2+q7X0wl9D2hBhwoTB6/U+mZ2RejG/1IsG/C4skbFvZRSYTdkOG5F6
T1G599PqtLqqpfLlX9vLY9gJi3ex/fQxAuzhm9471WiOwsjv92Odx7aCJIrvCEuTa3ZTm84Qlmug
jjD0hvm/xRwQinLM3xLAYys7NsBVKavRMEHYbgXx8gDH62w4NK4PxSaO/Yhk7AvT654TY03n326j
lvifE9EOKinhrp8iST8hVFcKIDpx5hrSTqSBrwqlx0Glz76BjP8O90PpxRXkenZAQr/uJiaePOh6
K2LwNfdNYl4FGU8NseU6dVY8zAiFpsZaS4WUmSs680LCwB7FXDk3HSodWJwiYDWm5psO40JLzYhA
oKOZPYCsyE1g8DV0zvI+rl9bCoHM473WOY3UYDHhg97LhtQ43ooK188VlCKcZ4XMoiXjUWjKKKar
r1uNM1FWFtW4EEOgA21rsYUA9sbxwlXWEWbEiX6X2cqbqE7GNmR+ykCOGuJJf7eUqMf6W/uEC3uc
+HJZAFjRpVjdKzb8WXdMQ5rB9SEGQF9L9ZVmZZWmBI3eFmWbVhQDYOARdvv6wKHxeFz4ore4lBxy
BUoQMyT0KpCJ/W3wMRSns+pxEb1m4cm8EUgyyQGorvQajAklC3yIB9uUhPBxNhxMCt2BAwSZ0x6s
YWbqiSfiBS9Pt+mnDtFiPBQZI9XVzTa3C9VD152pE153FjO5RgoN/DfviKPddyCao70oM6vTGcD1
JWLnWM1CcMZg27lRa8yHYXFJMRBT1qWRxjU9qJJr4oczfYTHbLqz5yY1yAvb4ADnupmHWR//K5e2
y9wbvAem3AoXHmHRKJVFvGJQBPLKXMkYDmuwYOXYm339MNvukq37QkvopbTVxxHRY3siEppzMhxT
m5+Pz70PsrSc37Q8qJInY2mWYGQhK/hSUqUZm0+Z/BTCxbUrqrZulsJCds6IwM/SuNa56SLIvJIC
wM3LJjwy/75whH/MlEAqkteQclLLH2AlihZbLaj+4HPeeiUXd9OK01BEcW8y9jv/tB7kveA6rjs9
WsaOvuxT6L+EPVvfUi/e5I/9nB5Nex6zExA3ZMXTHswNj3ciFdJjGXE2+c+0nDVbl0XKJDGz9rpw
avSXkPaFOei4tei77YFUP8vhb2eqttVnfIKifip4v+ZT1vVmIoNP5+Uq2HENcvEqQwIjLO4OK+xd
UK/PndBWZYWJ6E8amDNTzxzKU1ESHT+nEfOTvToxkdhWn3H+Psei1ugVvMKugVBxEhJ7aIz6wyiR
hZJgAKKtNiDA3FfBoSW+32Lbx78EbdL3FXMWFYJK2P4QsARvjmELvUOTGMQfdkzQrRbrz1CU25V0
F6eSY7tYjyiSq/ATYrvGL+YtWAAcolcBnePCtN4saH2XQJ4A5sdm0HR1mqFY9cn+ludhRLiKjvdU
J+WMU39m1kRRyq1u0gwVvNXhcsjgCpkTtfqZS7oF2AXGs27FTO0DWRmFWuMCODyDsCyq3UEuXcMg
g/s2SFY+rVQqVR+g9EOI7uFe4pJ5kthVLrpQ5r4fzjNFzXZyiOIw1Cj2dSIS3Yb2AsmIcrC9M0g0
A45CBclm7hisT302DOPPirBcuyzjmxUpSKrJCmUYYdh9hYWfllXfVAcK1AWuqdXOOl2gkmn2fDi8
435JOJRU+wQlbiklEWxI26VWNpxkWHoXI/azKYZxOo/2xbdWdGsEtm7mO6l7rYg/ieB3lWmgXOPE
oyew0Z7RsY+ifJ0jlsbj5Q78ef1BYiW4F1sRU9QY28bUHYJKgVZRz9aOl9uSIhVhFApWzgiQMUKG
O4Rl/FJAqmtbv0HNemdkKT2cqcgv1L4entp0Vz7JzuFFnkbABwq43PWTIdtfbhsuDMM1yC/JxxOa
8T98s66EHCkpswvGsRInA0sME/nhNa9XcFh2ugcqUd76Gulbil5aoAeRWHCes3XTbFs0SoWVRbm+
brgYyLp4nLfCRhftbOlBMxhsk9vppRw3l/cKq4nEajGPt8VGDegiMTOuqLy+eiFkSRWmA4C6R9bP
VbSZkTEtG1jVL/2dgL0GZJXR+a3FH6wsJDSJcQWTSnIzwlLM2m8LF/8FOIkeXXCbXG4WmRzM5ur3
FkFHV0HMx+HMod/TmOAqlgKhsqbzoJPOS8OKEVAq0Cv8pu2eCY95Rn7/woPefF5yjK5X2vLj+1FK
32WUKrfnxQzM1g14XNM7m6VOrDNOoZuQyrls35Hg869smx45K/G8pM9Iz/J609C0GySRzb6D/3zY
cyTjmyFlBHFGyv3JuueLNeKeTWYdSxLkdaNSoypbWviureAo9X1YB3MnSuIuG27ueEhYbgNujG3d
mWPjjTEVej17mJoaSaaAcw8qa1EsGzWavU2V1pBzPrIBJ1/9YS0ThBqiVzuLpVk7THvvCZP0hIju
7hMdltxDon7e2+e+ujZ+Bmidm9dcez/m1mRyp4vKP+toYB5aahdl3gK5v8PVnfuEneebHwRYgqpJ
em0D++MA4GcjJp+U7G55oKPr80wV8uVwyiO7bPzmm+8POUHhLbMrv6RAmgx79NbreEFwVWDZb8cu
VS6e+HBKBSUjrGHPA4CSr4xf/+AMd1QJPkHbuKOXa6lVC/JQ1BF+2xBZBUNJGVWNSwYaU9EBghRK
/JlWstWb2SvxsVi8L/5tpRL91Grz+ub7EiLqQ/ou3F/KLvwLTL6BziPR0ebeDXOuDUcUhMXBAoKH
qOemaVPhkBrs3lBFpCcF0UWxEOPNu9KmHqprM75t/sqQA8RefbMRPShCJ7pLBXRHTsULcOB1PGKe
AX+Z6sMYx1PRe0s6kw7qkyLp77mXTn6321LowcoVEcJOKdd1i+duIOXr1uDPYeKewwNDsKcHcFYD
owRkGS39tFC2fh26mWSnrvTGymZLuR8tBuqQFOgWGIVhMPfmivWkNUxr3uy/tceCnz9fEa6y5bce
BDNftHcNhBs58beQ/PAoUvsWWNpoXgBJvBD1cWettXpGr3l8qoj6UCzDAbKAeNdmyhEnFa7kN/R7
G3Kwq3CGs94YisjcDNizdXdDrYc8Vgp24z0i1JixZK/hyvlMcyO71OnD26TSRXi2olt48JvR0tJE
1F4unkW/n5oVQfCA+HXAhmuBShjTLx+dgpCU/7OQBPYMbsJCdIYk0zUg6t1i/LPxL+O5Cq+7yd5d
JENyr5AJt3yQXzpOTKZCdLnKQK81883jlS+LLB/Ex/gef7Kx7RVtN0RodH8MRGnn6KgqF2jWb17+
+rMnCbadtzd7vyduQnXOkaOzsmwIODvvimc1SkGTXqzHaAgEQIy2zltCPTLndKB76A4NRZj7pc9m
xt7Dvqxw1vuLjZx/C7OQxUrFOwuw5UHW+F96dwHZex2oa3Bv/cEt+sd3mCkllv7Bsx3NCidnnmBV
rUg0LPm6IHajLqSZvvmmDYAq5zfuH0IV8YHR7iAFb1PTiJy2fSi+MlK7d/Y4oOxTmsC46g1yHdXr
b2jX8F3lexyU5dc1OzelK508Lr/xm5FuMJACiVlQJXfQBveRYkm64lpwUXl8SOqE9xNELqRjG/C1
S4OCOqEYUEHUOlG1BngLiA1FjMwS9TqpbefYs0fTcT+U4BZynHhLS6CKQWGeNbWd55Kh0N214tyW
Ho8JGVl05xWaXfKYSmfhD7a9tQkkYG1HB6LDqUV9vbUC/2Z3BG/wFYDJSGiPfBJ9GHo6bmTTA6XR
U8T5+t+o+wgjuOLSvElnM+sS/ZOnqRR84i7DHoe6RFvJKxGlK1PCWsE54zGje7JSOcYwhvx1/Eoa
oOUdDjLvfNzAv0eeHQT2AoAhMM7nrQWwiF46qODQrxR0O/8C835rduRyfh46yXFV7PtnWPVacUiD
+NAsOa6uKNOMrHEst+MfhJzeQJW/vCGtiSfLCsi8HhjoMh8DkeWSqVWQAcJ8OI08OKQTUuZPG3SQ
Qux/ZEFNQq46cMOVIb7HITApyhJ7MnMw55J+960jjhPlvGB65fvUXr4y7xJ71jNFW8y3btywaXiV
/ajewGmVIINUzFftrIyO2ya82uPIfmsxe3sevijpzZsUXUh6NeYmSvO/YaAv/WmituxflAK+Ahl+
GMTJuJ3cQanb4saMHPYg/F0+o8U4r5PfjIymWFTPayonI1Q9mKCx+nxUuZCPOqTjnXrxFic4CQwG
Xnr3CXrOFkPwZXa9KtxF8wCIZP1EZ+DcEmhKQ+bVwp4luy+Hg14rIhF9+5SmCWNWwelxEKEynZfu
6t6lpge1fBaPzHy44LXNHGGvr18T50ddNKYZ3hPLf5CzPvscdCLRIdkHl0oGgVs3KCHi1E5GvdQ6
l5nKQZWDkdOU7e+9vSnKBtZWU/GrliJCOuEO8LqjT06PbTb/eyLR7tQlnBTXhl2p0k5RSoAXDORY
cW/DeAJiiP1chA2Z21dWxm+oBvnAI7xQRXvAZfSyFz6leU7bHpqmf/vglQWILZfeIBLbizdR9Z/o
/dVgUgMeFkyprF9r8sHu7g94EnlFsQ2xGhDX3AZuIStt5PZhBfpqwhZQcVFVYunEVIPehxVgM3ej
r42G6kQ+mSw+TLyv/SzCrwm/2ZKtBLrCD7TC7PVuTu/YNIcq4EtrRPmPfHioho7eAsK+OZ3aKAuV
HlUYOAS5yeW6mKmnfkY7xdagCN2iedGX5sKL/5cIaEb8msbYzCNYnmIclL6/Fl4jE+4ApCw8FO9c
waUPhB36F0giUgOUC70bHRgZJEY0naZDUjZvG/IaTRO3St+UhcNOj3ce0y/yuvUtN8RTLbcsDBau
vO6NRaxvthYZebUYRKqp+kGwq36JCC7/bfphMp2z2IKR5TOiqi3MtcXczPIeaIcJUDXEGLNPpwYS
goXsrR6vk7F/W11zvFxcueZftVF0Qz0YIBDNOE+TmbboL9pS9w60qFn4OnO7hm6OHpbN4p+w9PN0
nVkQdI5VHSGucXxpKGGoidtORT3cfvl7xVhNOrUOPrpSncCLPPyCJ9DjI3sRBbK/ILbaXnIfZa0Q
kjyo9u8mw6WC0rmiMkpdzkQFJfOEbzCQXmmfnpc3H6u3J2kP29nioZQCniqtXa5EBW2ogAHbW09X
qNsZYkY4rwqnrgOSV4ZV5Tvf356UDR3bEQJSjtSwrjtcSM69SxVhYoGXMm6lFTyeCT475Z+mco5u
3EkzTzY0DoxHXsEbfLr/9GF/NJIyVY4kQQi2mQ0kmw/XJLYv/9tHsbs/Re+qkZpLsC5LVMC39Yi7
k9CrU1OfQfKg5hyUiy9oAaCvKNJgzQt4Y/edg6nhC6ycoT2G2xoJ1csf7DRarf2ZkXcSPZL8226S
mw8qfWYod6qpO3d60XTn1NOmdcCTFQS6oim1XHZ0KGWI3Oml3xRMe0vI8gA/31KAUxm3Y0SY10s+
xbHnMXIsz3fn3UTioADJs6nNyhhJwo5nqd3R5N2QvkWDydOQNzfpN+azJgKTdEWmmNRPpEqgoNOC
JDHIVhd4F7aA41yLB2rzYIW75+pcdSQk9iLVVThgCOYY9k1E89kLGfWmj+Ry4EddlTdnThXziihm
fq6JIeaBloyPNPGWLMkkMXoCA7t+K/DZ1SWETDY9Cudh+BFqDv3Dk96o4lgimPLBUKD3EbVnIG4H
IOK+GqFezDy9kh4/CodEBE0Bq5ECzVaVVLMQ6aMJ9XjICG4HLgKijFeMor/pqX/jGF1uFaxQs42H
5R3oolsbAgTfpDg5NCnuAxXgdgpGtqc2Bzs/R+z7m+/oDkQdXkB1GbQBtAwHRR+xHcTuab4NC4nZ
cWBs6IOOAtNZXq7NBiU5drnyMhHBnNKwMEwYlu74pmTiWqL0aFnjVkDCa9W1NWwIdrujTe4U1LmP
ijepuDYwXe/WIDOOb54whKp8E5J2s/irqmqSOeoJXbz5j1UBdCmTxygcSn2y/AfqAWKDRuaFuWG1
1Oc1l7y1rgB3d8I/PBhY6j/IgmSOAm7d5jlk5kOUmc4HIQRaT0dlYaCfjL2xYABVtyLB35HsmeaE
McQqkQ2CNZphjENf0E92HLudULY0y3tNDZgbAyzrOWllHCz3vUSqeR/fhFvp7LIuAdOFHkTs1023
gxplRzAn0dbC+zfShrAHfdfV3HpNyqRGo5VFYyi+ZGobAhrKuXHanyUdgJFAyeB15+qKXhaAUl50
lCoRJ1mff+6CIP/uFqqgOVi4/Cmddb+9anuQ6MxEETmBldiPpGzIuxXK/ZliCzQ5W08ZVCCSv82n
OMMYHeshSORNVhK9GpsZiO5prKdQedJik6B8q3UxoyEVB4k4M0vaCGh6S7e27mo+5xCS6Sx7R6cM
7RPx/l3DOn/keQzZKt9VEEaL5oP9s+Xq1qEYzR2PLlxy5NsA7GXjyJ5CQYdiHhHe0fq09EQgKpYI
zWW1T/wDAATL/caN/Zn5AgMzMFM2ef+H39bBOrSetU/56FSZDJsP6RCCwMMtYkkIuKWQ9SVGg6wv
SYgrMBhTSZXogtfhTWHX6kckrs3bUgzhhSbbwGN8VWpQhueRSJq9OSRn59rZ8uDUNSlf0KvPt6Js
Ukp0QGX2D9as493tk8myqQ3HwuJxbOS5Ec74sOaJbY9Q+pb+vXdsHNQZImERiDadHBlCSkhLUUFJ
NAsR431YasohGzniDYK24Jun5O0qI2YCofjCT5r1XuWK+Q9JMCuGjXLTO4mGbvbbu3V89RO4UNzq
UTMYCQmhkZDlJN5AQm7z0fHuk/i0dp0MxWXSAfjaFYFlU5ml8a/9cWkI/kcot1OBTnQW9dpMzsL5
5UW0vvxlM+dhxjlHEXxgnGWWnzosFZWHJBt212ocGx8Gp4x/w5GUozHHqZjUvfD+EVJ7e/WtE4RB
gbx/KtCmMUAM7Ibr4DsoKWYv/WSZsNGohcSuJ9Tt1m2I5c8fg3jIrPZ1y5L+NJvFouPmMxNmGZQA
Po54xA+G7NgF5IOgDsLN13x25pGeXsQuI7uskVlMWOsrLXura/xjh4Ao5hXC7VK6+uKIEl2lMDus
OuZb8+P8C59sZpCl2peD5d6zoKHS6xaSDcG45XzctS15A27TPlGvY5tx3MmVTK0AlnxjEVGI41PY
vvLsw+DEMxuqub0B6LXfjzqfzd2an/wblnhO6KCCOm/+JryiePI/BUAZRmYDZq9tXw2AxY3KLToz
4FVtLzTKN+PkMTEBgihpc6foqUgGrkmREb8tPStjXtKOYvKzlmqAVE1Km8YdlBAKxGZrYRBDVRhm
rpE3JOTZtOAjwDiUw6M2OFGH3Fs2it1UYSuCi0968vXCcBGMY5tgQHkUoTlX9MORFaEUtJrHAXPO
OV2Ly2Qzyct1gY01nq939SKkbPI9Nqs4wIc77/B//s/zjbNFAmW9UTLyXlb3dDp5Q+FDFgE1nguO
EB85GCOxQGgk6XCgG8AWStIbh3f5rdjYsnyiGJdLi7lJaMaTEkTF7Xo+Ns1Tu2kq1I0YS7PXu502
IolGNDuKzcYnbqR/cf6B0w3J5R6M6olvD8vtmIj3yG2g4W7fKWj72YQxgmtskJkCPj/tKjIkSZTs
0u6vxXDYbaaornAZ87L6O4rgC6wWJhzeU9NREJAL90Fw0TqYXiuIyisRkbH2lsQnFB09cPE7fHdX
NVWz4vY37jryJfahzAbAUatYF4mbYJKRoRC5OwiVx0+CmUD9CyA5ekI5UpZyMwm6JErfoJrktS2U
0VubiCen5rqk9hve8MzBQSRgN/jxn5ZCkoJ2rX0Q2ADDfwx2ZfEtFr4ipNLL7wOKsyLBdY4HghB6
PBRpPJO3LuKrvVXVLhp2GAViTOD2Qck89bigcaIaVwStWOV/Tuy5nSXdygxw9wb5BGPmhwCNOIXc
idwAhgBFRkKomGukK+wCrSSKche2XYd6gwJDuJYOzajreD6UkthDHJnWHURRoshkP9+EMuki4wYr
IMSwbjPFz080QCBCFp8mSLGM+bSSgzZtufYfIuIX1WppbHH2CfD0Zt8Oxd03UWrGLft8fuueM5eZ
fs6FHBuyj4M9eh/dRLWlMv8aEaJiUxGUqv0SeQc3TWx54KgDNBgDUVDDU+fh1h4VH8Sda9IP7ho0
pZwfRQNeYZJr2aXfTyGZ5IfHTA1A160g3wLYtkraKgiqzz0WXb7mJOLSncn50OrOmQzr8YuYkuR2
13M+AynUijnxcDgAje8mOWedOaDaeqIw6ktRD8G96tT+j3bJ9G9pk7vsP86j0M0Ro8EZlUtSVLE3
8MvhBmObgiLLr6nm2YPKkKUoOE2CrNwvqlz3FZyrH30eKWSKP78LzMCBc8bqmBT7TFfpzrFnC7fT
WRoen8ok9d6EeTKyFnR2MS0At1n0vB1N6SjgWNdl7w7hgep8CY84UU83xCnJcPgachX6rNonbr39
0xBz8hxWmnhcNUEJYxZKUacfjzaDfLrzfE67SNOS0eKMZJVnS2FkWzpn4OXUZiGxK4XH/xm6eReJ
dPPmJLEU9BgC2NYz27Ck2HyZVY22/wzjJTdOG/Ua24+w8fU+ly1Vt4cjXxo+LcLcmq5siyjuRtVs
HG3cAM7Gg1q5+WlReX77hDc9vm7bajtyz2kTO+Gww8a529eeVTbG5wazuNAw8aLQDhnNmtZe0KJn
NDXcafbeAcuwhJJLNOAjyczusODdxZzchRToGBnl5e27rlwsTv+8c+pq81qI5Mcpy+UM1ySaj6mF
pXPKTRDr8k25TjkAxxuDTMWQdxKxRHi1gbiF6fQ9PtVAiDe1vLsTflnQv8Qedk2xUlnhFHrEp8te
vhJInyfSztBGWWORy6tL0G441cx02yFY9e0ttKrxvOfgffXaur4xC4FsSiiXrvafcBc9rpniKZVO
0tC8jyEXzLyveoUonMl5vatx5+zXt+d9qKZqu+5mCPMbRS62F1zNKB+Ry9cERSl6AKukJXINaqCn
EpomSR/44aO06BQl3Y4cm0DfQ0haMHBbEyUnRYmqULaOyNIKm22YMYnFo+14mcHYJUvYGyuabyIF
QiMnZKP0U9ozjLzj7Fy+8MDFM7df33L+PQ3VMkB9hmQwtjd8ed7j9Ma1XzF/vTBvKQueXYCsF4HM
AipRL+98zox2Zr0uXOaQa8/BSfN/vSHskhX8Gse+5KBYxc0yvVcMvQ+SmxvcDHn3vIv30dVCAuBD
cF869RrRGkxFP9Vy+zbga4a1fXJ11NJvG3Em+mkpATGLu88rJT26sPP7TTdjO1ft35bktWNQFl6n
BvTHDzG3Ysy08pym6kBxksCWuZNVBnPuWrmFKFdKIF5cD+GHkO+Rt9ZJKMD0fZAYVoOOwzjNNF58
VfkwPmgT5Cb/Y+fyZpil6c5FdG8AaipLCfTEJ8ZnpcTS1na0myPyuJn9xo4fzZfInMxeSRmFAc42
GdxoFTFiROn+s1U7jjPO3HoTGfQZyIXSeVOBn9PB3zbECNOFCsJ9lAzQRnzf3kaVy1vYoCx1jp7T
44DEHIKF0FKXkgEcO2DsMpiKxn7dqsRNgcX33zpOIwWLoldAUE4yI7YmPliJ6P2Kh3sodEwJWW6G
64HojxH1SoFfE98sHzpEuZOUvyXP+eI1jNgm0S9T/SW7Z68ItXij5QkprU25U+GJ1eIhpdVEW6XZ
gP+QGWGtbpLAwCM2+lNTE/3MF8JD9Xi4E3GVhbN6oOB6sAdkCctGL40S6e+c8cvmUBvbnrYmaA0z
5O5Z3dpRugAmxhC4DIcUnzJkW4qRnno8N8Djy/6q5PVaTEb4Lvv5vrRpyAoxPWZagfZ4WcBnreQA
5ezebH6X2M1smUS+uj1i0PjOV5P0LF3sXFdtmZ59XC//YEQgP78OfNW2Jk2fCn0sLUlo1zXiT6A4
XG4tC6xG/8wtikokhfcqQz8W3Yox9vtLuNUJT+jpl6tp7mfPLJYhn+k9VpsLGt/S+aHyN053XlRL
WD3vPYa4Ix5g9XiHUU75T8tbcJw6QzvRogh6Bg4uE0XFtHtWEveMIgSv8ZzdHyVtOSRW02TOYIlI
QS5iuebJf2zxP7ptVbJg7lcceq2vMhKB2LHuDgQypdyTpKRA0U4KxriNJeSy9qzq1ToxCGTJakE+
b7F3BvZdZj/8CMd83HLLP/kkZAl33cV+n0lItkzFNaIizg303sSijnX8TdyD3wK7u0GOMqrVfftS
+vIax3AvQHuHxhmHsMYX+MDO3I+MfMqT56oXnOE+pKcAx0yoHIsLIK2/femjnVEhPIsteccbv0Xr
X6eoNeA/20lu4o23S1SaZelHzbtbURAjHysYieN0LHeTRZzr2uAxOQabWCdyWNY3OW1r4ir/MYpq
WJWMhNuu8UZ6WZSY1yZmU/HupmStd74yQd63Gh/TY+n14CrRo8txNKjOWQv63Hp4vxJSk+4HWkIf
nqnUDorlxcc0qVIUB7URYE//h6Too9LGEe8LMnNIfKTxOzQ0klqxnM+6ASVb6FWJyKbwvquwYnR/
sHIl6H7Cwp07zZPTEGEkdlCz3sbHjS5n8RjWyCdXI256F1IiskwKwkgPDK4VXSP8ns+Lg28XwLem
5JiRart9BsB6QL48xfjtZcxpxXaasknJbj8JckH2gom26Gjs1ilYc0uaggS7lVL5ObblPvlZnoPQ
8EQVTJUKfJEEMzguAEvFusRD9oXYMJNs0V5RkMZ0HWzr0NkbHZ5aeAA+7zbgU24XaW/sZafyYmP8
R/dEBpyD1wJURTa6wnrEEbuqJo98l1da2iTexWJ5EYPnGw6c6hyfs7tzeov+DqzjwWU7PFSKzJNQ
3LANd38Vokp1yZPPQXgRQ/yzV6o/B6ylTdyOEYQzCFl0HshTdIiEUYEh6VNveGK9sMVDPQ4XWIfR
mZ5Wa43cQbhpqe3rGAaxyIynvAY/oHu93b/GDEXl8KDmPULBhzuFA3mZMSUlL7dmaRy8nvOrjG6x
3mB6LJdfTs/ZX58PEGnY3HWPm/Rb57ZoNfIx124VYyxNEG+lU+8gBRymxQ6O4MB2alv7kmLg7n8A
wXT0x/PYj8e35C8CMEsFPJOIhRBNaFshiCU+5Cv84zunF7j2awC1OjVAYDeAUGI+dExDgz6NiWUq
qYVXYv9tA3Qu2HO51SnujAyw+qQd1YvHOIqgOFspEwSC+YVkl6CwR8aGoUmsxfxtu5UV0SN+xftU
TwxZpZhT8BEM11fJf+3qR8nXXB8OewTJNvKIerq2ZTB7Qu/MTIji50CIYKVLFZBUerXUujuSwuFR
nTv92h1gWeIfok8t2412Dez0gC/SiMtzIG47qneo5OJwlScMWfHtulc7bZtzsaga+grabMlESlnL
/Ym2oYPv4VtbipUkWOyUFnVaPdwHTDgPv58FRZULzshqD+K0jqyMUKw9XIDiWTCrK0qU73mXLllW
WUSwSzt0DewPluI0kDFDmVGBgjSbGcmiZUJOIIPWoou1ZcteQx4y8Y5pXptSfvGiehZAazUiLaQN
4Jz3LdKByXlCkuHHjE1m6n1ssCjxLSz9ocEpP7DDZ7nJubB/K2Zas9n4MnanFy3frr86MOrGzNpp
D041iBnjRgxM8o06lPNF97xLSvUePp4j9GrPTBoUK6bg1MkbalhTLjQhESsoN04Z/s7v5W+6Ra3d
RC8NttFOonft9sfKdIbyrh/QzYm7ei8H1/h0SXekHc0MxhA7SmVjtdeHrd+AmQyI7lOiO5tqTZ5d
1QuCKseK9+ulK4xq0Qyj5nDzCH6FzxGTvKSGDK53tOyKHv40r7kUWGk5Eb1SS54LsD9dnITZ+UT0
YLw5GpRpD+c1g7zveiVb0d6gXFfn4YBSLjrQVZtnwmN1cD/O+ZlaI4A1qOdQlXE84DJ/RtuX7tAu
bxm0K2/NO91A+NmIzG88bQwZB7z35M22SUXLmKcOinSl14wImSMrRCRRwyyZ/K/F8/MXu+GP1YaQ
4/XC227P8uwxPG+NpVdrw5X9M7zhtDyd0TcKct78svg4pV9fItkxCfkibmUHV/1V8KEDP9k59u4r
bXH7sMkH35rBJH86CAk/Xmi00qRSAGCQCmw6IUujOMlx4QGsuI5oGNcV5u2JOElUgJHSYIc/oQol
3q9tFO/iZ7Kzn/ul8gfpo2pqALCm8m+mmrpsK0WwvHU8/p9oio4P33PKkIXLzauP7buF3MHeZOuT
6lw06u4kNbatal+6w4BGL+dQBVn8VcHILZpCiETWlts1lDz5QBlPMfMUEsRKpDRvJ/dnw14noh02
sbeLsDTyM9+gkoeifMA5Ot+E0/WVb3nZv/LrVwBb03WnFiho3cv/ucIrZxjrkobZSVr/XADzXGj3
3N5P6UWITh6LJ8apiChxJ9YP3EsjSajMKNEQpdMTjCkYaJMrh1qs++Nl1rEf8Y1qa6J42qbljFZA
wl7p/h4F4UpLKIoFuOXaalV0GDqQgobp4nKTxAvrlRjjzj+JnAEgLIBxdj71OwAZjJAhlFErlWMP
jXWunH3hiUan67Ae+WAwdaIAcTuLWbXhSi+Rtgbw0ZlIkyhyo1dSgxOpEpADQgSTg2whdSsitzx9
ecErntguKl5ZyD1FgSAZ2vW5Ch79EX6Em6cBuzovz0q72WAfnYb1TkLWVDckDAkwykG3qrMJhnvn
dMQy1Ko/2t21PK1CeldzxDjLOqlybJDEzpKLPkp+3vUYjpPTWOr0XtmGRvtZdZv+y3/tFu/5riRl
G9CzLknyFg9sw+XiFnaI4JEw0wkfpYLi6eGL4SGvHYy2YGi/T3G2actGwkmMZ0lYXqqifHmec3Ge
Oss78cOKny1JGoXLDHeEwusVt47y3IcVSDOL0tV/rLpjTo97BVnyNudzwOii2tAi3AnZ4NpS0rcQ
CH7ZrpHoUoqKiraYL808Cb0KSxZDQT+AWoAp1CUGfjLhO/vNUgSgxHNXk6zJk0Hn3TdisBsWhKBo
J8F3j1vH2SSWiJqANwxXbqh+MKQN8jqxD04Ce1UDu+8K8nhMwY3zrMXKWBfOaNevN9Wr3gsdi1Ww
DocwEbMpdb0oebUJ8WjbwXbnNH4j3uNgAMpiZSqhWqj3Y2hQWrZd78vgLAfC7/oslQYy5Mvi2vcx
Gvm3NI8WeAGi3DzO1nMsJQ3ez3w3jEV7m7/tSq7TeeDLKQ5P6SPRfyK/i1NuMWmgDngmNZ8XaVz8
gpXb6PLvDuqhbJSmN19SJDWnLLXBTblJv51lCmkuAMIFj2ErVScQ5P8pERKp9r62BKEPvVeyj0Ff
wa+Td9vp4chwmc2h1/UI+XOdR0VrNligw+BnyE/QBPeOUS6b+MaePAtiq7ZGhe2wasD/PMnUo0ff
PlSehAOSZ6ZQiIV7qfSKI94PkJrgAjma3xJmXAQhs61yfiKbxST0Tlw7NyG6IRlELDvm09S39BoN
vAaOcfT3AtOvpOgXrXpYjiSd75B323hP0jGBy/pvFjBjXQDV4HIMf0yynwoogWAWrBevxmzBcvdx
NJ/gzukKVTaQWTE5+PLJbRshrccNoA0px1VWqOFqwjOgUjs4lYdIZO4TTI1XWVa4DOcDoQOhv8qm
y+UkDWmDTqj+xv5ESrfGlkmq4SY2QDx/ALUZT00V5psO7d2/KxKljACl9CPkUdYywBTgkfQj5cT4
Gpjuv9yhh3ypbB8Hinno/anfmMY8ZYUliB+YdkZsL6OTT8+thRkyvA31sgEtAlkpVzOa4x5JDMVG
J79WKaaBB43LWOF2JLlitJ3mupZCraft15bm9/yOLUZjJQjj+BFR2GG27riUhWmqCDUnjQ530bjn
XfQc84c9y7HhBJp3pa4pE4UNBt46lzr0qqZXX8KvrtwKJFcBf/gELqACeNRcKtXh+0Kh7DVSPgzO
bPQwft51edWHdJObk7KOsLgrr+9HdVSDGGy5kdneSUBrev13bl7K10RAIzQtGz1kCSYL0O/+01kb
l9ZsVPRVC37lKosviIISgDqhjL49e/SHwJipiQU22gLFyKe5YQ9X1DHBbuGiVgR2og5uf8231W5c
/YvEBcc0rQh5xHhxsCqpjB2/SVQJsvLjPHWrxrV+oXICCCCxQx+dIiOUCRLY7gz69ROCSgXFR/sx
lh4bl/bq/G9yK3AvfphCUpK5FbWyigI4k1NjLuIRUwqKM6hbpAB+bmTF42jFf/WoVxmsGRq3BBmC
qq1NOmxzzmqH5nHvIl+A/tef0xTcfoL4EPBhkLBKHUDJ8WxHRedhuHbdmNiOP8TqZJIurEeOg1WI
kizDF15y6+mAMH3haOCWiNWyDFN7Xn861SDGCi/Gt5oityYjZrBzYNXczSZlSwiRnknIuEIrK7pF
37fV33LvYkv0VusjC97HcSnN0tMu+Hehuv+PXt15abGY39GuXPiNHMUXL1haEMVd3+614dUvcqo8
DEGjLbxBT64Uqz6S499c9Yra0BZuyKRuoGPUI1IJvYEscpq/EfTkbBJ05IFmiarWT0mYClArgqur
HMTgTfW+NNPa+JTIKQs+xT1NmYNbJKO80CYRmwLyPM4os1Q1yFNDnSs4AjlhE364d+GL8lQYM/pq
QxiRqfJntt+KIDGFCBMDFDDN2H50DBvU+qJQq8HAP4mFvLV048hm3g3nJQG40/uUILAZCiDwKA0i
87TbolhA738Wi27civwqRHsxxa/RusGP9j213JFaDtHuyysuh8IHKdfGuDliJpba/giVMVzbomYk
GvsP0FgSfu+FI0IoYuWaH/4LiN2hjYLyps4oKx3QKh0oq/O98iLo8aOZynPCMxfd2rEzeqGzPgN+
T23c/AbDfslv09mp3oJTko8FX7LgICSsM4qub1NfZMxLnayD+6XuszxDieosddasGoTPmbeUkA2z
uHCvAlsETaK5IzFDTV4rtQpQYV5A2ErWlInNimTPGKsDffLt5ss13nTZi8aFJ46myX8cuaFV3E3W
TeMADtHYorEryZ50MrfRGZPTQYn+cHuNv8x2mg/8FwK9NBOZuePj3IroG1DIOLTKiL84uPUogOBX
cSVvR/DFSbLWRbMPN7JRYKgtnlnOyAyMmzJvsJpHebV26aYp28MrMsLaf22s3uEGosvJGsZ80XKo
CTvZA2eEHgWEz4OTwRrbPooVjMZd/osiTc4wKqCn6DqdxRiFwDvlGQlAXH9MVnNcX2oXQslzsuhT
9yyYew0sH4A5BfT2Ja/azVPLWWizWpc4shp6jJWAS2aJfrBVF8s8lTFG9jQqn9SvNpQkmwIPJP4u
mDQEHHfr7gQ0+3f8hH2tUEp5H0P1EeGUZCuokvqvV6lwpkR1AUIuYE8f8lvDVjHaP7G29m+Tkd0Y
BaKDoYLlyV6rG+RjYE+0rX4vV4Ex5Wl9732GfHslU5Gs5xjjuIu5y7qrPMDBpALgEbXpTCqs6KMu
BNhBm/TO2E6Y8mn9qeZvizaFSMX0cX9X+2XAiZi1qza+yyrW2k7JFMdA3LiTTG6RWgEqahYvBmVI
XJZYD3GIShnRXPdzzQnnb7uWg+I3k2+LOsNd6IF+Xd5Z4Dg5KwUmR+hk7e1xO6QRJ296ZY6jvWv+
KUHoF8b8DfPv/SkVirjII2YlA+F+SdjmRVFjeChQZ5a1WbDlqFhDnwG4++8z173Hyhpv3pFbKKhU
DvtOIzyYz1EalIampFsqhbbBIF7OGNP5kyesAjD9cR73RMTTKY1+BIO/IhGU4M4Ny4pdtxSem/rB
CoDvU9oeZQu2sXNFb8YBYBDDOYTZdMrzIqumTxBlFnzzDjRKUoFM5sbRzwmsIxv0PwItv0lrLvF8
J792ww0BM/QPhbRA5+tw7yUiU/79tJCkW9IW2ZpUc2bfhfw+yoo/LTYldxrj813IQf1zFE2QvVXo
iEIDxYSbUiahUvM4279F8qR/jDcEhUIZF3d9DEjzCajCFGzLXSIME7faRLVw7BMoGhOaMsMWh6Ee
S43NGgA1ax3nBai5XeXBfG1oCXfUEw2mA+RXL3ylo1Ten6B8UWi4rejX11wXOkidT/7DzEkP3Smf
pK1wDX9P9pMJX3iGoEP7Q7+ifMKBY0EF8UUVZ6ZqH16yvRaHirpqXz2UzX0EGaUBaltmVjD03206
Phe6hl79GXD/DGJP0a/4ZJwSsBlaSpdRRtdOZADNDHOfH0m9EPrMIBJ8bY99lB3BZOCbUe1JsaBT
XHs+qxxpTBqonECqF9G6+L6PptIpVdp4HwqveUsTiEBzb+avyU7FGuhj85Hkc1Ux8HA5ttrKCp+E
ohCOWVb0xkFc6/0RncGdHJNnsgpLwy96yVbi7J+/vdZVcIloOy5eKYyawOwkMtMMz470vRa0gt4s
ku12KAzwwgbStxtMoXJKqWEaKO4k+GK6aNzVZVYerrGVRyEyvqalVNyjgjIK5IzbeXsuu7jLwFuG
tM7hjVfLXTD4IAcEawZZkkQNWeRVxS2kxj7HqgmQ5A3llpJh6hOGK1zUFh+uNt5jh9/050s611dB
RQmufqDdAPGJtZJq7mYxMQBiaaw/WEzhwAvxY8aSQWg6/VHOMYc0vJS7tsJoKwFkmaN7kikYRySL
0iaQ2BXasHyazT2p3ZZgx200N9fENZD0nRtzTm/I7+sFgquptLWsVrn5lYr07snuQ61Y0P8NcdBD
QZO5zrhCFVHWO+HLUZCNZjJ+umzqquTh2oKyOjlBulthOy3AQzAb2M26Ax3i8/I8wAxRp5EPB1ES
k6zLmLpELIs57e9eFKnFYOlAYT0GIxxmoQhZeQ8MKViYp9eCjyT+ooyt5/OtYfThuA+8C/Ybb7nw
Y0f/WTgQ1c1gRwH8UQ+5EC9ybJr8hCZo20xuhFosJnvg2EiMj7kWl2UyctyPPyKz99HDJGd7OW2w
5N2bk96svxMXR7qVbhOu2ZVgmikQvxSZHMxPMzEtABy+4HXxJ87GiyJjKvZbWIDbd/qapDgTg30b
GmJ7G4YRTsVjAX84lC9xuuxgU8ehUbIHP4cF8EINsfiaJRmDS/haDxx4EuVRV7H82bQGxlEEmwvi
XNtkIsDi8uF2qq1w5tTrzepe/Z4UMLVFvg8+tKqatE+ZHn/7NGY0BS/X/er5iQ7dJLsqQlmV0kAf
1PPWEZp8Be+3wzh2EckUCKXFLWlptQ7H/ExhnNP5YE1guhFRrOGMamJm6i5O1UEKuerFcERcR0aK
galHMHtvePFhcfdGDTi5QvgadkmgYBKH2Lh7QUwaOP8Jdm8zUkeLOH/ibAYJCf2eHU+fxjNW+8YN
JIvYKPTGz7CNUxIGhXunCHE/Uw7xVYK9toSZP9ZT2CkDtCSMIb10H6yXS0WjO8HUqkjT/6O9VYs8
+04RhnpNumZu5jsh9t1CJSEyXwWX6KEDq5b0PkKjv4/C5Hq/GpvdhX3eobF1ciYGr9AnuCc+tgtv
fQin7xQ9wrbw7maFIrD7YNDenTrQr2Sw6iSKavBDPej+dC25DP1zu7/Zj68MlU9c8oGdgxTTT3Uh
kGWMrlSXNK/jJdFTtUv11X/Xq3JwILGvQDLSqKpmYom21gDIj9ZzahFWpkaC31vmjyjwsz7d+nAm
h8mWP9MDa8Lr+NLSQAQchdsDKr2bjMYz9Z3GGI9+c7Sa6RQ7mnX5buSvV1nZXD7vDnVbEF/+Pw5F
Yd107GqQ3RqRw13646TNbM2QV5x+SROihWrfgUGMyqIhXCc7h/T8FFVn8XMmvEfLR0097Oc3EFwh
R9FbhSI+dfLutLkXW+CgQ+HW79e7qOgYl2/0Odl5TlyLymnLXBAAEgWVJZAL48lDfb5gC/l1g8oR
WC71zYUW7XO/tx78CZiyn1nZ6xoHNL8+27NcsayrhFJi9wm1QRCCzyOirgpb3nvbYUJJvTWJBiqI
LLQ8cho5Fk5LthaOXYl/HI2q+u/frCHlSANdUCE0mUnsWHPpV0lMIOWHv3rgVwl44D3OZX73z//T
tBBCGDxSzbsQbDhao8Fw/qNWZz19c3viDD+N+2BCIdhafyqKE10WR2h8Mf9Fwdt/l+Lkx7et0xKS
QOi7eaa2wQnDmJJFTR9BrgJ2WD8XEjhm85fnt/e/GzQL1fnpwyTyRXvXZ2ILrXyznr/nvXC00Cab
1VhiOCEalb/UY4HKIsf0dgtZwxUTXzQV1BAAWZpyHXtrv/fUA2RLWfNfiQ+2ER/8HViam22dHiVD
uyRls6lZCCNF8UBh3DgDNXiV2q2V66SinD1H2cbAAmTNjWH1684HtSCpM+Mn7bbERTnJRwgcLWkA
bfcAw2TWBKJeDcSBqE5gN/+p5RgCaMDR1sKT1yT2TZQAXa3jTna4ObhwQTeBYE+AlXSGSyiagvdI
T5NZrYf9FFssroKjFepBWvJED8ImQS/feyNy1D9w9uCpNLL0ieRAdQDqdcFNP+GnAnhthItwNkb1
km+YdVsdfiumEpCJxAblk4kRCE/d4L/9imlutKjiwIG3w7YiiLXLCdD4FpAgHfIXl+paeEpNMKBK
cGmHie8XYZmWdkAVER1bu7+NB6QZ8Izo+5Xq5t1GHFMD76uTuYfWNcv4WyRp+I72QIzsF6MDMJVh
XJ2m1+f2nrUpHarfblDR0J/yZJ5X254bqVVNMrbgAqUfI+qoEF9WPHgc4YM5DdgBD9hzpnf4GTdk
LKjt80xy2ywn2hHNAro5ZI2CXubLEj1EC5CKIkadSaQYYJy1JmwYDD6UnDpP71/Rxw1rAemQCSWc
peTbzJjvDLSHm5O534SSgAY9Dcq85AAwzrg2yQzqCx3Pk4sEzhAw3oEShzLXoyHgW2BSveWfH0c1
qg+zuyuFoZO7SkJvGGtgTMHXt29xaJa4s8l+T2gpFCFGCj6jP49vWwZ8Wiy41PweVoPS80/6CLQT
B51nH0KX0PSOUbhmHRBmCWkup3/Nf8Lm7vRhRCIbnOCKT3+SGwVFAiRleKRPuN6a89TBzEJohjaW
QYBJkNB0oYxI5ISCUYOoz0J1+bbghxkmVzh0V2R+i5zqM9eaR7CbyVCwsXwXkb32XyylzB74slQo
xjr/3UxDBBgyLJ2VbEs8kcGZQNfCu1sbR5KrpXpcRWxHdtqV/naUJ64/gDj+tz3muZW/Xypo/0Bl
9WZ9Bzq7B8kE5H3KekuN+DfXPgYGz5TblRakvnHPeeJrEFJ/hUbauhVHUwWLZ+IPurkWg42MfZ5A
j0/OfBIspIdv9P4/pQ5dujRAoQGoxFF7Z1v8hbp9xBluzzvboQSHVmbjQ2Gg+1oXKK8eBUlTke0B
5Se8whClUXc/8R+dyEnqLEaKcbFj125em/0c1G7QJyjnsTYIPaGYKjmJoWHBxERRhPVF3RhDeBZD
/s3hxIPJkidp6BGnL5rZGh9B4tewed3M8RtttBCin6vQyDkPzR1ymfh1P4Nnk2hwXyQ8tXGnmlok
JjFBdKFPexE63g+0BNiQMXJIvs8Z9P+601SsbLXGLVea3mtShgRjsXzikrG6SnHhAQYG02sYjFF1
x8/Uc8cZ4/LqBVlhdhIuWGNUBmvy2W5y8fjxVWIIgBcdByCup/5R3D9oTYzdif6hkguFyQA1uWxS
m1ar/XkLoFTx5Sp//CWKx8mNWn4J1M3a1DRGxPODQv0eubnTLP0TkEDrCH08LZslzX1WEIcoQjPv
P5pWRroN9petoQwQh8zLZsdNf+IWJxAgfofxZVViJV7JhBng5gMu9tgm0KdOrq+/TIB9v0V+Z+/a
mp8oTZ977Zy03j0dxCBsnNmzk4UnFXzEKI+sFhUwkGRP5ieWKTpCxthTNtNCHqxxntXdk9dHIeQz
04osbiSZNXNtZhK1b22iWZ/sbaBTp//mZN01md3DNmy3UKrz0fkgEnEM00uqBx8s1VBbUtBb0iLy
4Mqmn/7kGEgc6AfYeTLcfQ21cROZXyYNtCxpWNBq5AkmIIl5dMJKORBU+JuehNRCh2NzrTKZCZ8w
Uz7D6d+a3dueiYHm9V9omrgE68ElZPq7iFv3IWgiJ0dSVox+oiZKz/Vd9/m8fXSvWUIn/jhRllP3
bZSNW4zePqfA8mhJ1bezGxob9JBJMqNaQsAQcS4W38Vft+cDXUT7/XK7qRe93eP7n5bu3bpdwDg3
c2274d5svjcnl14tPUPJj7ZRLqUgMrh9npQsqPou5Z5An5tukInkOWDvEXfd1YcSIbVfTBEvF/Az
UAgBoNErm7CR8Wdq45oIk2GUsapAExdFtu+DZEPdc4Jq/V98K8o6tK69X1yDKG4hlmDdex0UQCtk
ILF5tiWsm1rPLBkH4PRRzOBZAcZSBuUbsZwj1kY7nrAAjMsZUDa9zlQ93jh8Zyj5juGXdmhmuQPF
3pt59adFsw/zXvtBHHshJGJj+GDNClp+NbCRz+xIFiR6A8WJXe2UDhVBZ0uLqkr4oO/kUIQXk8wa
dAtPIHhzBmu54r3sRwkWWDdoTip54vBdY0YDkDXYi0qv2ScJFw02dOGnJFGAKCVa/HUJgwpRrzk4
H5ahkASgWAYHyEOZEaW9uLM4wpjTLeTOrbeC6S9hzLUK7Mi81lBTXreHm5GSIv1b7U8aFyckYcAB
iyWEClKS5G1XaLrHv+a/vnPjC13KOyzeAX7uJxR5jt+MJOT98HMc/Bx2TdbmAnE3a+2D+agzlRYP
y/zyqV3aLTVcTFiznMmrlqUHOY/ZKZ8+onUsVFwZSyr/iNRVlJfzk/wvT1i/JS4wOiPWR23l4asO
Yo7retDS1zwAUTOGHA2wkScIPi71Rnz70/sfzCKIqY8LV9hrGhfOghfjwm2/uZKJKl9p4RREcu8K
GzeQXC8TeMmj0z+q6jyiNGidG/9WDubKc9eKNTkfVwBI0mynnaoi0Oc8MoE8za73jx4mzqXW6FS3
B6hp8BsAPZq73oAnTs8j+KjpMQbJribHepLiScLYxqbvd7Dq264MUVfGJWiKKDcQ31P9HCzLTnzK
16YVITSL7TRErvwm7xZLmk80YEUYkTF0e+BS/KDjQa0t/Q9KGJFtBQaEV/Oz3QqCIN9g7jqdKSsN
Z/Prvba/PWFPvHeojbaVBKnSd57ZprROe4NvIcK8pJzr6zrhg2/MDCOlPa4BVdViGBXnd48MzdKc
lm6mJNquEGUmaE26LIhsFhWzm0NbCF1BvMEF53tDZ+8heXT8zLznh1xUBjjzrqC6bcHXfAJ0AdSU
GHGKjnfITmHbjFqXkJIz/c3wd8tj4ZcNloAoLLe8cNuWfFHcNjEjdrMTcIrE6XBFHoxq8ltSdRHA
nnLtQNuE5Sh3kTsVudjV3vZXXI+nrq7rk3Lw9lNGdWhLmly7CBcmsH3NPYvlm2EO7PFvuBv7dXda
ev3A0xSKXR9flYveAv5rlbYm9Ud5zwE293Z4zf1fx2/qWVSPRN3iqH/JVS054j8JZhBLJiXcO8lj
hd+7Q+NhyY39A2kGqaC8Vos98mOFbNnZV0Eh7TWqsOO4FLY1Nn7Ajp/QYngt6poyHHvwtPNBMh3s
RmJAenuV1A7rCxf9CZH1FHzAreboGYrLAl/8k35FEYem//G0FBUUs0sjPcTWOZ5yOFmXp71vJOPl
0Gega56V7/n49pgiTgvGjr27M0HnPTho8MzLupsSeSEaVlKRHAGd9qkpor8GO6Jg1Iy51ErOLYo0
NhL7VIK7Fklypap8ikh7ZU188Rcf1yhpURzpwGNdTt2yyP4WQ2ioZ3ek2h7vCm0fU0ggOJkBEo9z
s3YA3E6VFlKelS7w5ej/FivNl2r4eqDAcFYOAzCJiTQjDYjGZaujlzakXwOPx5WoXms0LyvbeuTO
Xck3i3kGg5VXm70BuS0WkNxBLvr2ft3KMRJi9ACpuY5T/nccrOPKBQC+cGAUktXhXpHpHEDQWKK3
sg+2ASh9k7c9TKnI45yPP+OWzOLQYhI+47jeEmp8gSMAesZE40OAuFW5N7ndVTyl6DqQDG/pdIi1
bP9Wv2hSKjaBIFMDJdo0rGY7PlcQTo78ghGCMoy1lepAx6G5np7KkL9gcSANExMEM3zX0O6bIVTS
y3tZib9dIeFh1uN/bzoIABNJEjjGtFuqJ2SgVvR6broYFvmddjrgSh1d6BZNLGQrWwwzbxz8wVxB
dBvcXewjq3mVN9GmuCrC0lXNNRO4AoRY5SFg8VNF7u7a/XsiL3Yr/cB1aSKnMu1qo03FM7HJ904P
XbA7PhKDlRnBXqDJ2xTB3kORY8X7KTK6XaU4HZQorX6r3BbtSH5PxHDqyi9G+X7g9A/D22UAt5Fd
zg5vI84L4TWeQUtQDu2Sukkpvs+aIGTYmiIrnXzAuYNZKHU30hGC2oiFXMOaBrGgUFA0Fzwq6sAh
pfnNbu9GBFzUpIW4nut2fJTeJeA/KRf7IZNtWXla+jIJ/Fk2eMq2pnsrd5ZYq8lAFlQI84WWYGAr
O2aDjD9vyUS6dG875hmnqYuzn0vedyz1gX1iGltGJni0C2KdTpido8JZSJZ9Md7IwDoQwnbDQA0K
Q+sW1x9FJ4ecyRalc6rkKApsvYiX2y2L6eDP6tAiz7cfcQbwg67gy3Qj79AeXy5kmHPr/wSxW/We
IFyua31+sUsHUvK2yiY9H9qHkTtk2OXDtF8aqk1H/40lgAPxY5H+Dc/+K9NFHWnd7mV+SjmDek48
sE+cVlfNCMcoC8bszR/5+zBvXKTUaLAnI92LY2Jjno9F7oZE+eiJ7e7MtW5tVvAhxdg6jVO2cSik
pkt+IiIpt5qTx3lleO2WoXJXWMnhdEm3dWZEOByqaMs7s8cPzonM7uohOblG58VFHBbglBYofTVS
6ynfXA1UG5Iln03UjDCPIC/eRSmC8tk9GMGk9yV4hICa5sZPF0iUP7jmABG9V81FJ2LrOzbCoQfe
1MJcLeKIZ+x1Irp0S3mo9d7LKkFU6X272Hfe1tPJSIWaiaNFIHo5FZvlDF0wgvHNrJTpj5oeGa7k
FyxSeV8vntAiTapyoyx8hFHd9EBEBGaEBmFdo4i0ytph3wqnFDUQcX8gx4eVS07csAh0qs8WOZZT
QUMOp+3TJ6iAPwMDccjHQYz1gIY11H2vPr1yuhNu/cctBG0XIWh3gRlTBXJUPKZAaZtdrRFxvGXD
lji2u1p7L7SKyy6tqogcoGlZvUvBEXi+bkqh7o3z4Kmwz14MwU6D7Zq/n00bAT5+QH3UQIkCZuUD
GNl++fBS5gDBTkBYr+hAVL6aqa0GBfCX8/1Fc8cKz1cWUfgkmC20mbrAgWKKt/ucb2tqm7TnfRkH
jTYcl+lOZG4A9s0g9bXeqQilZwdVGiIwSzXLRc/jejuQD7UM4iXyHO7sY/qSjwOgpYp6w5uZOiz7
cwkpGVI0AXo4Ac5LOouCtFao9nshAXA03CoRoQKRDJA4ylx2UoPSWbq2YnlvPEx+XuULSkNtETX6
MxbFRmiD9cAu0DHffB5iA4+1FMSbP4m4sMo/GQivWzVn3/iW/8euNRLJNBRBH1fEZ3F2IIb0aOZO
GuRjkOP5NxAtEA+I9apXcwySZevb6x3lAPNQk8PRaKH9L1kVxN55H1ja+yR/wXMATlq9k71KWuRM
7O4Xtz6quKXh9075i7yx934+BnbvaIkPDX4xOp4LVSv1BkI4lqodBn2THqK5Nv6sldVIXWMdmS/N
TYBQX9IWgO+GPLW0raderaDn6AL55AWc1mZo6bnvwqJkIMkQjEOGEh17g47h/4DyJ0VaVA/TmA64
GeAhurHrWdv0UyFoPiF1QiHjwd71YFv8WIqPw7tJ1yAQFm5bhV7w8b9j0z2xQYzFpjTdh8kBjAmi
wl8jfFO8QjIGZDD+6PBZ4lfIzn1eA8/aEIrP5pgJ/JxaiJqlV+YT+GWroz0BcMuwwZXoubiQ6mrP
UU7DdxZNpP9rHI/Rcen0PfIUyeWQw2izmamlgK/7jaoDMa2QwSsTQkI6IuQYJxUwvYNpmWAH/w3N
3ISopuLMd1HBxpOoDpHWoFV4Qgi3nmnZMdSMcKS+H+GwnKTwJbfHl7jaruH/1qONJ8Z2AONARwne
eHwFIvKDtwl4AFcWWex4Mqyewqr5OlutOZ758RX4Uh80jOKx4JUuqR7N28WLEXMtKg3gGS0faFm7
l4Jbu/bRXMmxYfjKTh1IQLxLjMImy8kSc/4MQ50HwsMdRk/xAfkLyfXDbYrYMPFeCJakbTGD8N7S
nThzFU0A98/R11EBwx228J0exeOFNWXyliWzWBHza8x+hnzcJdR+2kCCT2Hr5GgM2ogrzuNwefpa
UARmb8Vud5PSAZiWrvkfBc++3bmN64VBRDQIshXAmR6dOZ3Z5oujgTA5TWaTAsY81zASsK/a7hEf
c577oSEUYOiNXn1aIPvtqYfWEOyDFajwg+bxi1046ZVruT1pPWghsNAYkV1pEwHxywiQyd2AY8am
+g+jyO/iQM+tzNNGz+Z/Z4XJO/OV+VwRexQcgsO2l2fIfZBr4z8VzglCk9V5x6lEL8oSL88UIY7p
7TEPce22G9Ajh2vlw32dzT/JyneRRQBMCUKwkwUofeLWVH19F7JF0/MnpDhh3vntyqwr7NsZ3JYA
/GNhlyXMY28UgzWMqcvfagrXJY1FA1uJzGGKTYJ3YbQf1KHFBExIXj6ewNEGXxmb8X92FmhDkz7U
3BSmSE4vGyXuExBo7G2SKwz/BoWq+iJoiyoEPIeyY2r2A7OQySYRWujmvC5uY7/3XvI44mr63WC0
It8k84Y9I0RvJCQhtdaUzP/qYLKCge8gIUc5DsgK0g0Mk0xy/xvVdGVhMVQJHN5Kl5xxGRXJwXti
OQYPHrh4OsrI14VhTQgsHzq89PIawrS4/gJv+EKdXa9n0EyjEa6b9KiA27PZBOiWmg05SfT1cM6W
mBBPRX7pW4Lwe/yj4dJjzgXRIvFj4VD3oyy/aIBk03wpvxAgg1OSAzpQUGSyrqytU/XSWP8AayPf
dJxb/enhGQvkMacG26XP8Oyoskgk5m62vrFiTiEQf9w6JekzAVt9j8qbJirJxn9lCDdtn2LGoEYs
6Thk1FZem5ehDF6jimRpka5pUcb89D/5hMPzjS35CsWae0v3zYlslc+v2ScCfa9aNZQsdIXVxobf
s/hYNd1h3RNqb1BXLJfJ1F5e7awX9a3v6EwFFM6oNe/XSO2N2h78b3PcxT9baFa5Uk3ZakiZpAQP
XG314H693matEWAhfC4uJ+KBFIANoy6Ty8DdIOp2q3MzzfcU8bjVeHaY93UJ/2/M5b+SZUgr2Sf3
Ab02iQ3oi+DJMCkmq8iHQ3A+j7RK67qRUVwOS4J9FJgixo38z5j0jFsv0G0luqWGzJNVGcOFBO78
wvRG34Cf2+bR4Mq2Djr+lo1VlNBfyjcVaafaHldU7BjCKmeeVjBs0LdOXb+IojaWYLVx1Y1fz7wF
TJPNJEhBmCBC36Hji9IuvCnuk+q6wL5aUXuqTmIzXdaKutkw9t/gj0cogMbCOODMlIYc5dUim5SA
yu5+bAZQjmoGyNnql51Z9B31wg+s/3+z7jjYGVjVOCtPUYVjN51iWd6PYWSWkEAKM6+nQ2u36eID
BAz/cU1VwCSoXLCAgEAXHfP7XEDd3MeKNLgMkFFz65nmuhAIDDJ342GRo5GZbpSUyiFYfU6rmw1N
2+sp2OODZQ8HXOKrwzKFA4AZC7vjssZTPbFqaSXNHZYL9iyEeovl0fUL+jHZCks92DfYMxs/8eTq
1J9VL0LzSN0btfRFWWHyp9G7naU01MxbqGEuAo4eUEO9ae55ahq1M+xwMzk8dMaFjFuKV2Ka9viw
/WDJtkUK9lvKt+DRoeLEJqSGZjUoHANo/oK6i8Qb8IMSeEG0IECIenZqWUipX8GnV7YK3pFmcrCA
DtbyvhuvO4OGuuNw5dfRhyxBtYCt8A5AjYJLRGjzScLDvHDZUD4WekqHNFwUKcrrXULGXPatHpIo
RbCS725gqAY66OGKF1yXkA4y4BwdKLG310ffmLVvNtJ1t7gT4NqLyqS8YEFo8rAdyb3lFAqWLXoC
qlEqqdXQxUiyFrY3Es7AiZ0Y1yXKWCcZgCS6bVm9+SpWqWPKBPtLGY8ol4aE4tF29KO1QuqpzNME
KUyGFw7T7tRRJwQhAZ0WRGaehJw1MpATD1TzmFKSewOCQO0d3oEeBLn3s4qquAjEmp+PJCve79aT
YozSUA1TUwE6p5T65N6ji/f8jhGpdyWZ0HK/rQiToqKFKU3amHciZtfQZBQ+roSaV0LphhnYzF8m
cOvr81FUzvl1oN1dRE/lBUkeZiILWUJw49CqnYAblGk2vKiYI5hG/UtVwNRDnSPzYEe5o3pA+b0u
RExMFpaeXzOGD7EEEjUaZJsnov8+xKJ7ZuTSkurE6BBhhuDFadt8KKE2N+szYqCQILe3fSOJne0Q
YxkMJ4lFKIuNIusk/xlg1wAuh5N9Jqg4hEfFSHnTqzgWCbFrJCBO6dfhGbANy4GjZvYhKTVq3deE
g1ZaMYSUnJWoDkyOGOkLIJ5gb6gg3BtcctL/95JrjJCjFz3YDjqWfha0n7N9B75yYn/y19oJhhDh
RZLBOO5PwNGY8Tm0me42ljNKVwImqdGfHgs1Bzsntvaz4OCaaS/3HEXyJ8HK7cZgYupdOdCcZJTw
EZrNnlC6ShVGJDX/ZuOmIbB5K6uAyVq7SmXBzyD13nu1cPRREhFMnjViDXlA4X14EpzB5RoFlxJw
w+9OnlWM6+vCt6xuPfQneu5mryW90sN3SsPdoQerA9vTb9xMnmmrj+ksCTwsQE9a+EkWGWzvjsRB
SNqK1YM1S1257crOUD3a9kO4W5r6cx28wyU6FxBVPPrs9oDLafKqHW5J7Eq9Qm6cmVhVDnhhVVKA
Txk5+PqLBClOIBJFbu3/NloJsa21uOgnnkw455BBd65FDk9cveuj0dWY26ehGxBhJjhcAkg+Vf86
Fad0DIfjCcHw491riHYU47mmX8gEIiFavD1XT133SpimuBNlJ3vxG82Ah31erTXfNALlTx9jRJbe
cmLJx4unsh+/TTNZjEqdL1le6fZgIqgI51u8ZY9E+EAeME5B74RUDK6R9mVx3hLh5LrkfxLhV0Fk
4E0IGo+y0tDje5Sq+svyli2V6LPDPvqLrqa+a6AGgmmYa637vvhETEVXE6pXOFZxd7jnGwPpRJwa
jPcu+UI4OvkXflBRgDc7WPsKf1VDLTCkYFt+c7+KIV91HemxRXViQQaY4V0goCNR+2Sts9OWDNV0
I1xOWJ7yyGuT+ihUVNUdBnbUMqgsQw6fm8S4/gEk4AHylV6HEM9wHCzkT/o7cOf8nZn1veneqEoG
OJ57uFh4LRK7iMp10DHtkmd3l4dK8Jskx7U9vmtMQxIk1OGX9IkXUYP+WW8yGjMoz22pR4umTKgg
2zO27j2BD+tgWTO0HG/iB/0omC+MV+Guk/Yl7YCXiASH8OtYB9w8ILx+7QDuNsQbjqKIIIYMRdjL
J22Tu8ABrCmrQDbdCgQM/Rra1c3N2mM5j5/mwsCB2cgJj8CZEKvbSUxgV5h0pKbawhZaOteLVZuw
XSlonXdQrAgXX2HOZyELMxhC/by7C7bp6i1Vl/QxE73dDkXyxBcMSkwXMHaNCRe6IN3xt614DdAT
Fd0aIDzW7GqeLdUum8T4zlTGdWK2v+xoyvP2+wR3egXgHiW7RlQgplwrrGC4al3M5a8gWzreDh6Z
hJSBqV5/AoMLHbueqn3m9bc/e3o3ywoDD/0okJ+3FZeaX8SyDfgwCVUBhbM+c0/BcvOuced/9fEL
xB3B5i8tddXTbr9JeHdFk024jKq5VNVqt3ctdIamUfKJdEjJBnz1TOuRzfGvC1k2+e8Um4Hef+S6
uxUc3fpz8zR1TRFs4M3jV0ePUKX/is9ulghmWEUAj8hPceMfTwUsaa61XdDIpsuQ4JMumtgXUSkj
TXAU++AZV5Y6Ii86VuAHJsflpn+EDDOvCQApLapagzoPT1RvUFyuPqa4+RELn4aaNDq1SuT3yGXG
aXOtDyLmkTzh31/xxFfPENt3NDnemRVYAuEPh7OhQBeG9ApzuZfeaQdJysOzsKGiJSupu5tYpkRB
xagmeFjbcyatGqm+HemeX2aw2PDTOFG9TLjrFIn5Lg6TloRaUQCfNtZcBCJgOUVHK2gycpUnV4V2
9DI6NyDzvlpCiwbH5d2Qj2382YMxZfUBzNeng+RvAluWAtuVFvYhpIQUOWXgMzE9w7siXFE3PgYK
egEFNfTce2DSnJsPfcPf6SzEsFTLzpBjmLpkQgcEGtBsIMXD9qvScCzciojXKRNE3CH/JlxS4iJ1
gkHLU49ZWbnE9jHrT89Fopj4nRikRZB1PuKGf6CG066iYp5vQ5wrGqcaGURmIIn/y6KCDOI9WVU0
y3ZzfgbGRVnB1mx8sMVpaHVBiI8wDCDzb1U3S9uY/yxL7jO+MYy9iD1NU1ka88j45Su0GBfohLXl
DOFO3eCW9yY8EeWfHOgUg/Zuzg3n3S+VONG/dEJZ7P5gMBbsg2JNzhs/mPxYeqxZ33QzqC/p5gm3
lUWJeFsIJqztOd7KPaNQ+QCavSiYioo7lkkvgxbya1NV/OG93X6O1HUuh9OOsyZxsynoomLx/Z8a
Wz3QGGxkeZwKjP1eNqm6Js9FhvhnRjTVOSDfL1y4h0ZtSQWaXxHTnTyQHDkLNr9fPcZi5poI6I3i
SLYS/07F9HARtrvT1bV548Fl09rBNzy/Pz0oOHX4jOK4iB18nn2QALLiqTnRn4Z9nnCr5LCSHrsr
ljQzd9U+CV8YSoHl4fpfaM4BR6ZLHD08kfeMksH45MBvYZ9B8IK7+n7udgRPz4ZzDoch82U49CtD
gLE7dfemErLEzC1n7FvAo2YkOJmm1OKcjbPbFHxncjZxEhkP0q70mHrgvRhNMCW3TGfMEvMGBvt0
VI0ObjfJ0z7EnYmsv71S07gx2KfW3/XzdDpayX0o3P/ZAJulzANn3ZJPpQZcOBsOvBwPelrQ8LNM
v8dLCjH5d1HxhwDFX7xNcLmO8OuxQ8gv5ZchkKOlE8asd890myzZozyPiFhr5aydwF/7H6GbMOWm
Gzu8t3++C3RFvfggpUGLDSLuBITO4K2iSrBY9DyXEDjtMmozPMXKwLmPZCfDlWWn2RCxAmmlDiul
9c5ZxWBrtUXutRu2KnlntN7lXLcgXcjHefGSbRuCg0UN2SxzQn3UZ1f0ejALfQSbD8U4swmuoD2p
msHKuCnP0S50m0veJ1dlmeu3ZJgouneIJeMhf9dC9R/MC3q5f/uFqOHgqcdrY27L3cCTd7lqqFVV
pfi6RFKmPxM4gIOttK5ViXOGb/T0fIR/dJoKBkrVXERS9N7AVVbhpSC4C8TzPkCPl2jQon0ED29I
39BTzBML0Po9TADd8jxdvGRM/nShHaz0BGN1Q70dxZuevJ7t6MkauF0mIlHtbgo32AruFBxwFVRf
wiFQd7QYYzR8AencXKAjzQlaXszkXDhPbvH/1o6hqLjdhmITmNYEyS750z/Lndd6XiqlZeQU1VJD
0kNG6eihChgmGq9k8R/aurTLgGNRiJ44Ztr7sVpGpbRaLvCP0YK64g+lOaNQbx29ItlOJbTatNW5
gjrlbIA27Mgf7pByjL6c8piDyTAKCLNvac9BeoAVGWE6PMGtjg5psm3DOgJ54EKhvCK/LABGlAJM
ZTmg0gHpavVuOvCAB8ogB3CgGEfL94U5Y4HuNfR5VMz3lBTH2vNzrHxRU5vp/v7mqINrHM/yH7tE
DDlc3sQvTHSYi3i+TLP50jaDzbfvw7BKRL6hNAKTrxiQ6hJ0cfW8S7bt60p/N0yTGDzdKRcBrKKF
qDC+gVcOqdLbxVSX4K9rP3GvEEAFtqgTUfSp0FGZH/gnEixBdKDljWtywF9o6VLFn+YufPgbEJMM
g2R/ZuwdbBWan4zgOA6uH8unnMCJKDLG0Dwa+8F7KwfhbBk/O4r5JRdjnxRjKwLCzfKwVK9UBryA
Kwi73RuEEUwRUYq3e9t2rXW+cxle3ufjU7M/wfYTYCtYewxp4pm6PY2XDCHdaNVu09j3xjkRXv3g
xt+aK/E3Ec4iHmkbiJUx4V9Ggaoc/nH7k42SDnc9p7mPAYRAmPocC1mvyo/DW8GC1rL1tj+mfXq4
USdBdJ2OJ/N54GBQ7tepqe84ngjqEMljTlsm//c6mP853OZFg3kGC6448GUW2FT/ys9OR5Gy/R3l
Kx67OMK/4RfFRsR1dQagbBjjziM7jETVZXPUYRm4j3IwfVuwFzO9uS2/HDDQ/RETbIIC71q2R12M
NA2Q6vjmhuvgheMxYIbWVylPGhk0SDaArP0cLCYYRCclebvx3c/jnXHmtghfSNSZIgmOUcfbMMwm
EmQkGanyu1twxemunnRs3wd/GTUEYHEU0ax5tF0eJGM0T4U52ffSYDPn/c1etQR8gs+jdOR13P58
if7tnHr+pyhUKs02i/7ahJhNLwFAZMRSiCAvkaJaWrCz5VIideq6O1+jlxycZzqhOjXJgC6oK8vM
gDoJIdbVsyUXMXr5paupR01G1yp4sZlAsWOosxxRVvVB+tsOnjIUMbtkQDrQhWVvTaFId4NeEcGm
0U4F2ew81a82Tw3+bp5n3/sjpSR9jcKX9qjJFpYCjnFQ/WLqZOfmurkkWcpDrYe0MKgDgSOxRuYI
Y7ez52c/Q1u/HnVqdkLRc/e7uo/Cj6UM+skKrYGU4wknMQEFMPO31TGQ3lMSsPLigYUHwWQhZdYx
/iIOy7Q4KXoL48Ywg7tbWTBzv8ff+l8MRp+AI2zIiVH5MjOJDfyEi9Z0VTKv5bqdkrWn8P2HginQ
aBxRVLxxKsU5WMvdi15RAtlRGzduZymFZ8ymRnL2pOlwfK0eufSv4abDwqjunX0CU2QI+5WW1iX+
xAAwC+QNY5z9Wc4EaV3eIBntJ4XjUX6SLxNgkdtWu98U0iqJC9/GOdQVRy42/uqEG9hl53fa2qI8
bGu/fV8XjAzAk+DcE5w+GcrA5tlKU9MtOnuLzTJ1mTUVrX5gBWg0lJLHrpyRH0P2bFW8AEeFQGqh
i8Mtkp+xTIZHFDdCt+z+cDt57sMTb57sTk5IPae7ASwZT9m++pmNsjZC5E4CCXY0Qz1UfvceS9Bb
Zw8XL3XQOU431zvgyxhfB3vPjj2AUmUCJbh0oN5YYJkP/x65Qa+Ac6Ex7PplyVyleOUFpE+MOWWz
i+mxTZHrZOt5/o075UUONXxb3OoNvN1KqbuPaMZTAqxQbnHh/KjXaIevMjDium9gcjpIbupncikR
Q+NxehgkUTXa3ltPG8dLNr9IJhvZpZQhscaw0tBWeDDN1/+LcvToz2/y9GND4MM6+4F56VofQCY/
xDA82F1z5xnSZoCcbKQ29a496hfanEtJXvTN3ik0Jbuc1W9bJNcVXa3o3Kwh4/3Xz0oYesCNnpLI
f6ua4+UWLICTl6lpZqOF5Uds/LAu9fNp3yXXEkvJaatj7YPx6OffWMdSg0AYl0DYROM4gi2W4UEn
J4gWeJyzdIXJh3wyu8eMJJGmsWyXY92ju6VWUy2lOK5S5150bLXURRtHiS/dYUnfKQinm9SLEijc
CMjnWzyfHdxsNo/lzt11RrvFXCUDil9oWj5IsoOe48ouk948C6XxEB72jTRhyrIHsthoajzL7lII
s+FgXm/TQ5aPgM0bplUNFRTKdY9Ojh08DtcIj5KYjvxQvxYkXK39kk2J4pQs6HXcq+OVRrWRnRDC
EkCuU+yo6HzmMd1mW7BPjY2NWZ5Rhc8fOdT5MrFQ1cEzwbEWc7TEAcZp5YeINJNDmOmL5LR+GyaS
zWLoCQbmAoMWxRAcN9noxMIAsXN9Y0h4niddu8+c6z1fkHZWbmW+fjK5R4d3rxHVFBVKuz0/iusm
zqwTqwl+uLgOkVN0KF8vLWuhkKdaIZaAQ8xCSzbcWXEuItpPi0Y7yhbF97ovt9xKDRYTpSZf23/k
zipnuF1Y0gDfMuTDF/CW9A0Fsos2mv/vNgzlNweSkMnddeiD9P7Qy7JI5z/1FbupdAmx0Mu5vLUz
5XtYcsjv56ADalQs2MeshR/+jFpWIGjehIj+FqHgO2mBxAhDvroTmpfT4+tXuSY6NcHH651+BZio
Z89ym04LXnQNuShJBby+SPLyAizoOUGsgWWHyRfaB1/RD3IkiOvJQmh6H2KsjCwxQbYb3Y3cYFLx
5CVNy/BG//O28QLxF6txnjDvfxSKamRFH5G2ZVC5yPhhhQNQWMRbinFJpG3IYg4JNb+/sShpQIDK
3sJVhcWicKZT7bpqeqIPiyZP4CmCzKF7VnJSmNbbA4jlNZRosTU5O9Lxe+lvcKDbApsm6IEP58EI
tv7TJ0eXtXcKip9SEJOMoQDKOz6/nvBB5achLLX71SG54CnIh50pc5ugkmx9tBHvhojQh3xY99gZ
+WNY4mfg23SyNmJ2QHpGePMclUH3DiyCkGhxTUdUMYD196DIP4bcvS8MoEPisRwqkz0FHJvDb5W6
y0kodKwOQq11smdlppuvp2Tx3Ih/pVec9nbrY5MWEAAO6rEnem8VICd/BY4hzQeqqomT24ZNXoqW
6uNIusGAqUW1BoprgXVEC2Nt35Dp3TRVRanli8pCQ5/iT25n5YV/c+IBqm6tU8qU0a6m6xIfsB1Z
nHqYNfME4Q8mTbG105G1kA4chYs18MhrxZ7iAWeektKzl7XFYEpryeB3kTJcv9oOHr0lAH7IHmg9
LReN+NAV392dHawhWihOVrnVyTB1tBJgRKP0lwemXg0d7ic7bLRMAPQ+4mktyMPXI7HSt2V+6DT+
dKFptcVcsOseH9sC780N6iZ9BxLt3Bi4ISDBuWaCfSTWUk1lVuo8GdadlH8T6v0i/fAdDNolN4Te
9mVmwJvavfjn0/eXa/OmIjrBCugmalLiqm0BQZYTq7jih48SYXjcRBfSrw1a3UbDbkFc7BeoHNLI
nFSm3deIzQD9BfaOcnFrnIBCuAa0a9NJdmjJGiz3kjpTss3IW/tye3xqFau1Jp8sRYKr0LjTtPTd
oKpyWf6okjpkzshlIIFgzTpY0fJjcua1DTE9jpqGoxgJZ3+njsTpFlVlV6DfLOpRtVQnDvvsvfpA
IlRiYxpYdUULw4IB0SWNkwNSoIgSPqruODAaHOJrv9EgUJoTp6xKiYwUQ5gmTD8yLoiI1AZpYeSi
V6PA/yn0TdYOSMe10lN3BDF5ImLyOSppHogRsWih7noT4nF2/1jlkZ9pKxJe52urwcD3EvVwgLGX
pg5M1UNA5ZTP0qGyIwEaXeToyCUJo7sb8ammozrSL+RoLVOwj3HdEgQYp0NNtNUj80DHew2+NiyB
j+3ke0KJgF347wkhWw7IpJVBGvtklkA/XRizIyY2L/8Z2kg5rOAJQ/EJPIybZqIE+7rv297d87Dt
MNtLCPwC+yOMe1be5VAlBo9xGda5Fd7k6WPUf64GLVw5LJAEs0rxCOG4GXxBEiPv0I/LpsVD8gBW
KrAb7lmYmr1p8pC3U/FcmrJggh+4vb2gyGXrs2SKPbLMByEtdLZ5yl6n9+n+E/UU5CEhqTwWFFLg
tBnHYwn3acrFlk0MBuPYFyFoFKGUuV3NuiTIXNxRzB6yXB7bjTptTLdFFylY4fllmQ8ezbQVf9FY
Pr+brQFcTBdD4uYf9AsDrOsgMkSPQgXNSYIprP5tjiZXU07Ok+Q/BbG4L+MYeIW/Cxp3SvObIX0s
RRv3Yj/KqKS3f93E4mE/H1ihbNxbBKSjZg3Fr2Z2fhGwnOFa44AuunzNhcCYu1QX37JQ2jBoGsGR
JXALN1fOGc6a5H58kbyBxYJNb44viy8QH+Hc6xJoUP28qioQ1saquTLsoThQS1zBefrB26n9W+kS
2OBNToaREqvUlrTW+bhOvgBDvoL2GSf9sVlcSZyLHGKktBuEpf3xCSn7kCoq4HWXviZKYUvrSu1Y
4ybTHa2+7ZEjumc1UvEqI7WSzNR9ovz2uGuaLVE4//A0r9kAcSXiJlZw2HAAFxh22Rs1eHTn3ZRp
QI8R1bHs8ArasewqFOQtH1wVj7j9/2mMywLVFQxmLJLpO1JqMRPs/ZOzc4n6pj/SDFxSjMfYqU2k
CVsGqfYsuo4dYAWSvhwBXOMVj/UGG6Y8Z1bK5+MuT3wZD9MBha9flSiB+9XJa7ZnUmCMo1eV1xXT
bgBLs9Yyk9Rfx+0cZVUgJYMgS7HAdC5bBnDLo7EacIR7Zr6l0S89flWXIr3wz9SvRhvHBsLDiv7b
Q4SEFB8kG2I0KTH6XoraUOABvUw43FvapWuBxHgJ1HP07TtHU58J6twRoamOdIOBq91FS7l7Hugt
Z+Gn95qx4ILIBesf7shQbs5DUUOXuVQIEDcpI2Fxh+Sl3Me1sWudRzMy2HFBUxah1UR+Rq6kBKDG
3fLWTmy6QwIIuOOLMrkcHMx4enzr3HBfKa6EeFRRe/+O+fYHBSGE+ta6BjFfbtUSIOAIXikWSNuA
G9eoIEdgoxKHeuNwLs7qCGVqFFVoeZvaChWIsQ1rDBjEvLT86RYoXIkVtitR6XXOQRbKbXBxkj57
TTWXkoADEk+h+Jb5oJGOQB6fvRwfAa49w1hjoJBwqKalqXn2Kip8cRerc5MuC8/kfE7vm2Q6wlb4
X2DPkWW1EMdwxfLD6siYuIaKQM6UHdqnUGxqtHJMMnd++IyXp/7wCxg+j6Fk/VTayUxJJyMt9qnt
LLBdwz9ry5xqyK4RtYYS9lrxX+XNVgVrimbV8jxk6KbhTOODssdXxnka63UCpTjMVksLChKK6yWw
1yY/kWIahfhMKgWy6BffPBvbt3Bq2PTFyH9/JKP8UO41RkSvk7Fpsq66wO/tP2UUKLc7FxitWQpb
NTNclTKlVUS74vM5VcIPJxeQFy8jnuyQvvAdoWc5NpgirJSUi06sssvklf+B70z4Z6vRI8GwHEoP
cILnFV8px4BsitifQ8bO7GiVbVmj/oBL7fsInSf5qcwkKibria5qaZL7dWArMxUKvZJVTv38w1l5
y7uBz9ZciL+CUIjeGkqMxrAlynIQ39e6dt+nVRiP4T0UC53PJOJ1Jm7lTHpZ/h7Z0Os1h9WYWxqz
m8eQWOETy/gmEYitsA+XVJj9pjsBLVGDz751iE/VWpxFxTZJDd9fONgtYu4BHPtISzUMikNEP7vM
lp/xPAuEpHrLbCp48DIHKhlQPM/gNmNH3/DgV899W4/Te6HjDbNaAzH57+g1waCg1PCcVf3uZF7B
4h6D3F9cii6asRqbhS3jjx3GUlHn890v6fBbiaG8nEj7wjIILEBC2ZBToY0Lc59p/uweyhW5YDDE
y0PHzfEcRXjLPdkRDS6vYxdMZoVFZ2x4gGx1K2GiizDjIUnTxVxAb1wwKNdKs8wChjH4ebAcX8fe
h7j+paKOlQfelR9yQ/kuQeChRF42bYuhilp+amEbVniKOdG0ldL6SW/cQbHsssKndFz+0VPaAbWA
yGaTKmwHQ89LsfEaiJr2VngNtYBvakJTtZnXzLyecShDXSaL7Jy/Ai9sGcmDBzLjuNxdiwdMwT1i
EtZMUv967okOOWWtlRVk9aJBTzBBgx+pHsvOTJ83DoU2di29ZYY+UyG+xfxiRvwS0zJMAh/Hw8bv
TOivT+pyhu+2Fa4wa4BtiOdSUAA4S22F1Mb000UDt3WbNnHvfK/66hOL/8xx0YqCps5eaE+RUlWg
hAx+5OrlHmFZO2rpSNVN1A8Tm5B8k7jrG7r4JFDQDqeTO+CDgp0PpBTFYTatpSu2RNK8NTNYkuzP
F1Mz01wcRnbqs7tGDl3WPCThFEOi6fkzn02NFnRMIebr2vobsQhVxYvQTYeqBO4ZOiPUDeQMdrR6
VV6mrxVK1+VCG3I5OgY7pdgjK3EFLC1qWLet6KKwxvpnNx1NxxWwAaVxQVV7UfDikHJv1GBEbsLV
V/N/oUMYd+GLs4vmRnAtoPuMuziSi6s1kzGJ9OJiZQQx9lX8Cp4uxPkGvuKZnEU2pU1H7+/MOstV
JRpQK/uts6Snosjv6e2WFFHseHnKdK3V2hWfLj+ilExZLGISvD1uu+dnLLnW0Yyp+6NaZXArLt4m
QmpJqlL7fVJkjBR4PuPm4rjA33b3Btxv4IO7p2yzUk1uI7hw0An7Bn1v4w0ICKuc4X4U9VI3DIRI
j0xYyQq3utrY2U7+2RNnW1yTLalteFFbe1B9NoWucjX2MpgHMuoSSf3/lnrEweT71jpGFC1eRRne
oHYdQnsjNCw32yHpEvaP9seR6IykIMzqgi5eg+4QHEmc+oQzbzfDVzR2nta72ofa6DxQ0hF7yKaF
1+XDUDWAUEju/NjoQ6Tr5XyXRItDV81YFesWZJ0QkMb4aW2U+s3/mN+GWKEioAF/rmIXDsiR7FoA
rJVmMRFEnPPYcmrfPlrdCCxmr2lvpOY3o6WaRUzhUu2UZg3KrvU/gQH7XYBLTbZkHJei5MOOPG8e
ErZU6ObMp2RzkXhBUDlnZMUPVoovA6BVH183Uh5DkB4aseO+oNthQQrK05ulNuWFf4MTN5Q0Bq/v
fEQAuC1zft7q4RWPjf8G9IfwWEYfqoVkj8ZGjE8jQpqsTUOodUlFpVuhhoJ9+GVMuNdg03rSOnpV
nOxlfOuiC8BsKKobXJR/yNjxSIZMk6Y7WHPP+6I1eKOKbgHbthZ2IkJF8u8e2esvIA/ISMbPT7Az
hgB+1wHGPZNXRX/5bq3sAsV9ugan529kzMMzP7OAPQ9ETZr0rcCMqwXPmnJqLUI509JdcNd0RvGN
AAceKuFXQcqNQF8PjIBPAHri2qfgCfCEnxETEowHEgDRjn3IKdz/giUnziIaTV/fc37x+akXVMyC
P4WCWkKUkbzWGYVMgIznqO/R/+youUOSnQu4mFNwx5y1dDAkquADTZUdq8LYSjH64F4/FYLhGQ8+
szT55++kMtlzuZ45L4KAyOwA97Y9QellNuFC78Onq4OjSg3ZbVNVG4hEPFz5M3+Ms2paLk5tYEKt
+8GwZD91LxpF5iJF6lzm9DazqjMrnzTxfmQGjkBlLsNurpE+ESJ/em26ik/mG9Ba8vD2seOR90bH
gddx3eHKit2az2GfzOJc/Wzrubt6ATdL0mI6WeRy0gdQRGu+uIfLNv6ZuUmfKsEH4DeN3WgkholI
9QRZw+P/lBmt8zcx3rHscyA4aWCF16N/ycymeO+w3S41OhmA9LMOMXHhktvo3G5qqm4Uv0P5uvsk
f9oCxqYYKMetz44jqYLYkMScQIzzDfUgs3qkULFlfXIRTDlpqJ/IgjUXDZBZJJgBOp1XE2PkOqWm
IFc+i1MAZYnQTG6moSvhiuA7KEL5bM9v3EMyMNs9SbN3KufKPEgo8gmLPal9qJB8FAuyEu3uMIjB
OBZPHBuT5KMXidwLyitrPs9D6OdbXfaZSoQfSkb6n/WmCosWd3JMNSqepeamaeQqVPx8gFxm772n
sN76tr8FbFtXY8nyh3OuATpAE49dMwDmdrKg5IB2xqqtaGgzf/Mz2JuxsSb1J+/mttDI6WnYBiDO
cOxUOdHp+zwsfsNcDPmteYhWCdK6YimdQePnms98KIwJutdGpIzWp2ycoeO+r84rC3IziTK3uaKI
LDC4Ove0qiOWzVd4LYQegJs9t4ggnyWnYplvaMKCsc7nxDMFT8YNI1kmnufrkmoSxeOtrR8vuyG1
fH/dHqVnJMdPxAjDj/0Bm11cMAs/HsPsyYZdXPhokfge4b8CtfjRPKo52iYtbaG5as0+WFtGX9IS
eLdttY4TUGvJZ9CsP82X8qg6B0Lchr2NO3Xx8Zq8aLd2k/whMwuOsJOoXfRoy1p0s01cvDRR4Rzo
hSJifrzRmqaAOhteG/d2EhloCyXpoScdHvjRtJKL/K31azCv4L7ahj9W8GCqtTxWd6tKJqGrRpB8
7Qg+DRm5TG6MGurI9zoigbgVtYqhhoLkAVlhTCFreUXfadEMITyR2zWawqy+K+l/J2rg2xEkMfT6
1kTV7qsKb19XVM7ojcvhd2PqyMDCrsy++k9khwRw4ykc21N2/8+EI/FlMARaNtVdRRCTnqfu3qpk
1f6VmNZvZW/nEPkDEhrugMFHhDeAHdr+FwEIFjYFQrR5mJoAblmkUYs91Nh8d7sAeJzesjQZsMj4
+RQFF4sq0ZHK8k5GGwzcrkeou+2vBnl0zqvGtXHKnNWMa4ziJKHwI+SDAhfZifal53f2LjSZFg+v
pKxEJgifq5dgOGYRg/KoPTxivRVGk16yxya6BvyXtIvjLCf2AFl9UKGvSqi2EG3JBK74hwilMgRy
ZCzGEJ5HjLq/GuerwvlI2TaSHRBnhslctq40hPPMBmbCHY+R4EuusjIcLIEFC6EG/n8A2Lv2tH4V
zuBEUabtSLmboW1sToDzkcuwVVyW66wBLcQMVvor0BT2Uqhda9mjvLqG87M4nUpfcKD+H7SWdoGK
gNgt3Yjcm5o2CRyJEKNnt5CAF/6B7aDtpfWS3GtGxPthl4xyerZDemr8ljz8riGBS55GCHuKCeYp
iuwR6kkgjAzUWmpInoOZ9OjPJxH/qktOhP61z+sOAAZXCc1CXS2r1GhEaAx5RhVXPAZpZlatwpq7
C7sYIsRsiC1bY8gtmzSJVZVDZ20tVMRv5AbW64jg5M6XWZW6JUXPnUaYtW5ARNzLOMiMLS3SjlGZ
s9H+M29eLfn6DrvB/25fuoPeR8jehSYNfFg7ZeeEmA/ns2mbJEdeYXivNLkWF0oUSeZ7UHcLCLFI
EhLl8YEqV1gNd8eIWQAAAJfcVxb4slu27PM+wJl2h3BbSnAPWAhW96EtdVUnZ1qWGJyuGbmzWL3e
sRCKkaLDCtqICmiuWm0PozwyS4r02mDiAC9iEkHUBw8yqPxwZp4r5lSBeqSDC0FLPglSx0NcJjtw
WxZNd94uzIAgJZqPZgMgDl/+dbYZ32BA1r74wB1jXgZBjLwPbHE6/2rCtwlPW3pbeK2/8/3+niYg
t7T7K9eNsFo+13i9NiRxgJKPIDC9lxuvM4cS+dqAjuLLN7IFnN8Mb7KxVhs/hmWFGrHZ24P8hSmr
hRI5FlYm/4Ckps7J0lSld93syvfDlNQ85iaMFTRlbuYxzJCDdlfs04ME0/Xy1vPZMO+F3AgyYHfM
BAOEZ5B1mQx4oGCFfpqEKFh4d90Es2rXZe3gt+AkVBO85ZrUG9NnCanvs5fURL50FVo6jPGTmMe6
lBLyWsHOVoj5uPu/WIvAahEKrIMVbef/n00fb6n0CwrfpkiABqqkaCJo0NiECpJRb0wcvHS8U7bW
J/wQDY1YInOUJ22tntEY0fiZrEHzmcAn+cmjZgrZtVvlcX2hrk/wUy8aSXNvOlSlxWlB+Y1CN+O+
nQ+j+plBxoWte77rLnUx1NNNh2l7hU7niVsmQ/F3KXrBULkOqyU2DlnX+BeRKwInB81E/7I2xLEL
TJwAId3NCKSDz4gB4uF8DMXbglO6oxehh237GvIROjvaggdP/ZClkq88JHCPNtWDKFzZ38RtRthY
0ZRBayPvxXK81R1jZfIc0CNT0ZeM8LeKbQ4PcrYUv1vwHfMnCEFtW4yn/A3WSXNovE1VVGl1MAd4
T4nopQxZV022NRsYbneqY3lIACOasyTkHiwfupSQzGPyXg1lDbLsZG/4Ohy6E4xfgrR54Q8FkTYf
pbQMEO79zol2MY3GQHBjul0DDn33CebkIEFHB2B0DtETTGxnUk/4ebLP7POqEO7ESatmSeKINL/T
awkQR/kcf7W3Vdl1gxBKyifdqoiwf+zlD/+u3boVc+zh7Fb9WdZFe2cOt1R81fQE4QDAGySY6xzq
tQvVqgSI/lQVrY1HUt8MPg9pYdyUS8GpZSDZ3uTNuFuBdlAkhBTJCEGMAt6VImnoZlssw281dkoq
gIpHsfipP1t+BhKP1L0R+Xn6xnPBjXomWhSdzvjzWK6AuGxcWmQr/4PQQdQuCMr35A+A0Qdkdq7A
2qAR/ZKmw9txy+aH1ofnYfdMx4I1m4CCRI8I7CE2UjUwORuyQr3kiiYbTgyShfzQ3O4+ViO0nGv3
s8Ng3RGcI4nbHyh8Upfrd6GfL+4zGU9JmBve1dd5c7pkS8LhlS/dZwZDhrlnQMhbaw/WTIh8a6uJ
M7EjkBsk6yeiixVlKacQE+MYfnk0N7UeX/gsPZS53bzrnSQOtHukrkyBBLrAhOvMIYDDc4DlgvM2
h93OId/mFr3p6BNttDZdhKuGy6b8KazfBei1up4Ta/GFPuOz00yghpeq6Smc2E44S5AMf0L3QJvS
XAIuIHX7swVaoPFj9OoOkZBxzB2TiDyzZx9CQyGDK98FhaVNizVnwXQJaypvropl67Zwg59xuA0Y
PAeoz270Vz0b9lxAX4NfhQfjVw4m1KM160eTB5/33GXl40PCXMB7MlzuYQn/oa4/pCt4D+FR61Oq
PChN4RLWHpXZ70qM5Lt6s9ht/MOQxT0LXtOPWIDxnyiH4fx1ATqFVSCd1Csle9RpCAc4+b7ulzyD
HeIqKIKmlCFjIjgZYD5PYPY5ChvksEOBaV974x16OnrvVv+umhBe02GrX/2R60oFSTuz7hVjovah
Uo5EQbm08+cbrFTc7vn8jkZJyBzdIq4cUXX90KyZAVGH70RlahxGPR8pBG5HLD2Vmk6CjlsDJRLy
bf5/kUg7MZD/0j1kSvEdtGEQVE06UuLUkX6UZ69lfiDPlVYDerzU7aJhZxxXJCVT+2TUVghbwXdH
ZZeRKWZhZbZSlyp2MeEQSXCUN/UIvD+eAzN0vfuqwe/rWiR+FkVDidfu+JKy+D97OdY1TdCtDEZy
4LV9//+i/n/JTt/rSCpF+tyvu2NW0ETQsTUo6huNl1iiu/tLkYpHWp44waVSbeF9vG974Jz42mxi
yC9HtiWvXu9bKlx9DgsI+qLO6S7ZHHRG/65eeV54btbmnAQoORgJeHbLIyqooOkgq8WyJHvsQGgk
VdzYwvwds04i+XwWhClaMl0sHm7nCuw5LXxxguz0o8d4w594etxjttJ4MptEInoGqdREYDvsWaRL
Bcp7lsvmwTHzikVwumvRe6Nluaoun4q37nQNdVCeGdwwjopo2SoMiI+Kl7iSjOwXjHkCIB/HXADH
sBdE1ILEWTnOxhnaw3lwdk3+OVPwcKbGd6pBYmEm0RvZleKHfLTxn7ahcr4Gm5EoCE4OpRPD8ZXM
xpPTWYLSHyIxLb+WMOIvGFKWOfAAB8dMIljiwi6ZsFeXiZSmj9EIs5kWjHi/AUXvKho8cekIaMAS
Y6d22DZchdsAmdw2QkUOBvplXJROqA/tLSCXKAJ1/0LbDn35f9c4F5TVbMrH/ZcM2UMF1Xg34hI6
3xHHhtFSCf0QAug4Df38KBmErUOIppgWiarh0a+2u2tSrBjVe/mVAEnMkOpZ/SWwE4sbPCWPyUAh
dLCSuYiH4V/+358eGiKcdXEU8T/SXWJ5xh+o4jKMGP3GgSYBCmmTMOANITbrqLNkoOmWvgV1ZqBh
Qusao8M/zCu7JdnPER4ub2/PbwWk5wTlWFMNjCtDF51j75Tz9MK10NVdWQWzquRZxOaXYIsL1RrD
AsW5YzDjVzWrR9ROQZFpxAxBHWyEp6stq0ws15OV4O6th4XOlJL6U39UfRN77dBcHNPW2OTS0EuJ
7kDb4YElmGFD48wsOsF30z6H26wlI0lOZQ175HqPFpjgTSjjvTILKv6dIP4XkCml4Zu98fFP5I/S
0E9gQXiqC91fhLcBSlR8/yf4BWS15yYeoLTPWjgHuTPTIunUjWL7jS6WyP01huYQct43wUsS0dgk
f2eL29+m4GpXCKgdtGbt4Ur2tXADFCd7GrZ5Og03TM43ginvF51CS5h9QUGYpDPebd0jOAlTA7Xw
OzhFbRjX3Md6I+Z4ISaVQqudTJw/AJsd7MwNQ/gF5X6CZfdkLBUQfmzvMJHjOPVbzw0wZJbka0Bg
p2MBfmACZwgH0NvgmjO0wEAFpZOdLRtxzGq13ta+QcTIXWYMOfFcKaxlXiFjLLzs2IgiZMHfONDh
PrpFvegVs09fGZ0nMbOzNv98Z9t58iTGPd5MtQgSJ/IysnOlHqtU1HMNBNKJjrzc8EO1SykxGDEs
gCZzMapMlaAnjmY+sm4xjG7wqa3QslDVgZB4HHVq7+SpaRlUQg6+RNveZlMvoY+ESROY1L1ZMfFX
lZSJ/ucMpIcssvGk2aFLSpvO3/9sYjk9uTN1aOHd37zDaIa2kdCusCg9ug2bl0gwhVkUOkoOSIy9
OJDzxua0bBrExwzF+Lc+swIt55KZS1DbRP5LUelHHGOVyaqzhEOnXksJoHLcPUMsh0cnQlNyad4H
Qe6DEQWj+qf4faM2fjYvwZckr5v1slPJu1cDRP/S3yYdtI1fwRxd5Hig95kEWkb56OHkjDHIeDWa
+xj3s9DKy0+rDOXEja4vQ2gOuq3c6qmXqrIyldgtCEnyhs5Zxe0Wyd7K5k3zf2EpdL5yxtJWhIXr
ugPgfNsQJynR+0yb3sZmb2CEgCrU1/F2vyNTWYSAaMTXozUETd/ieYuqn9I4AG5i6LA3Kf9kPpWO
5Sl6TeRqpZ9l771sv0r344ZlmxYsXa2HYTgEEmwi7/qLjbGD4mTzUDd9VXp+osfcnb6DszOap+ir
YJxGx8EdrkQ9N7/BQEqs8qccnFOVesKkjcAIyDo0l5XuSEd3er1YAtkFs2Qf3+8VgfjEZ0EHKWnn
RzWwuRMqNmob5TxQh5JsF0DXSDX5+A3HZiikIoJsyg2JPwQNAEkjOgNUSfZwXR4vSF8D38Tw2DUF
sELjaF94SVoVt/FiN1CK/mqWYKr8bjGv/Fzx8qiHBdf1SrEgchA9FKY6pongO5SrY4F1YR8pYGqN
RL4fCh5Pq+iklw9QtO3KHdwCP/hcSfS19chUshlH5kuFf/uD0Yz1QxGFZ3j+8W14bHvbpqEbqgLr
Apy81gNsvZJcQVOYd+YqEv+q90TqvIPL9n0pUYqF4gORw399m5gPGk4PNkAF+XHpXwRifbYJwl0V
Y3gdu1TZIeWdZVXah6hcVZ71/BxE50absf+h9Q1D44Y1NFb06unzapGgHhL7SY4IBSrjv0O3UJaP
oWh5+RqCVgQb30TZcbs+V8si+g8MfIVYXfMZ5BLyu8FpCfVDUh6fQdOzPpfrdVtMH3E31D6k4xoF
F063V4mc+5CAUwi3nbixyeC9mpvmsVL1Yh9ci9iyvHdY8ov+3F50Ot0mYIBcWiw6k79xkL+y7PLy
/N05O1/joU+GDQhdCGj+unqzMRNLF554YP8j4rmeOKrAAzp0zb2lnrOvOiVCRGoGlE77V6Eupn4/
z5SKZTQFSX3G8x6Yxrg56INHjKgbUa+4gMfRO64a1zcNAn7bpjl6Ay6X2lyafRTdHeB1Vs3wSVB4
fmlnRZ00o9u4ptNyPjngkFHJnK5b6OQULSIC2AHoRphwS1aRi6kRdXO2T9pQowVvMso+8O5DB0A7
v4kNWcZfrZ/PYtDXVDj8u1mgd8H/5t1jwo3YNjzotAja/DHJVUFPN7gkhnf2nhhinyXj8VFlkrSQ
pHXq0WpeU2r+2EmGiTOQpGEOYjISfPbuwfUDwsgFlAEDAYH+y4WggNTOrcURNa1XMKYFt2XYOSY4
iDylbYd1JeMwdW4ZkmUmBbomBYsmfUpiFZiqO/yb8sRAEHwW/UQJtmX9ii0GR2tUKBZc+hsue/E9
grRPP2FARd68sshNvFRVRQ9zX5lxVzHooMkuU7vDKnv2Nprqg7qg+tT5mFt047J+N1nP2UdL8mmV
sULDTUV5UTkKR76cd5hH9V1rYUOGCBuuXzcrk6EyRlzi1wZk24jHPfCXvOR9XKkeKIa+JF7VOPBA
ArxyrFg4KUMfomGPfQBqEbb6aZtyIRUTU5jRc0FuiCjZX8fqyl6ebSiqFbMfw71yabbWyDiApJhv
sln6aDiuRO/Kg6yKIltacptNrTHsx38MHpzl4wW0fKK7seqAjiUUpyZAFdm1xlfFZdftU102REDb
O9xDr67e0gAGwPeLRQ5QkkA/q/koZ5m4Lh0UYFxgW+p4HDgUpFaVPhBlegicvPx1kxoQwcU7NW+5
OmI+HK7+bSviU72J8/Q0oaPkWRHcBkFYEFoxIAhQLnsDIHTCW36mXdlh04Xq6m7cu++SkwdsX4r2
7Rp04fIWIY6X7LxrbQwK90Tgo4/nNzCovY5fBs3SDwqLrCRelR1+Z+czWaksxzykeZLNIKtEns/s
P9+onXzs8pXlN0csnzoMu7HZUbc5Z4sdZrbzIOlEcl+is8pi1mhOba5WA/bQCakKRFK4J8MeTNHf
+XW9HpKY1BU1aRoAxu1Uo4kT8qqr7p0MuVjrEU8hKcnynTdmwoC9ghleazIjwkAN+2QioJbDArVR
dfjCGxZo8onY3l+jXzDHU4t6eN+YKR+Pw3qFduULE6F0Dz/Ty5Hbj6CcMIFvCOFvRgq75oX/iUqO
f5f2WjA8x8sWu0UMQGu91hRHfSQ79Uso9PbVSLmxrHNReltB/hm/RZY12j5N5hCnmDQLG5uSgKfK
ZsSctS8CJcV0ns7RpYYIK4ONzJj2Ltgl6baeGHWgAFteqmqwMgWIofDB6N+2xynAJf1i9Ug2VjCa
7EYmH+I3szjbv03xrWCeUTkCJpEmKgTCOgxUZ7crJAaWUJqq3HCB/OUCFMgGutgvgU59T7DbxzAp
Qa+Z+NmDMQSOSaKicj2dAA/uDEAm1VUNtHLOMDlzDyujaq3MBRBHP3m5/lRwBA5bguPx1CtyL44o
XxDGmswIvxvqIMIsfBNZliPskqRTIfm2CSEf9AW+0oAIt+1wXWDT28bt3pItgACFSzK6aTXG3wWL
GOdw6CoejjCcUfZmbVo5O8pgG5PzBOVA2sDmnWmrNTZCwRyAU0iFKFHdt7Yw6ix1D+haPQPc/VHg
mp2hl/zrgImFUN4fde2sygiWodZtubZ9KMCTkJvZ8NAcfrPmrrVGdVZ6k4NYaLinA79Bh0xDTkfx
ibPu4RdiB7SI+VXpLTFR43Evir/ick7jbP4eBi/kzh2vy9GOGpgvBgQLeW7sTFi9TroNYfBdAANa
1Mdk4EviMkzDHssOo/D2Hc7X/7ubRfakaX3GsUTa+9Nb/Wt7G+W6bOJtjQKT1UTNy//U0iPxirVA
EDYMJJgqAVRU2JCJgkUI6aUCI48xVCfBvxSOJ+k2RzRTueA2jkoKoHUnLCDjwtBwXHx/SXSEzvzV
f8gYCCJA6qt/rX5NsN+6aTuCqee2SGKgMcfxgFNGvAkr07hDRDVwjkSNFobuKRdT1Q4MmzzvD646
jos09TJ/FbPLWMKdT7+NUksfxeqUZqS8PJg1Y45mIB57t92moLuEzCismuAIRfhSvpptl5S8H/wO
DTiNo8eRdCads6pVt8cxl/L2L8s2VuSz0za9zFIwABc4MScUFt5bjd5uzk5PNi8D4Elw/OWvfgEG
oJDgYWmlfV+Nyb7RWe6CohnElSpCRBFaVBdoq5NuU3wEUMY2LsUZhjWvqgZMEyHvEU2g9/EtRPKb
zQr1AGNQvH+4JALj885MUkbgmh1bnHi0nA3zRwlZHccw+005/zes2WGMoR7HDPvtmq2iLXpX/Qfn
7Zc8xEZujmX5DiIKgI7dV2k4AlQdmr2ZJozAQP/EXBOye8eOko8qFYkVmNPs+AZJqjgn5hJyjm02
LNngGHkRhS3p3yK8SuhW0Le2npyu+D5JDo2u+BVjB5ROXTWpRqjbSoUh37Auc74gB3MGCtc9dswt
PP9cKkuYGLmBnc1YydBXMUad9T6wnBvi++TZJEmnsrZVafuQMG74874cAg3AVJJjaaJq8li0XMOa
L8r5ipxAOnpf58XbMeQmbwjeP5zSfcg5f859I52d2Sy93Q2G8uLt2mvfDkI6/6eEl6mvhYQs4PeK
DEbuxKLXVJ9cfRlXNIWwORVb2pURVN9WNw9/0L3p10tEZG/jg5s2/yFKG9aUqWjaP8VDUfwNqJLS
cjeF9Vynj2N1wlSdFO0WT/yBGT7tBbMsRBA8EcmwyFNuzobFRChgdXU516AehSam0cT2f3YM8ufs
cWl7ZLrHLAeHDHj6dtBjUxEl5BeKpcxXrDSAt3irgSAulFLjuY+1tKmih/JkuJfzeLMazAivP7Mw
r0BRF4P0KES97gMCZhXIUI0V/ImzIzWGA+vCIqOdOzPRWu3/++OV3KYpJJ0QDvx8ebnSzOwkytRJ
bP1/Ued51JNYVi2EN9g7t0uiaBLuewwO+dk8hhK6v4JYrRehN+zJ1kfui+yXLCfi1pKeVrlUfekw
HIXVnCnD4llrZ62mKzffzRbJsu1eNvotg+r1b03BZIzyJwusi5siYWJkvFj9JvvlV4s0Ih30i8yP
Ml/5qTCcOsaAz71PfbDria4Dm7+3xSrnMWNL0ZZU/MQsTdjbHEaS3QfXZ9QQqBYbcLywDXWvqqzs
shaixAbNTE7fsSzajbd86WEGHS7vaP+RW7F2HlV1T5q0INA5TN6u/nIg0Kbes9CBQ4QScu2FN6w0
8CxuxMhIDz/I4yTK65TJ3ofzTexH3zE5oijXvJN1c/pI6mAEQR/5XAc5vSDVwLIv6ANI0sh4g92g
TkvVlfis9ank74aroFFdg1OuwAqDqcrN39sKs1y+7KofGHGoFs4YA6YleHJZi30NGLrRS2Lt7W4K
9HMjO783kVNFwVh8VLG74Fv9tNOmRDUKOS3ni/OD7JfqdW8rFTMH9o4gm+WgyhaZJoQPyPjKao3v
8RYcmSPjmT4gGKMnXT4wOcIYPG8OdTeEifmOFGkdTvHKVaJFyDjtmlc4Aaz7tNjlFE42J32A4Mey
4UhkHaSYtevZP8wQE5e5b23W0O3J8tt8hoqQ/31hwxsutcYtrsQQxJbjkozhnfhnqHdEJql6T8m0
hFh+6cV1Xz6eonp9FCNxv5PZ6795h6lNZPu1jXZZPFC8X52TtGv2B37gSpkVL7sjwsehggJVQ8Ms
SrgJeSQwEgaQwW0UGpStID14BGIgg2sJXO4hP0SjdG9s/8d1KsGmbyQNSXrfV1m8qsXJX3WYUm7i
86oNG+/Z5v1y6nU4NzFmq31AExklPP0x7IzLMuDv2ysL2PdNfBsFL4iY5/HlF7nL4cSYEaaihXIq
+2thc844Knsvctw8dbvK8syQNa/OXaLMWo5esW0v2bruEq7731c4q9Y27nh9XccXthgrDJ/ZH+8X
ZFWgrz2Tp4IA0AG87FEIrZIVoxlMYgEvoqEJs8EKPGE/RIXocVudfV6ewOwrpEuWaQw8nkNHzQyg
XB36Y590gueMevTAP93F8BkaiKpmE3cluzULWV6SNxrIjpO9AspwYH2GoEssmXK9uAs7ZpjS0qXb
QLre/2MWrgTGjjHnnToZnklsAlmBG0gB8+wuAIjKsXyLoP6VZ+s0p8PwubqHCTy2w5kAmuoXXsWb
09Gj2zlRm+Szl12PqNy+DKJKT9nyv+3Q7FpKdj2ukrWAcxCa2NXzNsUfv16cDr9moatmCIyaCLHI
bVgyCMM9BCtU1qVApit1lYKUDn1OIszf1rySiG0OVM/E2vWNsFmcykLbynSpVmJ4afZYTei8BziR
/QB2SMeBPmTcLFsLc/zjUHTLBG9HPC0j8sZsBkLRjxxVrJynQsPoTpO3grGSjc0T8CqKW6TW9xZJ
oD/3rTycJXitrkDLCHkrq4bYMqHHnI94O76QmfrecwRc5AwCYV0Dw+Z1KrJQPofT6s3krVbp1nx3
TYHkrTKPOIg1lgZpV4n8YwiuV8BJIaaWfvQRo7xvxpv/3T0Q+EaMcO3p7rrjNgZhZvtLfQrU1W/A
sE4IANvi2wK7Pvgga9+eNY/V5IMzhgQ9BxH/krWEm6wsnF/CDpCveVjwQ4qg+c9By8Q7UUbRj509
Sl/NjecIQjwyWcT7WCElD+tDjkCADLd/UT984sFqpT9Ieo8g7jWJt08rKqyGyo7iITnsbJBCT15/
rfTdFAdhXyTWzxVYdtwnc6Is66nbmeT3syTSV2hI+s9b+MeoqDgoc/IFfsIh7ixrJJ9IeBLa7zwX
shoerTTFHbqeqWr93S9dhcTzxpcSbTlJJbTnB6FAe/kgH1akpAp+h+jSCGydwmlFlz9kFq9rDHYz
foflf47e8BqUCZeXBzUm7TlvWybD1jGsvYLAAF5v7LvcH06X1XITaaNf6d6G+06p0pUtYyOqzo+F
PkGhU4rfxPgRyow9Q63pAuCoS48jp5s7IWA5JkdXZfb4tOLXJk4MYpfMxpoOFCRDQ0AQkSqGdU/r
mwSN99kRBxk18igw7r4b90M+eV+uS6HF3DSMZHxD66ChIS747bD9a3O6kGM9MREjsFhJ+6FvbFri
UaRCasGs7Wn1ZbbFliZNng25cbevCGQzbx1PlEjw3X41yUT0ufVdyqphzadtLQREi31sklj55npN
Py/2LBRL6NoDkgGv7cXBUwaKcLNkfvatH/2XSrnBBFaenr3IPvFeZLELC9sM6SlwqQyIoJlhE0FV
HyEtVyPtqwWatVCWZXQ5KYA8/e+sJW99fl5W6RvZ0laS/68DPM43CQyCU9wqNUTLC9uUKVcHb6XF
BUMyDtpa495Npv2OMMIeN5xYuwHDywTBTrzcGnYtrHdEzCkvvzNpC6nB6qFgCKasn4ELLLJrNv5n
Hp9anB8RWEYV33iccZX70rRCj7uLyEcj1LzOnZtEIYhyhofj9dZPftD7+6AC0ydi8gkKayA3C53a
d71taeH4lymhpoKeUiivIaJQRUjtvCpJHmCyzibOU4Lju3b7VorZRv33jKvCjrdchAKO5qDiOYgC
RhaxIKxZcKX/2ip1dILkeHnpCsFFB/5tmntiFclWv4lq7wLm/3o17F9PsCfLI2c/UPDgmcYizhMM
wN94szlDb6chHOM/nXtoJj0GlxtydCzG2MmjKxVR700YlI6zbqBOiqCK3CU5gxLjgDNCflixIkyh
sMmGf95mFlJ+d28mAn8wR6NRJiEaNbik/BK2ICo4RXBmUwFTp+rtnJ05hEWJP79H9irtaqoMY2kX
EGPOM+bDtwjzkwR2tVsriWGWACvmHnw2QxvcJnP2fRRPqTVmaUrLe7/cs1bDsKBTWK8XXyVuCxF0
GZRRu83gEU6GbGmMLvC23ireWVcC+hmOuiFZ8qpv0ZKzCf4KwnnK/yB2gG075XTLIb5lFJ2W+m3l
Jk1geYh2G/mS7e2Mar8qyC1nqhnCFKF0Sl/XKFY82G8TRGzpwE1vs/IS4UKOaeCOvA8N54ApE6xp
x+74wV/QB3YQBGI7hx3VOMUFyaxQN1ZHbIzY1wQoYEv5Naur169gsyJt6iqqhJ1tXzDPYnpGKeiZ
o2aQq73s72d+3i64mYvww16ySaBZe90LhIC+FysW/CqojBbHDAN8eE89szZ4qNuFOedxaV+39w+C
Lw3iMFDCw57J4uE+d8BdhZ1Rx/MXDOnsdlu14V4xCOUrpXbkhNC57jWIwZ9nSHUiyev7JubQvCIE
SE1q8MMl9KHmd2rbtUPl2MNHx5OlylI2Dbdo3ULRZ9YyqiR2XWH2xBF3jzWjWmrj5djh9JwBLGjA
GIau4wvL0k4xADIqU+e3NYyVBZ/wqemqCbizmKqSufbQRam49RsAMe7BK0rIv3s6vykHmO8OT+qS
MSpbnG5mcbEeJrkDEWx+SDJ2pFZRLKST/23dPRtvAZZVau9H7N4/fleIE+9ZGSnS1lXxQk4FbARo
s4Wd8k81khK8V2CxoY7wMCz4U6PPsOFiEfcLGAlf+MLQnGAVw2ShkU1i0xZFheJcel4enlc7dIvY
ugPgIn9rsFMGPH/q0OtqC+vNHHq8xbqYNXO3fnbyjxXnAnvoueoIco2t/FUrQk3hAeOTd8IVEzGC
qjn2QUeUfdRcgfuJ2pVE7/L5fyZhnqd90IloGekJ01eDe29eFFv4cn5OWQ5OYD/Br51X+JfubWOZ
Mb/i87kXfEcB644jJ69EQPhipR0IMlaaJH9l342NEKVdysAOGr1IH0nYB/DlLZzgigfxEa4EiCwX
roW6vLIQSgjsqv8RUVG7MrHm+v2ArQ/AHJOGZFSdiGR6eqZ7Sm60NtK5R/NXnmnAhoHTsFWSuHxX
NYV8uiByunkdec+JqVhvvSNqK1s14UnYrqYF+Y9SxaWqzBOFipm+nwUow/AqZe2zD6tdUf4clZEb
ivXOXZYWSUE7KjMnxA9UTr56MnXcNlmaPxvdmMp9nWjZ3CdyZERv0+K1EoRQ9aJ0b2DPC89rNegm
lYwUQJB51Adnog2z1QkxtO3Z4MJFTETsFt149tQ9seYQGT9B0swe/Y6P4QnQ1ySgLd5LqJnm1Wrx
/sxUr8/bdJx2mRnLV4qBiqdhQow569SBCLklmSuxL6+FVF5fSKxt/QU97oY/D6xfS5y3xTdD0zc1
KoBKWHiU6p8qRfURhMqEKa9794j00HmppehnKvzVgsijdtDCMJ804ALwIh6iWh1lFCQ4mqSVmrod
Y5cAuV3jt/6t46DnrMFpaTH2eXqRS6+meY/SCv6UQGhvVcGanc8G04aUi4tMXrla8IKjAb1+xfJI
3ekyhJWz6X4aOBdSEuxF/infxdPFSiR3NDhJFhnxNbAfegqbT5kfn9S9LyqnJnzXlIR1JKtRAyr4
YC/Pi23lcNx+3aEeRiphTFH/UVVVzXlyNnZg4maWAu6TU0tzQIDc+cUHxoBGE/o/JZG/n+rNQ5xM
Bj0Inuk5fxP237flISriMubv1gdPJ4kg3rZpWAsUdY+hAaYZs7HGRXqKwNKSYv49ELcs/TmIsBIt
6DTFPTZng3kb0HZX06YW+ET7vNMyspeKkxpozMsCvLJPEM9h0fLaRFXK6RatG+xctaBQoap692Fp
B6k8hYlODAcG6J9ppfBQ45MLi7eijfWWtTLG30M3hlBXVEnrT180A6GWLhB5+UBbSrTd6RaDOSAm
uaaROoLnd9HdxHiMJih0eGyyYIiHUH7OB4/buM7cPe7KhYkSXAL5WE6dQtg7Xsp8B5MkjMmqCOXd
Wd+pPH/qMYiSOa8Xf157BgRf4mJPFp5qSOeWpdr8fGyeSMUZqcBktOwsAQ0EqcRYlau/x+a4/Rfx
c6BJe2dwjicneAypwPRG9mMTY8WVSaBlZIHA+tFy4BCQ/JV6ANHnp2qLq03m7ArH9VFjrQdEAXgJ
ZM0JbxbZyYUDyJLOh8O4zbGhp7DIVeAM2fYZgHyfGzFBYn3tCH9KNQmUB6fZTAmN1EYFdHURFEtM
fpSp2tc0cNwEEmzWDSScLDYw43AtoBM5KfeZw0O4apbJuluTTpxSkRfOMQOrvhnELWSBSPa7ENm8
r/wnr7B8PwVahmIjAAhG2bD7fj8JVPke2oj6TW0hxv57aCs8+qGeG8Zs/u/fj4aZkz7vEOmpMdH1
WYpinUQsTLpzBQvIdmBa/f9w/Q8rqpdkA+lG7OWjCt1CKOCviCB8sZnhPFN/V6Mi/vfyyUwnIRAX
HVjCNFB3JSMjzCMuyh2wJxHimhZmzkke79LxVU8gRoJAK2wf5qlKZzlzUNzsNgjPnygcxXx/yhbL
zpMyeNHa7Zd1yuP8/uRhhWBFW+57knytLSTZhG3Z4K/fTclPIPuTNmpJs9FfMW/iWXPWvc0vYpmd
NkRJ9MPY/NlDKv48EKsyD8oWlSQ9x4WYyDkgfR12lVgwze/oUwZjLojVlZfYhuSeeG2UebZZ8ESx
LxXdQHv/ViPjO4E475ib6ONayt9nyd8cm5DNsaZ/4QxRmpFfOOcgbxWF3uh1hdoj2073kudi8qik
HdhqGog5pqnSZ0er9HC4JNiXk8HaNC+RukLELLSrg8KcSoX2D/7ksdeXGPNI9OkG2cecsuzdmpCA
YE+F9UpCWN3uIV+xNXrzE91+gh62P9bDVX3BDFkr/498Y1/c0KcGAyVxLiXk2+J8PGa7E8UYCX3Q
rYjns+82qVUbh6QQn1yhZePOgSN3GDyHPlcY/qCncJ1Qk1hV+buUl1982DPk+0O0G8/C1f4NnJrt
Hpk4YIxff22NgfJ1FdPler7ANPesG75K1vaGa5hhhpV7JiYjrUTZ8idVvyCTn0jrHgAbY5BFAON9
YRL2VvEnxPOr3aKnncttbg23oVjBS9EJrZVIh7HaNjTsPBkGzWBY5IGltkPUVk7geLXzbplBflDT
1g7zR3rD712Aw5yWKQyK9/pS6/4OzN6aVgwNHYqjzyJdDvNJbXsRmI/OtIpEeflsanGgkZ9voPyf
Ns54PfYW0SZIdCJUJliQOhHOUVV47Df0t0Ytd09mf+J9lua+c92ACrrxbFLOcLzhv+Yre8ENH7P2
2NQJWfItb+rI9Fjix8fO0UUTufqXRRq4z+c/bfTIKYu6LarvYR3Z2FsZBYjLjmOD6m6+Ohig8PD5
KQveYgWmU/cQfVkgOfce85mT3ZUlBGrZllk/MyM0XXpOq20g00hG/KqKf4QNZa4Y9PhiZ/J3JxwY
QcjiJs25cW1daoHVYphvAvByK3uWgMlhBJRE7FkZ+CoVTtrvm3Wc1DcGBea9hP63ic4iSm8ZHiX1
1NeZjbUWdcN8DUjf+CaKHaXeKwdJaBpSTKWq+ExXiePpH1II1exBCiI70ifN7ZXFGHmalxN64efd
3YzbrobpJSSOtrTAbv0P/mT0MgbSKapqIb1GxtNJ3RQJBrxVLJnhvywmu9XmsP6wTewH1j8KyZSp
u/eyUEcoPyO2JLCg/9Xyfo6atvGx4QihV/9CtibpHuM7NYjEyEgNTi5lmPfaywHXouQLcSEkIi1+
HgpIbPUPT+6EsKALE0IQZrD7+eUMBwi5BqGSWdWu0xLyiFWM/aSawuJiWMIxfBqy83/tE/jVKpvX
EpQqgPo7snLaJmTTvvunOyiYBU7GTPehgfwEmgbxjMfxMlSWmxKvcsF0Zl7W1x/of6w6nTWjhMzp
Ak924tHJhSzkHTMq/cTnwUI2/ryOK+s9vf9TUTrtdnHMyw1YXhJ4pupZmHjbZb32ktyzSZPem78l
Ffqy8nzPLXUyWk9zzXOO0CHodbN+rwCwuT4HBgC56nyo211I0GyRIWqIC2Gq2C1Pur9k7qvb5XYp
UPeRo1Ql1SQY1Rp3MqR+qx1lgzTnH/9lpNqHhob06z3oM3tucBGR4l0JvRZc0f0TSbDmDSSmSKHy
fy3KKoGosSrOmzvrU9Lgv378VCjksSDvItEIDf8ZtEVS04fIXTL+47kS5iwB3LNAxTmSaa1OMjjW
Vgr9LCSwjlhCgNXtjZ9h7iAO0jC4FjSpfLDlfssSbsomDrNR1zZdjhXsRLejivrdmXoBIprvpzlG
FuxbFpBRev1s+J6FvHPbYJuxRD93U9VOBT9tt+YYcEp2vDljwCmksCD3EdChsPb6QiKoiJSp7xbn
rG1rxb2xoY3/ZAUmJX31mr4bUB58s2iL/KkbAAPCgXSGxSY0osPsmT0c0X1suQPuolrGN1P6wPiJ
jKYnNamGJ2FUVCWajKdBKYNn5pzhddnGwe8UD29Gdfp1Fb0CXz0bdyFU/gnOeDQGtMFLTr0YIkZd
mi/sPg3FZpLIjJ0eIsi453otMif/Wdch7ea7bPGrnAXeLHyX+BEoUGnmknUxxOe/znjgvC7qT62d
7joi0srjByRmY/6t4Q4Qw/wI2QwQVrWt1B91ZEg32q8Bb07LjW7yUUv/eu93AB/r5WRnA1+wsq4p
Fj68XXZUmi042gLfMOVqvGMzB8H0oxR6+sn7xqe+3ffD3TXd4WE3FsEnrBuO6u69EMU0mha1QTD9
V9wOnGHNpWITMtU5KfoMAtn1hWGHtVN7T9pBldg+MHhk4Nj+zeHzspjO3IMWfdF+SZFL0KxLoORz
fDdIJ9WrPIIspRUBIu8XdwnRVUNmLDYwyy2H13a+1+J4+NInGLvMMX+vDZuWureWQ2W/2Iebwqzo
r0bp6i8fsUGV1xrgR31pDIeWqgukqHZf2URlfkcnCr8JHB3i2RRHBNNzL7oeXPdoEkzlB4NI4GkW
WkF81plqUgvaC6WrLeah0EUdjlU8ymJGnLSuYbj6ka7gpuK+zr7W3n+Cnvo56gGgfV2sXe0dVHiB
ciW7iFZ82H09O/rss3iouCZc9+FVng0+s9WtmyO7aOA6A+qm21mpvwaPMhA4UO7yVHe8kANPkG2u
swa/T9/I5bOrTnDYJPt3CpNm7cmyUTcgnflO3DeRDQL2dPx9Zoub18BuernnBZwJ8pkzfZzwkMOs
O/XAiJMSHwuFY5Ci6y33IFGigi/1dEJQsdivG1Y1sbWaGj4NiyiZQdnSvaDSZdwBimnCACSqCwK7
V7tQVu2P8p5t0T2CQMuM7w0mqLZq1URGUqyU6YFn/jrEzhgMk1gST8cBiaSZGNb4ZAtQx8u8/T8X
UiRoJc5qX/RKMrOTn+0ZA94OOU6J4pFU1UriTjfoqroCpbpeKOA6QEXBhpyF0D8ykfH9B0w1oA6e
NL2Qsth4N6Taj8gdbwFi4QNG82ty6MR9aEq/PhGAShmFiyZ17T8iWnPanrnPpO++ZYH2KwL45zS1
3jvH2zEku6dOXAVIh84lTJLZ0WehbB2g1YkiZggL4n8W8hTYRr5G/2zcsXsdHB1XeC/IWCy3yToq
/l+CysuowjvEOmBpCzjzj8ZgwdBPE2sazjdSrO9DYGwr6vGaI76d/DU30gHy4qgIIjs9g+fltC/7
QTOinmHt4gdMzgBhwElruIUBghfeHyfJLyh8YPzyQmyDIgjj/CZZR6THM6hPdgNTyf+8jloSDGPM
F9SUDMGka0z+W9e70KLYFiQ/i/TawIURChKFnt+uA+/1sIdXTBtiZuCpOIaOfFCK3rw7gMg6BqhJ
4wlv1dVSan17BnALJYdAya2P00GaJxmKossY3nmWj7pBs8nWOrh3uAuwu4SWfDByd3KJU9wrblax
607tPKzy7U0IH3vQnj3aUDNKEPTqcC0j/rGICM83UFFXtuxYKPSgsjkTL9c1/qCtjtJ/U7N8MnB1
fqO0kW2tXe7aSni1t8q/10NrHT2l8jkUtTfIyOxQ558/lvkmhz6doPsVGGUpz8/97ZuCq5IkrpSO
utDWdQenKCJ/DiVfT+k6K+RkWwaCJLS9iziUOc9D3BA8SY/JkLdTWSuOLq+FA4/lIatId5tzPcg7
6nfmhZnJA+9q8Lmz/V9KcA3QHmJ0PM8IxGurp9DkScF8BqijO9+md0FLWFFAtzaTpl/swh4d2dVG
QI3hnKdxaqneL6grhqXXoewmlmmx5RHOJRHzdVBE53Qq3O+uz3ITkIl6K9Z7QpfcugDBCefd5WP8
+xh41M3RELy1W/miqcCQTfCg8izZAzmuX9jt5kH2tTXuQea8/yI7aopUcuIwG6FP+JV2tC4Qr0as
kPYh+otokmYV7E+jMnUOOnewrvjrfv3K4Ljy3p11TS2Pd6El/JmCRS04aVksvHlpPkyMgTIEHJV6
dxmnFsFX/K+ANjBwLbfrFcatYbUPYTSIwMpjFsvk9wYyXtCzglO9LCGydh/k2pNK9RjAuG9IqcTQ
ez0IqVAKVMYaHqz5duRkUvt/jkvGzhkcyzELWCHNE4U3DIFopcshMQDud213Wnd/uTMRoaZfb2/R
pumM+rXxBfNvl7qyTOIUrnV+5edPsMElELoPZbFCp/BB8j6sQj4cwIWyOT3loluzvVnMKhtmf3lz
vKg9dB0bREUa6NXBG7b1N4dFO0QsoDByXg08Yjh+7ZIJ5GxA+xpRY5TPZhpgkUEUE/ark8VDqiRR
J+8wcI98DYIjMGpoB2nB74HpgktTKtMvKG6mzsfLdkkU2mb1R9s38YqVHIc9x4zp8ImO82KXvqjx
LfWjBfAkw7TCeHFI2qbpnEFXOWY9VeCmpOTMoyC7Cy+BZabei+Rm3+Eq2kVh062JpXUgxfVIdJwk
wiPMQyabgi91B9zvwbWlZt4nv9Y1MsA6YLedAYREiUSlt5dyE+cvgbKVOaV7oX/AF18P8jqFhA2l
OUUKPnrR/yT3YI1KP1PWxb63hUFAtPQLnKFeYytETfHHt90o/4llZBGBWWMGGscmYW9GADfkXkoM
OJzpITj+MLw428OhhvzsBLPI8ykBd+w7od0hgMaZTkCdvK5i0JPm0GFMZvWrp6UQRGLBe0+3w3EF
1hDQDJPcAB04wfj2pgOtKFuokSitFgWVdOaUwwPv+xytxmMgrvl6vFT7Kcw4mvz9kEhOOyGpTz9z
JZixKmh2RjC646HBLAmugS1kNlmwQGtq+ThwRbhpeEFcmGI0pBMAt5O8AQnm4Wsg7FXrfyDC1luh
0CDvSlDy7bK2W4ZSY2mfmhfB2CGCUl3XRLbDEMWHgHiDb4ymnAryLtgtoLcXkodX2M+3+9VRpKT1
ipl/m/H1XXhgZQVRUCDhz4mkEAA+ycEuEeJbQJ9FTfb849sS5y5LnFbhWazONKyY1VlnKxdxHtZ9
fNClehJ8cEb0efQ+L+NlOXELjb6sR8wS+BiWOCwPNcTjNhiCxDAzmqOgWGxy4fzIpIWFgZNsJXBO
p4oZnQ5G2ES323pTX9VpZnXlAZb+tYVSw7cS2UvBSN6K+1fJwn/9LWSdaYvDIBWlosqaHWa8P8El
6Bg0tDBSupLGi3h/Lire3//WXpg7DhkFrYRzNarWG7eN5Q9Imw3PK0wCa9dIDkd4D/+TSzllZbh0
cCV+v7jfymuwkGn9SMxaLv/MGZ5KvKj8FTFUCqr7jSwjy68MlLyzpmIy8r2PWLCZd1z17MTTWZjE
oVEoOmq35PcsU2BtntMlYtUuqh391Ea/u/6B0ic2DXaJHJAxES86CvmkO1yDijGpVimaUcZttjte
NnQ8n59Dr1fKM8QWqABmt8LxefEmVyE1FGYDO/KMk6pGCXkRzkmMvefRlvuCSj68wweV4xO5zzFx
YDSJd2eulz1TG9QS22HaDYoYK3lIpZGN7rrKx3BRhjprwO6s9RvEA/IohmB6884fETkX4SvDU1pW
vPFGR9cusNSNNajcEKo2xrKENRElf0o9Mb1o4UsXQlPCZ7ZwPPATtiQvkxAt3UmPe5zsD7RhZriH
FmdDo/JK5apxeEa569PC+NB5nXCixBz5oHlpdLI1BwkiZezjCaTMrJahHhmg6vYr7nLLi7LNmDSK
G2EA94ZaJ9FhiDrJotaWznBtGVgQj/r4XSlzuLTbdPOsQthuElbdyuM+lSIydtxSnvB7mPHgYieU
fw++BY+Z26Kicvqv58YAwoJ5Obrb0NCBMKWKNP/IwCp3MsEo5cRDiPFY9a1r533aXHzbVdJS7ipr
9R9yvI056RCNLbjTqqJXv78MRYxjvhRQ/lWGkIeSdVtX/7rZI3c0FKE73iMyRZsFed4UcCZ4ieDu
UmSb16PMvx4gFKk52mvohVVwWiHazjqpFLkxji6VyjjK7iVHsJIPAulmW+bPNusXFPXebEtPKHYA
m88vum39PYL5gln6j/g07UFVWCUPZmEwNI1OcbyJlh5yEFOa+pu8TKR+E4a32o0x0hYNntNaBm/A
fkpq/HeFtJRHMb3m6FanLtrC6ZrYpodwbPDat5LHYkUDeHzkRLIYYM3HSOccHQ8cpc3K+47cacco
ZFyfLsrDxHnEjepNg6V3rraTEeWx9c1i5YclLLCzPkccV5KwGEYhp3LZZ1KzQ8icYGQNQndUcth6
vV3BiBhuvf+IqS2DzuBVL1LJxBgeXndfylj7i95W9UNCFwOrCNJxI9eYt021VeZqvOgqyPLNmMEQ
mHE5ff8Sfhl7BeMUZU2crZtxnXn709sVlmJErHIS4L+n5ZpDipCHwDeOhElFGecHloTAyuL/TvCJ
UKwFWnAEMkGKN2xp67pxysPWI78EOg9oZzDTCMLnYRInfQZzuMGrH5oNnWcmo9QMUIE+bAIO5Zo/
/JPv32tOdjFV8X9TCwAv7kaWGgWtdnM2ISAtfBGxX+PMDVXcSfXKQyHx/INGoPnHCF8qU8wfiA2/
7E5CKPL4pJuZ+/BfzeftCBENlX2sgqeSpNSd+Eye4AzFzczbrAVSYN/CPE2pjqRdoniW24DBvYzS
fF0nFk0ivi6tjIMMa6uR4hyjhDnc7iYKHpxOpT2QMnwqhaac81SO2DtpAHxF2uSCIaAkRk/qmJ8U
1kxIZNkKQxxfQiPZxCujXkFTYyUF4GNc8uRiN9ysINDfAU3f71ZQ/8T5HprGEvIjyfqjjGa8idtA
6pTahuEZW2C3LLsrRZZA3L5hipGO5CB05OpZJKS08F5CgbPXcpnK2xk92hXS/5hG9T6Cn1NkFdEt
zsgRKD4ezurBcWEqGwIEDlONgHmmnuoDXSieWQss/3OOz4KqA5KJD8TzD7sG/Pw/4kK4a+ChihTn
s8jRlcOjQiwgkysKbOJsdCwwLDLZGntiNgWQZ2A4Ss8Laz8r1h4+Z5cpweFgv3X6mCLoAh5ptyoD
/OJ3ldMiTYLTTbKgpghmnOmqmDpEb5YofmkRmqCP4UqMAA3uDeIwpHxbHYa+NjuvTzaFkoaKvH/l
8GPMRcFXpqaxfL/RYNZx6jibCSoAjWuukvBxaYL/P5y82QuEk0cos3Mmq1lYX1GIM9GGUM7KCWUr
lehnhMiJUUpOhUddsC1WxtVrFSo1jIV2Ecvcaez+MVVT9LE5KqWCGaBA9DBETLHxc9rW02WAvR52
hO9l9D8+NXSUxtDQ38THQcj/VOtQg68cGYYjAOm+O1Xn+utAjVRJqznRheSfclrAb+au8iOcBkoL
w8f2Pn+u+fcTOvXEod7/WfZoNwZaO7xUpzBvgY0zFbj+O3wjQUFww/yiHg7nwhU7Ow8JeNsoK9dQ
3DV53eNu97e4rpszWDz7DyS7apqE3u12gtQ69CDIEZ/KtyrHHuGMaEBOKJvkjzdYKJwgWrF+eOuT
ZWiwmlpcRfqzfPO3Tp63s074ylF3Vzo1o7N6ivimS4AmUjc8Jp5SnWPw1/qd38+0HCjiOWJUUnX0
4yzrM7uITwC3vd9Rce0ZaIEhrcgi0wXSCLUEfV09psYbIT01B60waVbh5SZmaw+gFhkKJS1/wFrJ
43MNgQJ8UAVtb+DOvuSd/tscexUWxURcF7CJIc3pKn67dApR+wfOC1ItTDFhWim0PbVjzKG3wasi
ECJ37LJnB0UJRAyPrKAFCToZ/6V0nL/h42icD+vHhihX5HeCNfD6g8SL8a/rQBsnIMLhCbkZa0+l
fgn3EnM3YwGWejp+H5nheStYpyk+u02JV5QQPqXyTqXcEmKOhV0+71McxAxbO2CVH3jVFeH1YHm9
VwxJYq7E2oRKiIqSAxYmgzpL1p+lXlLESYFwS6IDSAYpICUoAslBz5mtMNMHbg2xP30CJjqSvRZa
iLovR7jaOqKxcBUkloD778Peek+RVdKu7uy5EomZSYR87f89cRqnUVqWoAReME/pjuBYwLczUOcb
lz5w0MCBx7kR0iYnbztt8PRQEmBCCjNPheq8X/qC6P0Dgaapxq9UorOhIF2F2HqEFrzyfoOApzOh
0tM59aWtqd4zd/5rfJuBR0LZTLrvcjMOxolHFciuk/wE6zQ0rESILAbxcRawTiOjzXQa7ywbQ+TP
VgqQpzqlodVAa9hfq236//SVsNq4XqO1zF0MJ+UBNauJvOb6054mKLdxLCxVNUrn9h2gKqAO+ffg
ocXQkB8aG4Kni0dEKjBTK9gXO1jivXeZ/OTYnnJkU8iNxZy+B+I8MRPLxqIqSMTpnZLWY5rHfVSs
p4FH/a94SLugRjHnWBVuoJbcRCDz+3bfu46RQ24wKk76LwFfScRokyoBcJoFa7kFlKB0fK6wvRSQ
PjuIjdVHWHLvKG2KaW/Av17B7yuUZpp6Pr1J+nDU54QZKfj8jcAZAS9z5Vcuod28Znl3l09jYuWA
9UQFUL1Sfn+dNv4xqZZER9XZOW3Zt9w2RQrGcvN1YQi5Q/qM5d/8Kr49g2Vwar9P7ZrDQjazj8c7
c6Bp8soFhIhLzsB1IpIRYTqtjTWMHFNWKbq+7VsSJsZj8H5cybVzTVnXmRqt7Qo/jc8ABsh1pg8l
T5z4QtJHSr7+RqAOjGuvPtcR/IqOK3NRx86gPN0lfaFAc+zxtdPchFpQ6aUrEz+rYKiWS9xUb+Rr
BTkICH8M44K3wySA+hxkZJQS/rpPFH5ReSpORc+N99b6c658el2EDYgJOUSMK78zBU8rEVbLvLTj
X+8+fcXG9uDL+jiqJxsyeIVumJComkOoT1efQRMxh6mVFEh4G4bOLv/cp8veA4XIx8RQSE9frEdH
4FWXivwXpRQmZa9pfraElXv92vXUE1Ntw9xKXKno2JMgcnWPYN9GXVxzx2em4kCd3ARXjC6fbvuP
t+HvD8STPctSSxCcM3rbLNqkTiE5VHkrPJfMjPawipx39LL7ABxkbltEiZ5Z1etjRPdajU2+5x+4
kOknV5ZsIWnW5qf8D0+wZV0k2mqhWDzO7KgHi7uyMOYi3pxlqAC7UTNIlF0aOozbB73iLNA8Rigl
Kdgkb9/HmcVt2nqIIcBYRUY48jjB2zAxouRQ93EJE4+GqqcJaVL+arCkd7z3Q4krm1rEGDURnmQ5
Achfd082EXS7rfTEXdlIHvX72t4LBgs3TfNcADH0U8ZCuRfUhBtAWY3+DPEVMhNZR6NAYUzBkYM+
XjDVYZuz0w9neJf+oZnqsU1CyfN2I5QikDsD0NpwFGv33tHEX5XT0eDG9QYTwJe7cgnKz2tm+wrX
GuWn6KB9sQyDFPqj4aWi7bb3wyDlk2Xq2s9cooCvOsrg/tIhtZPY5W+sl9jNtF/b5WTzC1X3SJIR
5sLXgxf8zJCI/sCpottiHP/AprKXHaDIExG7w+FtGj5xQLY+COYwjY0fnc2j4l+96Z+JgKn5E4/m
INVVW83Cmrj/eDGQ6zqGZ+J61dwTosW2D762Fxb6nLeTw6YtY8bjCga+aD1N1HfmC0/t6qEUUi4O
agrIxgl8Kp16ZRXQtMQUSY+d+9pey7REP+IwP10WCWF8HHux0wRd2ioq0kAHBykqtDrkSlO3t8/q
kjRiwpNHevcsy45578wkVtflPl4ocLh+GqFAzLC/2Nwon5CjBdcjYvF0xI2TFoxNQWMo+yMi2OeD
1Y7Jfj7Flel/UVL2HrnGfgg/MBIba2Koa+0dxE/jZEfXOoaYLVuVnrZoh+I4WI8W3FQpN6z2zo1v
yWAiIYOzBR43uqTPFG6+i0PVnQXdLqsHS57pkI6iQf9l7vgOSbFV4TCUWRh/UxdOCvT3wJIbdLvH
r4pPWlPDVl/G9ngB9jN1l0+azBO2hQdMdoUIg5/JWrwhMNo5GO1KSQ5sZRyMEkfNYb+ympOJDB6l
3pC36x2h8tDgVIcq/DW1xPgiiy1xfAF2S9GwC2fG4seNT14BhQipOKZZue0iOuKsCD79OXg3EoZH
mH3sLcCv/o8/g0G8fgrULz3uIF9CVIIE6zS3u2B0bhO5uhdlkVugxy8T8UmOt0nlDPo7UlRF9JHA
dRSgTqZq9AdwXQTfnFU/Fx5Mww1HZaI/Mf+1bUlTUzdl8gGREPaKn+zBF4JquJc9vKC/khjfuMRX
+NjqsN9RaGH1unv4fiVcvPEwoNQeHKwlr3EM6rYLEISOjJtI8llbs8qhoP8AivUhf1KH9PBfBgYJ
0KTqUAr1I74xcTiGSUI1NeENz+xQznIyUxoT0jC9hd6yAR4di7QJKM46g80F4HDWZxeIg9snfGDQ
W0mi/SzH37CqnqqGxlveXOVHqbHTP1oB3cbFbABmvG/ccHw6/mQxmKDSOh4SijBxKVwnrS3Iu6bF
Xs4u6Mj+dNCQn7Ijkm5oYq67+tVxvyLKW+5VkSx7PKikmefpkokMXJZQepmstXluG+/U7BNNzSQx
AUneKdN8k7JezqBLUiMezVvDpCxGGNiwBUP52RmrPbWl9DDohjedWO3tPLBD2SBZu36ygceULJ3l
jyrtb6YIooeDxOYqQT1p7ElcaE+nTbVFVmJS6zoM1YluZnGxHErmoE/AKHw/2Uy5jS53m0rLoMhG
JpwSa/lAtJ//skwAycXnscyx90VRk7luOtH0uHUT7WOiwr2GkrxNswFZO6nfLfQ+qYXAVCiyNMGE
bRqGUP9RYnCsh18fAy2v+jc8BGbCD04zfESWXbOCEY0tCcJ7oQhAIRsv22PuHwyA2O/+9iz44ivE
N1lOtTGgDKFUSdjJ8hWvcyf4X7B9ZjqiZG0maqIE0nphlzGxI+aym7NHFsFE66FK12vUnsZVHeRv
dYC0EReG37y0vk+JrnaXkgOo1HYpjLVJ9hhVYXHH7eRa9+HYJF35bCOFIgBIlTUWxYisjOCXvULQ
Cwz20WzIM7rmaXXhRXqiJYXoiTySBdAg1P+/451txxgHMCBw/IAQJeDBGauoN1hQ2NbwlNrY7y55
kt7UwIqZ8kS5LHu2cxYJdjabugHyPw76UnkAW5Y8pStj1Ojszutg1obNHJJPfKZR6MRBJt5VRqNJ
rb4x4Zt816cthWJUJNwZIHBs4AlJwFNjrmv5Nj/FFUkxk/Cj3ygtW9xts0zd6xYUwhk+b9SKGpB8
qzrmvJcihHyGUgKJcpZfmk7VxncY0TD5RFg3rIgwDo2PZdYZfT/hmrMZi5Qc33o+hUUWajBf1+BI
N3EX/g0KEPyXoVCs/sPabJZES8lZRVrzO2bLJFZSy0Zeqdmjs7NP9g9/YZ2PTgKjkI6Hl0gQ2kJD
J9ajYkwdXlvBB8a01frI4aSqiH2YYEYu6PMh0aQkZ00mVXSzSmLQRaLZ6u+l6Z+ghcWW7UZLUFw6
WTxnQmYB18xUCHZACu9qowwI6GCXHCf+IE2uduDVBR7X19EACgkKiv0AH2Ibhp3OTz6fkLpiNJCk
mo7Rp7L5q71Beq3j8mcTYBldKCcH06ExfeMDn8ZRofC0zW6tqzwWRzN989AiFrYtZFZtde9SDZMc
dlGw2dvGgxwm07p0syOQjsoSdbZ9K7PvRV2lIUDKkElzyQRDv9XWFBBJZiQf0i0lxBzGUJJXp+ms
VlnRGVxR9Xv9L2PHxxUwImSmJwtySghwQcwu+2hDNesqwk+OI2klihrGt0oISskrP9aCX9kQ8VfK
yFkHqurnxRqXaBC0xsdNRzzNCOPE3UQvNIchqMfjoD7xdAinDB99GD3mfE+BgodNz6Y+CGtQbH1K
QAuajLSUUzksGUzey4U9vly4/oM43iGmUuSaVj4yKUtrSuyN+3X+fvtOYfKP177vI8krXc8XAUzc
VvjE2caL1WhOwu49RTy1afjPBGI3+dbxo+jiVKjBt9WcTgoZMJ7Rm+/0Z5TA4BS01mja93g86EB1
AyABQl5XCgUFhAQDZLWVV+4bGzOZH1zLTYpL+r6pGOGP0ile2DhZhXcWw1fOcMwdRm+D3nNFzbGg
iDpy7cjwRJfb9hQMcW9EUye4BGttJv/QlH2CMolQLgKXeyK+n9Tfzp9+MX0J/zM7meptsRiuyjFz
2bkOmkMr2O5F48TmIwZMawmuWHOT+Xacp/MtjY27XdIXEZHxv6vUBN5YTXC237AmgLpNv5BtY4CA
VJN9NUZ7IX55Se0W+nOhbrN99XjpBNfzDf+eeEW3V6JYV5lhmmZS6elqbVBaYortMPDUfia6GHTM
BijfP5sHIN11lWlO8EX+GtWdWUUAckrLfOpRomWT6ANRHM5XxuBttfrE7kRNL81wZkeYNNFv8zxZ
Z9ynBaUEv66I8oe27W3Ca70Lx+9ikwZG2uLUpD+veiKugdYUY5Lq150TYZ5tNzLuWEEMA5VZH1Mf
cbZAdEAasb4BVRg/um+0GBiUX24Btj3DsfZyHVbtmOvJUySoowOhy+yud+ZxtPtOruURefykal3T
sFFGDi7cSTxed6ffDz+Nb0HZadVdtw0gCZl79LNDic07mlsyDepu2jPh75Agn2XIwgMnweCIgH/S
bMWTDaFe5DYwgTdXAys1/SVhqf9ojymD+PKHs7JjkfscKLXDnWpvuk1kH9/E2T1Y2iF1Iu5xE373
8ZWpljm9XKwSU5fZSsVAlZ0RgC2oO09nTwzf0qEwviMguYj74wdgo/PppQhzoeq1PpwypyHVpOve
JwMR80geQ8+zuDobhOy1efMMj7aEQMLFUxHZC7lgWo+MyeficB8w03izBys6pFLFkeGJUFUOQNpz
KRWObao/4W3TEIYZLcCGuoE6bc6+da/5l5pAPRHKYdRMPz3+01FP2dhz/EpBi7zKkk4rh+Pl3rT0
SspMnvopinrrV8T5d0fEwiOzAh0nWrdJEic4lZkXLEGZCCDuiAnPvwhyn5KJ0nSLIBFyQz3+1/JI
FuOm5uqPa1p4MaK/kBcGDVyexsEiCOAMrT84umsZ+t/kxBGQrtn9loOJl/KmJCZczZhUR5pYd8dY
BXjQjLYR9Kq355N9yBylqQfOkReGdylYO5KyG5PxjfFt0D+C/7QLGuohRsCRt9xyniA5KDE6oWdq
Y3/ZEPAoUqx7n7kfetvwzz1dHRs84djX906Dmi0xm+N6DVOO8pqK/B8aEVcqDa7p500vo7T4znUl
r0k37vH0n695Eo2JoJbTq2iCEagl2kKPDlSgFiH3O/U+CB24buLVbL2VG/DyFloLhpOTfGweeKTW
ZMP+pdi3JVVJZu/J3Jr2VQeuVnGcVRHpbIoOstOnNQecX3NhpiQYKT6YdaPgZDrSsT2tq6U7ARSP
GnGKegYuseniTj4B6acp3Aiygjis9be83LAMvoOZUhSjMRw/JrJA4TPORRrPHKtz4oJaNTHHbSNM
S5Ip7sra0BRzeZaJNtla5bL8zOZjciVbOnuUyeW8HTgoSYTJGkJ6p/iB9mdXXI0hHftktsd0xV6q
pUdbg7zl4MREUOzq57UfUxwhUqUlSf0Bv1uFQFFcDXhVlwNJnmoUV7a4LGnGlK3qopI4TGdXDepN
+fDgZfhTFDcXYM2sbxDSmpLvDwv16PKp+4/7TrTrZ1yBljtJ7YT1WrxKJDgEBXn5iBwiaosW7Pom
HvbEAVVGWYl6krNV19rChAclabys8zQbo7K32dx4IVReEPCJTMAiqdP2qp1zJ6FFBKJJuf/pHizz
1cd4zzEDQEN+yMVVbGvnxNaDK8JLhZWGXWfOSCsJdhRhDcpYyMRXTwOKnfDHeJOUjER7uutVIbmT
EpYd+mT3FYI68TKlz6Qb9oSLTTqLNFFX2fpNXaQ0blD99TxsDba9iw4VmGleZWdIjcD5FEFlCRiC
If1eH/fmJt9JPjVBcrXPj2pI5wpZG63RSC66nedVTkZ0XMrAqKeqMAW60V0C5JM92dZkoMZJVFW6
RvsbXpQUg0bvm3dunh56QLKhXOjZWiHaMVfq8TqHwXb3dY45o6agNMthZbJH8YaFpfOHI/z6GM/W
WQ/rBiJG1mOGjenq+yRleQQRLDbRRafG+6H7iMuntwQuRCjrid0YrCOkrbs5B89urfnDBWcmXmhW
k7GkILIh3QAQMVqJ38m58U4se3W/CK2AMqiXrGcwpvllN/wsQhc/+3ed9tlDXpfOWHk5O+mGxSiK
MJpCdS9qEXiZp89qbfGMHDRuGdKXYCWCSq3OvXTEQVVJ5Z5S2Lc+MCceZ9p6TpWD5ibwR0neItVq
oOUSZOP5rEV/93Cd6yTWLZBTSYqHpJkd3zRJyTL7Jcwutm/K+HpmgTm5ZJt+OPKivvFPUZs1Ae4d
7RYpQzL8ydUzO2YJJvKzGK44nPfxyr6cnaSXfHPJJPDIq0+DF5fTzbABNp8ZxqIHDsbFOvf8fxQG
GvlsxI6EEYpngF60g2VNljZfWmneT+Fx6BHc8ZG9TCboXr3PsVGR/dlFXCXfiAC/4f/frAiLIaFq
21CrPfifIS4pB/MS1FJkGub22wj76HjLkcZ7UfDTvfPbviCWx4c0b1yI3jwX4ZSgtDSCviwULcIP
2Lo9pZFqY0iTGHg95jVdXnE20v1a5zkITaTgu5lKbriM1DXuimgpn9j0PTiTN8Emdphryx1CICCU
08mF3kJHgD+z7z6reRLnbw6e7H97WB29Sn9D50LGja+BUGS5SAtfSW8PzCGvHSYBgK0XPNktzoi3
+IiN+vUArjLC0da+beO6jiaufWFpE3VfnSjns++6WtUWfH2pbB+x+N/6sYTb1EYfxlfTN6Ch5jFn
RA9Y+HGzRVNjEmTTWnm5ZsGg2GLwRF8/ASW924iiZ2zrBWs+mq3Nl9w4Awpu/UefsTR9N6IJhbez
gMg12liGRmneW6bToQJc9Kbzg5tNb9SpIC9q8AHJmzYhB/pyNYO5NgmYFoMamHfWBmh3TBDzQEEf
hjaijhFKwIDNd3Nk8wlHwbr22btvsBaCTHhlaa9KA3i8TIFgKznGrclo25AIc1pQd0Z9pQjrStMC
UWW/bzrtl5FoNx47aUaXxNsXmBmhVvPkaVBXN/wBFJVwCfvu8R4OfyLA8qhOnesuLOY3GED9CMYS
kWaHBFaLxLxpRxaL4t1kfkY5/mNlOhg1Ktu0HnJawoB+yqjgr5kiqm2hgXCmkz7r+LH6yQy5SQI9
5QUj9opI0bNrZUaWArGDwXNt0duWZavpRNP7kYRngVXBz+eidcoak3gP1k7b4t3JFnTs6SD9kQpW
fZtGuCyVxRI/ULAEmASe0QChoKjQveliBhtVN4NIL5XxN/3hvpMS27IG0jIUpSxzxuEKtCCDGFHH
AUkEz9lK1vaMo7MgwiyY+uJWEQ3Y03o6gFgI7P7Gg5Wy6WvZhbGnPIwiGNhQn7SUc8vgF0LCS2o7
O+bHpfMtYInnMmfa6GLdBYrHUXucgLpKD2i9xCRLAB1yLna9rE9QsuuMott0owG9kNnfj82ArgeU
Ylfl5jB6R3bmfwkSN047KtE/gULHFYAcK5ICix949V7Rpx98NAMcZDzzt9K8qB5v1VCgV8WF5Vh0
umPVBz8nkwf0N7w3n1eX6Kk5q+d1y3JQ7yBx4DzXm+WKkOfbo9WcZJ7fdjyAva3lKlDgBFFFSlK8
Ymoiito70ESEiPZD9TCayu/gYkAQYX5V6QDQHA5r5b2yFcwPvumez2J1x7HR7ii9ianczBfcEl8p
plUL8Xrcezok/Q/JTjh7EamykZDFCLTV8HGNnnksl4UwVSXqyUi7AfyyrD0luoa9VYMRxDY2D8El
ODYM303r+8e3eo4B4WFudVXd38kI5hYVH1wbBAA9H87vFsmQpNJAq69TO04hxUvTMX6yhDXOcVSD
KQTlDQAz7o35VybFcVkhXTS+7yr/WlVL68oTzji2sVRMLmfs5AcDOSU8nUmLFXfTGvg8SSQam4Rb
cM+3SLGLeSVCJqToxBoQlORbOsvGeYkmTZhaulnBHMZNIMa+/2P7ORFgs+vwOH7Dyya18cmmlgjM
Fdg3CfaxuNd6ZwjOL+xmnca1AZjqID2vXAxz092+8nKprJoPKwGYL6bIOdxQL4kFRBZMZ4qwDjue
KiL/lnQ/GTzf8HG+OaOWa32rC7LQceZLZWLWobVzGEi+6OReXc9Ufkm3X+4YKHSpQ0tc1SYcKN0y
qq46JD4HJ83Qkn0R6xzxbzypq/eDtfSWpXjLJ1c9mvJMW6owzp0ulWzoiHawxUgZQArsQQydo4ii
6HFkDzfASD4NEI2HNuAqXqUT7faDQWGvv7dN+aFAHh+oOO18jH1R0jKaaEl/7XaTRsV4qFdrduje
O49l4KLv6KKoJwPXMiyEbTHu5jI7Wtj0uPZ1iXcdCcgqM/ow6HCszabz/p/8Pn1xgr7csN6Dramf
hTlVl1aNOPKVxzcA1PjFNkJKtS9709UhYBVNEG1uFCzvyg4f0VX8mNlz54jHvaqmhaQCV7qxQDtr
60cQoF/q/1eRqgEGOK6DKvIZMOyCynS+4XyxycxExXDCapSVa2ZPKgDW2eWwKMMJsU2V39gEaMKw
usetb9ui7Aewf0uWoNSrCJqznarfINctIVz6AoYlbbuAvVqG/Kk1TzABtBAc2VZAW0Js3gZYga6d
iHnmW3AZb5uYWeSDMnYOA1f5q7s/x5hNj1A4CLQHW2TZco//sdzE5CDk9FXqXlbSyoO8g9oRXDYk
cNMU01Ltt1G5uTh35FjmlylfQx0Wrr0FPHHl/1btSGBtfTIgEmBeesgWc4IpsCpXjc4smF+xAcxS
EZu5maIow/GsVopy8/NwQwGlk2HJp+DmXPFnmuiR8dbxA4eNKMTuu48F5geNXYckgu7uW65QjoGd
gQA4wQYrwwu/hTKHoAcAz1Kqq2JLH9nTy9BOJq8y6ZEVnIWKBgZG5WwCyhcRUo5UfhZmmPUKJEUj
bMoTkq+siqCt6hr3cgnjk5v05swvuCwyX4pNsWNbemPigumZ9o3bFOJ2CsBIWdWBj+ORIQGTfWif
DVjgcu3KVcwDmEHpWOVIAmSOkngSD7PRp7eg9gLoD+LrGht+Fok6kztce8ic/jgynFk20Kg17uXM
PBL04hXI9DFbhlCv1h9CUr6LeOikKlYi+okGqrMlWkH1gkVOV8TxDD8AC/pdmxfn4OT3rD1Z2V+y
iRgy1QL5R23sBqKXlU5H3bdNgclmX04m2ghZFm6vAg1rxPNT+UgNZNVzKrARVIGC6OkxjMC7dMLm
GkDyCxEIx2CSTo11jpBTuJSasQxNR8Diu1IiwKmRJ0cSHwCG5GYBvjnfYvaZWrNy+eXX/wW9ZaCP
rYcfnEIif+XAi6TqWMYecs7FMP2vrzYyXWfmYRC1r90xw9zLsICja3/ZM23daSBwZl6kQWBOX4eP
YyMXkSaITcwkk1DYWGRkAg+2BhE1EYPEDr8g5WHqYhfoZ9u3V6OZnWnHnTPKPbC6/KDOI8QLj22L
GXvBN0EAjMYjzt29sNib3yl49kFvWOvukm2AppdnJ+HA72CLYZb5+XYWQqzxW8xUYtTdVJCUXoAd
HV25QZzlhdct6LhSMzkg/IaGo1JOEOn59Jq5ikzW9f4p9YRbH6b9yDFqA9gqoWeUhyaAeCgSt/eg
PQW+aGZ1VXw8PH85im+VSZWCa+L7eccn/pzTSTD7vOGawgNYXfnz/Dr9+XnnPFIoOT4fcu7iY+Lq
qVa+yqwsxDySYtAXPXDsgS04qvpY2k7GEfOhDdHPZ9TCUvv66HPgAgwZfHyo8Qxl4L+w5d09fPr1
C+GEIctj1Jphr6uig9AxiM84ipUc5vhXn4yDUIDAotzoh3lhOAeGrwltPwDINcS7iQ870QSytrIn
3F7Wp7vDRRyhtZhNRD86sxgcIPWm6eWBGZa0popypsLFkcZGbGXlnmOuO+Zc7XWjXp0DrfUnvv9e
4/fgalWeV0FTwK+lfeMdNq10vDSHa0GPkNJsUWIPtEunUwaqQZTZPPY+nkw+WGwDig6+Bc4Dawqp
5AydNlurT1MU4oKaQJdIIqxSijiPxez6lQj+BrmGwW/ZSpFP0TSchf60XgkY43apZv8KbofWnmkl
2ALPE2FS4HJHrlVMZPZQSIDQ3CvThtGWL24fhuUHh3aVOh0FFSKy699y3VP876bCR5/k1nr1Es8n
6j8z94/zZjO8jzOspwwxqT5t5vBySfHGr9SaED6LIRkIqvnWnEMtSI1UWNy1TS05v0hz3O4Lr/+E
zGtTqxrdKNBfKux1RDc8zAikAnv92W/BG8stmJ2XRexgN+aPKC0kTm8f84917BjD7ByO9HcWtXnC
nmd+z5PnVe+JWApdswwr4yduI3vb7KgB0EB7n6Ubn901SaPCXC2u9KpRTaeUGPpx3wJrS2s+OzNj
M22NbN2m92IFoeFTV9dbQDiYGG3XqbH2/JNlSLJAnDwn8325ssRFnWXmpav7z4bP7xvQ/8mb0nh2
zp1WPEcHJJtydCLzO4sNylGU2LMQC6rTDfke0MLgIvtMhInBV6BJpWbqk15eIE8SK9uJfuyycPGS
Iy+XF8pqZexBNcXdQ8T3VIJSK4G6oywgZtF9cpYuTM2w4JubEsQJnPtCSr6zbQ0tBHTFG4N39mSt
eFPR2DODKSdvUFHMR7g1I+pdoOHtJrBMiXAiOy9265kuA2+HzshDsRT3kT68HTTmBpr0gzN3u82k
ICsf5iewOCF4fLXg14KnXq4mry5Uh0wGhvWS/Wf5YUIJvd1pjsGkr3oCqjiBtKcu8GBn1l/tbhm2
P+YyBWzI/71yr/SMLtwryGTP+tWdO5VHAJJUUP1fChLFpKIMsCduxOpc9HiVZ1QXN+2QYB8Olfws
JUBKQe6NlxKsGeVu0f9L7jYZVAg7ovloZaQw5rFAFlUBGKy6VX4kyhY1j+7e6cUshV00K2ivDLd9
D4RZ2lrZSCOQzUvcRmwMj7eEJ9snjf6pZN0fK1B0984o0HK4y6eLf0aUFSkJZmOGRuTHCYoKg4/V
wJEwIrRRqda7JaA6mxMwdV1baMZqkYDrweGciAP7N1Fg4azYX7bSOQHIVuwengcvm41p5ufBRpRW
3adQRnBX7pa84ULiC///XQv2Vi9WsuUtrjyCYRTQTzNTm6R5eDeX7a0YhK85qmDDSUwTzGPCuWar
0dECEHauIRtzM2XHDnYeMrfoifIujXVfa/j8UgzrvK5B9AdfsOCyYRRrntBxBGD5Qt84do6Cntns
4dG10ZqyOD3T9SwGMvRW+8MNunE5kS8P/39hjae9/XU5738neWLf0s7lMjhkMej3+N0eWtSh9I5y
xnhhmi0dYHmzwVDN9MjnABIh0WV69tqdE4LPUFcYeqei2ZuLeoxEg9VylojzGlW/PBUXgrsEizLo
oLBKfYfmnI044xBdKF6D/5TGdjoAiBbiiES8R/lt5GG1b7nom0UDS8R+z4TWq03sIk/1lszpAazm
mtQXOI95BSBWcNFIALF55PMvO+sP1Ko/2gqOycNozJUu3wwCVlhEWPFiFSPgkv8Pd6qIQ5+Obaj9
6RZatsOpf+cRdXNRSnl3D2Z2Czb4yFHK0c/FIfUB51DvxhgDvjBsz2wAb+Xf2qHNG9jb/koXO5fg
XFYV+2H+9Sirnfql+pDqtuL4YWckShB8yB4+5U6sIPa1SptVSlSvXVZBl//pdPn+WJgL+sL8KZa3
6mZ6Inuc/iiMZ8Jq/iklZN93tzvn9h+pnI1IC6w1OgAKo/76/w/zbfSRRX9Sc5kPS+qXYbTfLy1b
d5o3dImnfIHARYS5mCEoKfEqmst7JJDtKut4NwWq9irmWIyGfh/LZQqjHl1zDzhqBEqfUxEMTGTp
rCrldL0jX4dG07EQ3Y/DXi5gdsSYVEwPRqkNfqMeMajwbDbqGLGnoAWBGcO37Ux0qrqqQaQ5niBi
ltWe9dYJkpE+WyF2Jc6hxrkOjVcEFVrhaWkrbJrwmw28dYddbk+FIreHei+PvthxIBtouz3ESo+r
/vP3c7qGY5azrIBptOp1TQcIznva2xWj7EEOBda0S6FlQQefdmTvJfskEMC1UslIiDzIIc/Bx5rG
XNetP13mS2rkBcyu9WapEXByZsdNXs24tt9bBDr0B3cyJ86MOei8pI2lE69LdCgw+ZXeICcylv8n
xQuac92tGhiUfGCiWIfz9ID1riJBx4GbpTldmF+zHKYSnu5C4H6rshSwjP1E380ZkDiC+cE2sxYH
JoK3nPZluL9wKqqSBBCMaM4eoGptARdk8gwHdvwqCYjACWfLdagKCsPXICD+3KJpc0KpFliQUoAw
cP78qjpC9RIztVNj64mr8zdniHnC/SHQFHVdxR1Faqp7tStoBw37hikAV6qpk7zlUkCuE4Ttxpuf
wYA3bhvjIec+CT1Bnykj0aEu59RcggeSom4NC4kCn7h8XzJnTXoFWYa6FnueD0FJV8JHm8ZbGTo/
AKUgKmvWIefBBkbw/phTU/9xfSoCRSPtGc3yX4pO+p9n+geWDiNtyxNYkyD9seOkOMPR0RrFyb0C
gM+afX8jTllVVt0fgTwkQYFA4Zo8siENQp6uwX6y4zJhz10OlkV2B43LhqOoZ3MmsMptCXpBhxsw
sVJLsNQzYg8wAcUkDKLWEabxRlkRaX7A7+POxDOhDTeo6Tr5+EYu9JQ7nIJb2VBXvaPRIAWqyKYn
NmdKB0vbEVFxHEkTmM3F1mTTeA6dkz78xf0p9S2Is9kScsuKdtpWAJsjxfznJJ2W/o0aCh04jCGg
g9u8es4SqIrV0osrU8xFyPvOKSmp9FPKACD1B+HFaM7BsiGkOYwOD3Xoa2vfQC7cyd9Rp6MOTMmS
kBLZeVyWNQFmQn0NPxeQdJsROL9i+ggF4P0JrbGLKPNjXC1D0TNIMpfQjI7TguSQby5kRCYgdseD
rm94kbjr47M2VlaubfKgTMpwc16D48ZmfYiPtiV9ab9cu9BIlUpEXmvKrBTFEmofdInpZJtoUl5U
+Oy3JtsjuTmNAAJl75ofd+T0Dx6ODGSrJz3d3B1uT8C2P+OH7rtaJ2kEY3H7u3SDoyXTbSnrIsuG
Tvkl8x0eymPkprMjgn+ii2AQvacAXFoPJGJ56DkSUH2Y5AdSnDrHgUAjhRceMGazH3W0Y7x/giYD
A7IGuSO7Gru4IRQjbgrU/6BJzv9NT4FYqPDk8U0UJCO+4lVyAcVaASFLlCnxellHQUPGz2lO+37A
qzvLskF+GsHmnJf77lAXm3c6UW7Z6lP+mwjBiFz8F82LOktZCVQe1gJLC8VLKfWM3K3QRMYhpmDM
7DeSJbIJ1IWCX25r/HMUHvoE5i4RgI33G8Yzoq9xUZbD58NQd8ZMvmjuG9clhNoK0sUAMEmpMO+l
npdAIcfjYbAv0Rler1yesrk2a0zrezzQtDMyhCYF4ySMB7wR4PnXDgh9f5i/Vy+2aClAjIs/cKrM
x77lcw+K08v8jojOfIxXT0fp8llaWJc6w2LtwCqCo4GHco0BRlGy30+632iWMJO317Ou7WRyFS4N
ge8XCmOwzfJH2zZuh+yFusFwc0Zk1hWL4JfYqDEhFeb2OtP42FaKD7NDKBpRzOlbS40xFCxS8/p7
vmLR/E8JiUJLHTXcaSTE+2i5lBelDMRTRsYfHxIWbQUCAYuwjNz3fUUps1+WY3emDwuLKnrM+Oy5
I+8U9u8OEXbmgafOqvb5LInKnJTtQxzg3pt1jGj6szUA5BSKDdx6CvyGjuT2lJUq2K2ApGeTOKsn
UirJqXDExg6xAwusSwiZAzrcJYrVg6DCseigVm8KpzjDNPZSfj7bj0JOcBXw+UkwKGrto3HAxyVp
HKl3OIoq0YdMgbb8DEwd4cLrQVaaNkhE786IsPaVmffzuHYskcrTeN+C4Vwo4839pGcNKTcqV7g3
iNQALZw4wSoTioQZpsHWD17fgKn1Ye7PVks8j30de1sHSjgISxK0DlaO6egzpvBGbVOnjy7tQ8V3
7HkcmspVuXzLGwT7srElNxo/YmoC7StadZJ8GDKHC7OZ0PTfMQPWol5bdEkLocIwlVIkLW0t0ikq
+EoFEsaBZApzKlLjnNxmAB1gT3xH41V9dw6kFrjEHruCsW/3N5OkgDjeITqT8knOHmDvqteNndRn
fibmp6LueveAIOnHF66+eiqDuuvUwpaZB2zrEp+jkBcDQKBvxAIcBxl6Pk8EA+Tf+Bs4QKGzEe1h
iyKzZeORd56Huiaw6IQ2xBo0vB2aFnqChP62RaZmA9rfPkVwtZq2l91p7YO8CgV/yXysKhcpPtYS
yl6lj9bLM3MsKbrktCkjipbBFo820ZV+F6KdXXttE8NdtgeKt2uFPpquNcUZCdktoEF0cugSve2e
XPJgsdfLYZXFAEYPi5Rz2y9j8GjZrE53CU29bD79fBaK4Ir4+kT1+e5KtsFajcQiIzWAXcvSVP0Y
5qb9MTBihJi+biH+7LMKVD0Y+Rm0Bfut0ioZsmOuWRQGKjMZNPbHIDp5H7YUB5ncY277qKZpnkzV
SJ4VOlCDjOWWGQWRSZng3NWLtnQ4CAyljK8EI1oZ7gGp6FX+VSO0cBUn5PDthjmuGnjDzxVc+Kbb
0vh1n3noMMWLxCoUaRh2AAsyBFPY8miXDV7EZMi915GdgeAFbWomwm8ZpH2UTE4sJw1Zb6KTrA+y
Qw4g2lPWkVEotGpCK4gICpL+iNXezi0CjlbLANMf1jo+n95opCvo5h7VK4bJWgSXYqbFPFoQgzTF
XPFtLv21J3b07eBVIaAwYGIqtNQODmQFVjadKxK46EFkXRYajMNm6gkFAe2w6WCOIu8f7ly1hJQt
vyojIYPpIO3XQOlUATcvAYLBEfD+zUOnPmTrTK8/tGEXAWAJfPQ2wXeaTvBqVkc1oqKhG39oeRuK
e9UZvC0fTjVD+776wSwxlB2dIwxmEwhxKeWwOipRRb0g6RlpRDBUF8nxIDmMP7SI/4QP132SbW3G
E0yCLVFdgCIBBSJOsB370YYqCjl6ZJcFPbUaf5cHRiW/of1IF+yzaAPeKkXaFfzi4T8JSd6apKkg
7xXgS/X7afA+sXCHFsED9601UJuOojqwqWAo7N7bZnfXTTAQ18QC+JhC3sEk2pt6016xTAhCl5tX
P/UFUVy4XrU78Qv7mcD1SvAgDGTzIo0lQz1POoJpRmY4rbbCm0IZ/Ak3aWmvLbXIFibM8DwY15bi
cC2+e8iJJXigRroVB9UtGe/8vohDt7AjGyZ6ODqZ4is856vcsuKFyGV9ZJQSgqts/o+Au3Ch6tbn
Sdtce+hR1ffEjZjLOKv2vqIaG4jZuHNemQnKiGU3kWXfrrX1l7CyGmZbNclaVPC8uD8GkIhJK3Q4
KFFD3ZWKOhA+f4kc9icSy6CT4gq8Qfmka4ckhSZSh/Q5HSIpiXC7VGsjvRw0J8FmMfpLn6naA8WL
FeATrv777GScdIpEKUtB+YDlNojWpMD5uYu/Ox+rWw+3/7/ALfQdEYgSNRy0TA6YirHTzEoOLWU2
gRw+0FlDsExSBpm3775gbFBjQc2jGC/Qw+UfX2JWL/4H/IJSf0mnm12+gAZUcy87ISkTtxKLkPo6
RQ6uq8KhDE07fxZpvbbjOZhocRaYlr2Sfp0cDGsNbIWJvEZs1Soy/x7FLVNF2clKyGq0t+Zu8d1J
rOuw77zl1Jp4KO+VzgVORlKhRDMVXFmYIcFi88ajL8d8a7YWEBUDxzkIbp65YqU+Ep10Wdw7qAcM
7y0eTa8zMp8ljiCMF3j51t0RCxtEttJAaCBZhjLgfVB40yObtuU8Vd/RTLmNdVWik47q/ZASIVHb
a3t+9+kTgpVUnnG970EYqSJZgFIbUxvQgCNC80Vaq3vDVIB2/S4tX1CbmaN0/xmAiVpHyzRIwLjS
PUU5KKTmtZLSThFcjS86s/AiAL0uWAEpblv4+EHUDZRUkaz4KvQ/GU/pzFZvxbenF8QtvB+9WB0c
MJzkn0xceXloQEVqegFY9CkybNsh9j1VFHGPUTnyjsqHHThBV16chASQuYuQOTVw1q5M+YMc4sLL
jRifLA5tfsa1EuBc+RxScuCNQR/tiGg6kbIq0+gaGu2o4eIO710ywJaJs4uzLwHzA+y77H1hEakV
dckukVx/iuAi1mDieezPyJaUTouhalvBhpJSkWvfdXyEINFNm6LSnjwzwxGI73he1Fu4+nzL0sp8
jEu1/xb5UwtMS1+uAJfPBXeJ9QhougCy0nO2F6EkMMsqGrZsS427avlrx/aGG3GB31lrLz7JiIBS
mPJAjvtjQPyYXVKmV2KseaAjUftMBQg77RA7qLjFKYdBPNjXczuM0Y6Np94J4PvSOyqtbVN0evfn
+/Zw1xL2t+oqt0Oi4lkSW1sCAYb/2YyeFDDbMPJjG+pJPg4QVrwlIE1yF6DSwgydgJpVgiLovplK
xDFi6uq2MT+AsY3S+49mLHR7HizQ9TmDOGMalyi0xYa89UijcmUIGkjxHcHs0JTc08EDpyT8L99D
sGWRCOw+6BXRoB/q+rPqiYUV+e2hGcS6vspPzxVlxlK3pu3N1HPg6PD0tza5sO4Fzqz8zP00KeWg
9VnUAEwbW9pBSBmiBuR39mabRvNEj89HY/Uvqe1eWf7SPRUJhRl+MfXjUnXUcdJqbTB9mIUfCAgz
V0WBykcfMsEtYsZfbauD76r/M0KYP6ZKqc04FqWdqcLk+ONvX1WbMQgVnwY4gFMbNCXBwuzxcdMN
04joQpPWSdFI4aqHjWiR0MdE5VqpDTfw/vGEkYz8mR1iI9XT9lHc293fNRtbFC29shxd1P22Vs/Y
4E8WCcZO9/HT6KnRDHVR9lIHiAF4ZBOHrpuVfuR/kM4Sxwgwey8lT6GbuZ5LDxKyaH3pMkQLiejh
Qqe5d89Mwqi8F/pJOWjC+FyRAVlIZ93yyc8vQMt2OKR5+LD842maQoBZvkXIk4H/Vr+yGj4BVwF1
rWY5FvVyH7ruhFheBr8BGMvNzP7pZwCe1xsk0BlAmWaW9XP8Pk6kQFfGvVsflz0+7qH6SE5tcRt0
ms9EN7PuN6tn4nAlkCE6PkmcDx/sEuW9cWr02IppPZ4FoGbHu1xtb0YRtQ+IocGAvsYwi8Yub7C3
0VXlLZAmo3kw8bXH1Lp7BzwYAOeX1siC6DGKgqqVSq91y4IqRhOd9u9OCb9UUw3QA9Pxt/lbQonR
8EXODkX2e9xcaaiafmJZK0/mnQWWMYNQdVBa6Relb7c7OJDBQTMc1SNJ1WWvUJ+fJe3kPw2Th3G4
cdzufI7l5Z/ZB1ia43b4hBj6Q4T1PuAqbqPEgkKUBhKsbrN3WbFaH/DxLAok4AeYCTHwTuoXwPdu
ZK+JPriSXIMc6MHTaATEJt2Y/0guSQbMqMUc54EMwmk+HV00ArLuhlfLRmZesYNi7iUXFlQ6JRMb
hCGL0tYYvzN6TZ/HbkGzxuWQLrxZ3sSDq/3IOM8qrYXaFLOJpjTY0NiYQgB8bLUrsW40dzWYrjh4
f48GKjoZN0aPa578B06DXWcSHEQ8SU6kABWc9yWCqY7v4ItrFzhy79LMN7NEiyI4hZyB+YsWRXp9
mpdN0Ts5mIoKTJ55GcXO/6JeNOfkLn30Plc3eHHU+YsZtAueMYsf/hd2yRB0D7JR6cV/yMHikEyQ
rpL6Qo+h0JqFZ+FpXRQ40Td5kgKDTOGcbukEjzQ3xONCp2fHMG8bE20Ho+VUPsQBmhLQ5s1beU7t
zoc7p3/icuArCBCJ0p2faLq/2fmLTWTNgiILoFMn9xfHBN3TJSJ41ZGnBapdcd9H8/SKyrrLqikp
ayWLxSi9+8jrMdv+aKF3tkMyM4WbqJsmlm5PbmEibn/BjxZZtwtoDrkyKmBc+1/8ETDxq+JCN92F
mmJeeKFRy+i/Zk9hJggNj6TMyIMSWhHT/HaiigzpNTe6SrIiVI7TtcAsG0kI3H2Etm5Bb5YHXXY6
Owu5LeyUjWdna2HqQrze1lnkpwph1Jhwx6yYbb4dNgtjUJplD7odwmMbqFkGpXM0kz4ixYe0REZb
69vi66QzeSkszrIf1oJ2LGe5kCDzABKHg4MVaqh88FmSyLo/UoNCC47HoUCKpGaCScdCQjCG6ktn
NV/PJdqNOQ0gMvCfglnlW9XEOQ5uWvrP3t92AfsdmN4hTOJpTaKMN1Zxi+s0qByvB6a5sOEfH5wf
B2gqf73yruF9w2R2Pn//BDD30axEzb8XrR4UndtgeKfnkO0qH1H/TNKTrGmw0tI2NYaLgImSwpCW
E/+1a04LfOE5NCEZkd55B3OtPlJl6CGkSnufO+B52Ju+sYDcEQ3lAW6H9KLOOCyqTRdppemaWh38
KhrPMP1xSDG1xU2Td0oxt+vdM19KOKanpqVK+b5ai/LMOsk4jJ5MKwOWpd8uBsgG2jiMNwTK9q6L
gmxA8mrkuztmDiOUdCPEqONnKbOrFgHCVIj6AKuqWj+sqNlSh0Tj11ws+H7qnIngpZdm6QVXn/Nt
UcE2z2Gylmlf/WoaciQAnQbE9S6yJE4wLwlChjTaY83yhOdnKmBbd81pLgUzvi1bSfGHAI82vVMq
aTOzBCHmfT4k5YEc327uWAqFHka3fTW4XFUZBjZJTTnUlSOqhm1irvSNzTDzYSJbDUytkjudpIMo
0A1mOtH++NHEt6KJPbmkpqdXh0ikYINAlycN12V/fdvj+MxmEpIXcToTa5CuiEG0ReQVvBCMc71w
XN64gge65lBZTMXsKwY5dwtsrBA58mYa3rczd+PLuRfK/GzPfNJQ4Vv2s0QZBfp5//63RYbOKb6I
3WpPnzXDqMHm3QwLmT9Hkdq93xv0dVUiiXBdygR6BpKtN3B7xPCOqwUndzr8Ker7OuNTxCvhzKQ+
lxV/KNLwcbubvs0psUddNA0hCr0jQAcIWLB1YcwLk1r8Ryx4pRiOqiDJ1OE/pqDZ5bW+Tn6kDkTk
RqmDZgiHnKH7WVWaiUsFjZ6hkVgaOUXVPbTGWoAb2BueCDXQh0O7SefpmOKecpMaJVaQa3L75SMv
be22oVpKIeDTTWx4yPirOnwge9a/3RXsLRmxfTTG9GN/f87WybMz2sMTHjAKqslDB30psfI9obIA
NuRe8s97sdkgz3Qi/+LnEFqaeWDUykiB7/QqQD5c3Nz/vlF17m/avNHt63EEC8geib4rZFc5lCs1
SvOjf7eTO9XADpfTxlyNrtJbECprKk144K6zWujd36HH7M70+iNjZTlXkNE8vBDs0mXVMRroA6/+
MBhkgFO3RchI856tZtvbk2geNlPM0RuzqiJ+ClEwBAwq26zvkHkUI2/Gc1epobFSbDhiJpg86EsS
huNtoEp1UQugyi3pifsvVHB9Pi+8T2C/st1ywXJrfvX6TFAj+CGPia5SEoq+AbBt0FznVZfvXfcE
3RcOaE87QXv/BqxKfisDTLw7El9dHg4XZVcdQ3qChjfeJLGU9g38tgaKPPJ8wbgvG6MsLwFmJd5F
iDsnxd2yD1VGrZ7D+UX0UXkpSA6+Fc2146sp+wVhi8GdzLkc8Sw/mu3n+4fbbDafmuvWhjEzkkSy
nTm87cXW3zy++Ylfb7VMaLivJm3vqiNprwzmVEqjEHMdvHnkB3vzl04b31NoB8QFvIkKu+qW+FZK
iZRAYGVU1vi9BT3MH2lZkNqFDrA1kdhxF5MxI0x2MoD7VZ8wjrW1ZA8RPzwU+kSvdrtIKLUmdAjA
iBeYxOzdBFK2BDAVQU3LaK4jaXlZbCin0f1sJdSARSCZabAz/4Xn4K9L30SsYV6/SiwTKsZkxxYt
U+FbdVMuua8AU0N4GxHrDXOYGtnqxl4ZOwPOk+mG7UFYKUIqNwxb0R8bcHBKV5IHJbQNLohqLLv8
A97WtObLXI956TF2KZrYhGdkF/aCJFFHqtWGW+QBeT5Jm6XKOTu+pg3BNKownQF0PeN+dm0rbT2p
RaqVw4AR3HxPX46k0/TSuTxKhxZM1PtK7wykPFb9Yy+Dtjet7/Qz+acOWGsXu1d3CS0FJNRlSgit
lsbIpX2KLjkihNBaw09x9bUs4VsSlRy90qPdnTXZrorM564AeNE6kmhNMR+1v3/pOJijuDeV6NmL
hEIROPMHSrPTr0Pj1OWekUJwqUuX87TAvQMKOFWasWQBWuHZaDXhNO7STmGd07rnoq+1Fs0CNXIt
RM5bVUMJOBwDu1Kh+pg6zgZ+KNgIpljloF2qyr4DBxs99g3SVLo6qO0aH/z4io30TVHk9ToKYATY
HtnSM5hy5wyt3moF1fEvtW1+ud2fznyF9Eshldo9pPGGtLYchqYGjsx9dIUcqBCdD2tmzwT91OQE
TGQ/VBuJQzh16FOIwYLXy8IYFqQEdp9DR5LAGg0zVgnqkCgLuztOjOSX+W3gTqdQrCuJXBzfKeyf
YCkUNgmtPTIwBcCFw9GtNhRo09XVJJlNJvQ15MSbin8lWEQZndnhL3Tffk0uGdIi7MyyWmPQq6xU
vnuXJB/EMBFOmE6QdiOHV0rZftf33r25PR21tqgEVGExcvVXT9L6I/QHCaFstMc0i5eMBs51toRl
Nvj4mAcW7VsYrj5bezNQwfadCBme8Q2QrxJaGrm+zdVWYjJXLG2peJy41CAkwVGoRVBAZHo1b5aT
WVGN0cMI5/Ae/l/ETtZeybLsZcN5Gvw4cahdltBKaM8IM/xRmwJXtJjH7jCFTvdpuIOCYz7MFylI
IMbTY5gkS0QfduZNrf6GnS84j0ZifYJpVS7vdadlomhfJQ57zayKRZ/Ie61nOV3ur8ByKB9vUJbB
zWj2XyY9vN4vgBa9jsOQOdLDveGTmQbG6YL2p6Yt9FfwztEubuVQD1DU0PQdExb7RYISAHpc4xKw
4D+Fk0+CLc4ENwBStpMQSgdfZmEztyofX665peBAHyvf6xz/tnDlVPWhspseE2aYuIqTJ4l8WTc+
TrQ6uLtzI0sb0OHa34WZiDQ4yo48y/M8LwDaQ3SAyRFa94PY/Utd+RTgl2BnuSB8GUc5CHag6cp5
nJoDUbKhI8PagAUS4qaHvKHChk7d2wsdQz+keUa33RL2EG5WacAALFvOdMSdJfo6Z0mV9v7Q+kFr
Hey79sv5dd/yTOCgr0M7VUT23oh5snpk8avuf2ozcgDFm/g8UYEuUDhv/nCC3cVl/hoiuRqruli7
KCe1umy4hLD1IPh16WjDY8dQN7hMBhiMAqL2QKRQ/XYXV/5HREidspqc5EcXAXbCejXOxqg99Tey
i6Jzag4YY8Nn/FielbL2bp0XxtuGU4t38o9u1+dk5TBp/pLl8jrCJ76WwtlLhp9yDX1cMFhQq4k4
aVclbI/4E7Wsu1krSueZW4tPh7UlvJWVSW7KaqkLQxT4mIUK0BTggFn7Nf4aN5VNq2m5cLN30c6U
gp14uvmJ1nToj0aTvtIpu/lUedzs5RjOekkAlDfQ2108q/KjqwKgRs7mxVZk3dp4GhoDih8mdqNZ
q/n4fNuF/b0XdU0K5NA7QlnC/hY0Ne8daEu+Y9F+7TzvH6oIR2LZHdJSsBtM5oj0WX7szEsmv4JF
l+w7lF6N1rXDdA4qyDUd+fR86mZri+RnXHSqS/KF69/SwfB3vh5DLKsA1ZtDuAWJMJwPwcoLbjGb
605qud6ZM6TBflHZq5jJqVEumjRLFT/oAgQamDUsQKfVu4SQYtwcQxw3OCeXUtenRTicEnvfAZb9
sIaIVplCUUSo/BnZ0KAnGmXvOV4v9kWgZlCH4Tb6zOkDk2Qm37Czx87l1ugV/UcR9srbPcHqUVrV
hwGd158OKhWZASNJQsqFJk+fg+MEc2cjLFEwoTYDms178TQuEYGnHY79GZ7EKzyCFPxRwcXewPWV
UH37ozbWKfoaVEXWTBWrUE/deGLMXypCNmgZGfns+BA4zCFTR4z8hhGT6t/wuLxHZz4D/K0flytG
q2zAbbfUOdTXTcmAwHS5kwIu5pbZwrgLQ85GPqjIq7vWYQvVZCxpyuoZsj1r8gf/Dr9MA2CLZHLg
OCTRxe0aN1Y/jBg+rzNEvhzApGZmV1eGYgLZ6YozDE0uVwdg0+aW8tQNgXt/yyA0rlPUOrOVnuVf
plVRJPGPpLhxUngvWMit4a/W/IQKiLOyulHOWsnqIp9XPy3tkYP9X9z8OzLeJy/DUhbWbPcJVwdw
VxfmQ8o3SaliLUnGPAsg3wrnzWSIDFES8pC18MKE8QXODLl60Odrvynn0OVpF3+QuK28ONESdViN
58bNtGDbMv6vnp5CrJZxeD5stj2mQNSZYDPIlg4kJDlDtHeVc2k3fcg7foZfcXp100pARERJpX7p
nf0W1C4YFjo+0oIJHr9g/kZn6wYQ5lkfnVh3WHNxv5Zt/x54DMg+kVZJTTkTUBIR7FXEVPvUmBBt
NeJD0bEIOwWH6R1IApuIvAtpHEuIYgwdNCXYVdQ58llvHQLaW6rddgBK0vlwZN1YcsOL10BitM+w
Sgn09bZBPezXroFL1MQtllLnr+6Vx3+aol8EnZVdUKYensv61dJXyFDFOmsdkiSOxIPpQQZI2j8v
hA+A5fCYHP0KCN24bUUBG3dZh67okr+opUb2/dV7kRftsiQNpUiC6pm0Cq4E90PS/5SPLIPvb+gc
qWmHZO6tTH1+o1EiXt0bRRvY6bMJAXHRvAR1YbOAfcCBLBG2cOG2CNW39Z0TORBC4Bd4BmlviM3c
pO7BrMy5IRXPlfZfR2dDqeMQxq82fYGeT678B/DZPkjcOs6/gLFURhNDKmThsqs+R5BsE658ocx1
+7lzRlHFsoNT9/YJorOm8GJZfNNogLJ7HM/MVTKsS6k0qzue9FKg0UJb44VUy9w0m/XcPY+CVjps
wv5/jQPfqURPbCn13wKSxFhlEksjT9I4gM7iF4TZErfsJJiz+2PgqlKoxgSc6YJPirwaXLNfXcdT
so0jJ7qP+CmMuerf5gi7T9u1jDr6MsxkVK6qXwYlc6aUbWRzkbUnGg+9oLDHeXnrmU39k/vgs84v
jSt0PBKU4/q8GC0OF15sPXzKwW5SOXslql/L0eo7hnI2+A98HTZjr8gla7o+Y40Kcdz2LjHrjgPy
MyG3FNcV0MEOFqyXFjltSP12OTM/C2NtHTJk0lydgeqpSWjKofXYLipcvK8vJZ98Hck6XZGjmJWD
9UOxjBkQgAEkGsb2MEiIzWm7YQpzcvzJ7bb1iypF7PaaqKHJWIQrw0T5ilv8U2SKTRV2qiPMQ4et
FqOYrI47SDkh102VofCfMT75F1ur/XIDfGFLDxl0ehSCxMc+C3F46HH/3JGsxXahLW5MIV4Rke8G
PHqUiD/9RXazudIECvsbo5pCG3oQRV/JRaT1mSAlq1+F86cWE9N7uwms5OxJyWdgkx4PcOrz64XY
bkZJ5Gt5BbAwPo86Kmn8ST0YAj9lOKJizCoNuTL4jG44+rMbbgcd3HC4A3Stj8SPePRsjhetPvVC
WytTeqiB5hYIFAB9VS7tt3HXuzAhFUx7de7xo8RbW9CommYv/31/cUj4gFGqg82njcDOItBgucN1
ks/1AmOVWfoAUxiKms7axiIvMB1KsZjnscJJrFlta5SkD+Jalb0G1j3Zf+cQQv+Ye+d2Khefzk1X
iSNOGiHWftpRMjd/acRAIaxwhCOIH0sjUvXLoHl+qKefZ1q4xRXOd3b0mSLC707rbtd8JrpJigbf
YPNPoswNDpT7dvAeG3abYqFRzW1/fMX1wMbYwtmL/+KfWLwwNaVs9ZXTEjAtGzxBEg1bzNNWdo8a
JOaCHDimw7hGaAjsFVNOWHVF+97yaxf1eQS48askBFfP5isoBAtKajedStj5+3qVmPkk2Xxl/FxF
rMvER8eKwjwWw8zLL/7ZCwO4AbsvrHYoiQX0vFMREn5/BrnI0WTmKfWeSIuj02KW63CgJs1hthPZ
kKSIui92KTjR1XSwNDw4aIRyPZF8VDCN+p9sVVU3RxsP8M2gTedmZtWyX8OAoUH71Nv5FyLrQm0w
jb6J+wIcL9aBK68dOGhyFZa7yL5IIbyviK4rBNuFS2wfORuY16H+7bPMZt4WLHKZE4iJ2qneCwkM
8ey9x5uaKJq03M3gYytunjvchGTafMldLYWAettxiUIn0tYOeUqMYyKwImDdPyTLNc3brBrHRXdV
yyYcd0pOQYtrXKWT+/otkS2IwAAgn1ATN1BN8+DRKzE+USO7q2Xyw0qsPIyb0+HCdyCS6whISrz/
SNGqyjaJhCl8FEk959fRgHYZ66/yJ+creZYr+a0TpKlMpB1FAfHOXdqqf5n17jNUTNd3Lsam+Fwm
diK1EMaP+Xy9o+0q0PYPOyQ2yzawLVT+UatynXVu+kFd53ikf5pPfI0TcrmlpGzPjyz+ivkh9QUS
xTCUMB8Zl9oHIRLrt8+tyYswc5xyeka/X8D8H5jgG9syIUDsgspmBQOeyNIir8nl7VwTd6IgcfkR
JkYlLvnK1qjl6C5zI5PwkIaHp76ucpFHl8qh3RCoqttHwWzXbF1fXTxJdaFDzjWibkmx7rQi5GQQ
S42tWUWB8Z6M4iXGVwiBZ+DspQiDbAySVmiDFlQAKe6ZAXjUWm6h2x+9x5cLvMnuIagsD5ZBeYxO
dW5qgyTOM9FP2hhWn6CJp27EFKsEoldjXtmq8ewf7LrFXFd6ea+vvWZxJ6lxfcHnth8FpKcDtCbE
DJvpPm5aDUCuLx03mAWYDmiQ3F/TTNzFQS21OhvrtZfxeg/Goyafyxccwuz7mXJNuKztCFTwVRF7
WWulbn/i5dSYDpEbkOD7bbVclazKviGykbVAsyKg2WZSRrmoXng7t13KmxYrau/foJM/DJdLpA+a
3BjFYPraCh7zzsAC8M+JyF5aTOBD9JfcbsNytgfEVsGB21KgdUk2wb/QFvscjdHM7M4K9sqUCwDb
AW558d29xnFtA/0xcbni5GB3Jz8Np00bRPBmBfNmfWoVikyIXBykZ9fviu01ctmocY6l6CqbEhQj
C3oqDo8qxKwV/ghU2yNGoEoSZd/nvnbLpX5Oabc/QT2uzmuPk4wSmDmPQdgPu5U6SXAOuzPUBeKj
01Z9KMbVES5Rm4tjUHvFv/RIZyaSzEyQIY8yWVgijxi4ruSnAxMWZ02sIpH+FFXUmhkY+Bcnb8er
3In/NDr61qgBQ1BYvgKQSz0sliZjBOM58HkHxRo7D6GgzAe3xvKrItB8206dbyRqyRIs8yYZiswN
CgdKKSJfxpQZ9qS3vK6+PomMgbjE5gBzrC3bzUOsh74QDqKy+07FioiAfWlFRC1Bg80Fk/PmpFmI
D209R424v+704Yf6oueWoHVJU+ovf4Jz6DvpW0R6N7lfeGzeqfvltwo4HXaoTPsQ1XPSI6WZi4we
PtuUHAZEeQaP/e7+gAJN5N0d6z+TeHVURJKBBqhlDz6/16UCF+loAjhJb6d8qKxrSXCClLwsQZXz
IEMwQCJG1BjW7p5sm9/SKiApF+EKktGB2E9ejQ1l+FZsQOqwa9zURF+gC4FYzL3jaNQQAR8MUL9Q
ypWUFN8BC0Wt+dc97FqLoDJMr8zNpqoZqzszE5Oipl9FDFfPI19U+rQwEl3BzPiUlGSxDvR/i84b
Mr9xdBAGyTcBVLi8erLhqmgEvWoflv4YhcToIjaNYzk2OLb1uPN04kHks4xfGA+ZAcrI2Yfx68e4
b7dvFCBIprqftfkA9AhmgWEPshWLsGLSnilaSX2+J89aWvDFkJl/zKnNR/mJrzp8ZQNgozfCDQ3R
2mfKuBtInNvd2ToHsr6ZPSVWBCEqk5SOCy2wCcjaCuhvD/xsVJ8w7pn9nOHem1NXXQtqEpn+nddl
NNj4BHgT0UwF7iIU5KhM+AvkcnasDIjD7Mz2Ow8SeECiSr594j1SIQSlpnWa+bgjw32MVAo/ybeM
imBbQR/8wNcChOEfD3q27k0IblCqSjMh7VfA0eTXzTn+a9E+I6Neb4To6TG2IYXEiLELodWp2Pv3
Xot/1kyqan7uDe1cSvyrUhI24iDqWItmaTr4jFdKKOLuET61UM80B8HCbTeQO7TfQARYVwPEYg5Y
8ST5WjsWXOweH4/QNAGZVdNnJZJUqEYvbS+vhg8qgXPPP+qyC6CunH3KfnwX8M6sH9e9g7oifnlg
RVDU15ZK/bj/gUYstRyW3St3TkJxXZlXv9EDKFMUovnGN6pa+ogO2TyZyac5SeFHxwPClFS1AYlG
qKx+cxu3JYuhjELHUqmANVQa+Nu1J6ZbjZHYcexmP1Tbam4VvxL9fo7OX4Je0f/EhvcdYz4iVa4V
BP1N4pvfEak4hNlOI11AkljxSMUSU4ukCxdRMb/oOWHke2Ywmof6vqvAD6AorRBt/UF6VqUU+igi
endAT5qn284UZqFAI4zYLOm+28QBhMsPZzUhWed/C+jgAXn/VDqVZ3A7B9nWTchUeffzl0bPRT7b
TAg4HfRH1liW3iTzOWfJU4/avXUn9cSg8rJ8pbS7JA3DmaQDzcovytvQHLcPmlsT4Pc+n4IiFqUr
OrEvyIzR45DKqwaDyvv+QQJbQDqKCHUQAR9MDPwRBJ0KnJfdiBlOneYntiDasZAoIEW8SWmvKwkr
CD6Uf9JlAZcVXWTpHFqZt0o2SAFLVIaDmqSW/gKcCPz/pNpQ3gITa306fhhIB5Ud+/6b/Q9KqrUP
snP4v4iHIJSj43hLPuVbTOKyyG/K/8Z0RAnp7W4/y3/JyJ6RKE8w+S8z2P2jSUvCTIbDIOx1hVYl
xbsae97grqRJUT5OWUoykggjb55Y1TAv60j14dk8swKHOKBM0axCdstwO2A7+fF+j4o7N9P5G53E
E2H0y1niY3WfIP53Fk4eQDIAKi5RCaGiO9qGLi25ulIXOkiLHy0IgqspeoT/SUhtC00aSmxXAqFU
BCNkgJi0M0fLLXSWtFlzgNoM5kaFihb9FaKEcQWkuuMT9eY52G4/A5kMTRbJRqnX0cYRkq3tBWJh
zufKnjfv3V5O1qCt1sWriYfN2dV8XpB1tXdciGm7ys9lM//ydFoYEd3le7TwLdAYlX6PJiKhwbXL
n4HQQ79cHzJ26Ehke+TQzDtrzeUzszaYjKW/0tLq257z9C4nHLP9MMLQxeXMUUoaPay/76bkrX/l
nNC5soXoOCR3+0MAk/hauMjEFyfMZDFW+Y6MbXeY4PHroGBvN9F3FPHCAxTYrqoDJ7ApfX+VKE3j
jNlwqMAaSL7l8w0kfq+qZ6E717we+LlsoJWmdIn+ut+IKT2x2PaLDD2gw2k2ypqw4HjT03oAmgSn
73Y6UpRbxvPY6bDI2w2teem08xRriT6MrKfN6sD4zf0o49k8L5fdCgfmLDyZsO7IRVycarTLxVIu
WeNlzAIgQhDcjwauVNmSUCRJrEWI8Ne1Jhu6AklyJ0A8mARVRXohaItathoDhlSjXgoL6a0pIhZY
KuV9yELEG5YkqWrkXKVXOpp0fUksdJ8eSPxWJE0t3iBDuRtl54zjgcp9DtqKHYwgXlL5rdiTunV7
dySWptsrIqY7DXP7l0ldtWh9fzLxR/6Y52XdbQY4d3/7pvQAoEAdm11LS98sz1Y4nBJTz7mWem/l
r/CWvgmDS6qtPNfWxxYsHxB8Uyycd6Kj5XxFSFgFgoUJ7MCS/PiCYku3wmQpzsnYE6152rJobOdS
gmi9p2k3AsMmRur8BbpMx0+SpBm4hDNU8z3Lj3PnwsFnSEeQHSKf92BiUnleGdhtc7LXcwLP7Bdx
3oaNnY4jSfwQikjljfQMGT3jIXMR0sQm0O9cS2KRXUJP4dcOZFjOsdJkgaNzVF4LB7nD6nmhvqp9
1TnxYvCriXlZNiRlEeiZW4+cUkMKXRi50hv6jXDmRCyVt7qzNaQUofHcKPYaR4DoqC44Co3wiq1Q
rNbZhfZWn+SrtAqZiNFdvD6QhKGsxS0l5VH8K8sYPBYNGHdlNkpvoy8AtF4BtsQLp7Tsh9oLbHhW
9S3es5+qlIs34j/ymYYMKNugNaeLd0KGe8+pAmsCyvHE2uiekgGMuBO226ZRuaUo3Fox33oofGk8
RegGfV+mgAo3x+gy1uf4s/3QsjagXFOBxAfHcP443/Ew1UEDAoldZa/ha6zLAzNeoqNCBxkcQ4Ho
3FaTz4vRVc/bGRiFtfoJWDPCg3f+7Ot87u7jFi9va2XOe91jYjb4mSZ9QbEeM5Dx7K2kRlcjADKf
6NIsQkmsk5VDHu+4tNQf6+Jm7IGk8q/q9QOS0+5huA0jd5hQHeDpnz9azUTQcDmvjhyBcP5ZS++8
6XNQYLTdpsgam/thWrBZ9Vf4tdYrTFrWJsG2uukeruftxZ9auP61zAsppz33TyWUuj50ePNV5fn/
/tTEgOcHCd47LZ9S6GNT0R9xsf3Ipvpnie4hx2vpkJY3mxPP2S6haNNqWT09dHZaGGDkeTgYutrj
wFiC331qbLEQkafzmAtzYPz9704car6cSkG3CXxWlol4o7SynsM3MfXfrT0moSukBpdpADe/F7Qo
IZd/zIakNytUj5/acCveQ0KHFzLLg616W6JVe2AduJZ/ik1feNdUrW4OvcghBKAIBhSInW6eoHft
Yrwkj5mdprlg5nPSckQryqQ+gyavorC1EgRIyIefFUTxHC7uho+IsPiDQ1N684s8tIdfGtVYtYlo
VsxO8YQmzO18mK7vTUzSp0X0g6FYgvKXam/FZb06lYyNmBa2NdpVOJUvtR3DwLVxWPQzI5pi75y3
Ykl3XygBSIuTtl2b0KVzVVj76op+U1v+vVfxbBE/gyhb4dUeYLSJJV3tMlwj0UyP09JvARb2/1Nq
YwWv5u0SChPzf7oI5+KOO/jKd+uVGRV4pa+KNde7RqFCKh6PGeVVoDdihytjf15csTnclAy4+9gl
3P5IbgL37IsJShtFvc9bV4cWjd+zPix2aS4yNE8pbqjkpMGvGaxjq2EZfRwyQ8hTTmCdZSuF5fy9
FYvXEOaGwM26SqyW7mkvCSUEU9ZFI1Ty7Tm7nrA6K8SYlyEltxdytZLdibxE8sJpyOsDy66bXlav
l2KcUIkE9SU5Z8KjUIs0L55LZG+3FDJJaofXdq+thyb+qwDctMcNjQNTRLqf9nyrUO8OCxmGBcmH
95ul8dC/cquZBrlooveFtqCLaFCZ+H/s5ULsH2f74vmkJze1m1dtppi6zkVosroz09zMwfBUlMLu
aCyBwh0Eh8PCNYckewxjSFW+sNsrn/MbhQP0/HCXw2N68vpkPIv0QGhtVX83k036F0Puj+R3eP8A
kf1LMoPwOVHcP2Cm+9L4U4gpPZL+mYKhj7jVqE7X1Rp1B8bjFAvIizwRlWduA2s70LcYJO4bBGWf
7rnP+ph44ZBqgE3NXp1ffohrs271Tz5aLa9EQbbQYQ0KRQ2XVfwGbUDr2/cnVQ773QsH4WoGzMHa
Oh9mQlg6pjZK+09Yf25yXAGXi5Pfun60M5xzVxJJ6L/fQXQNZqPTtMpX1uk+5fGQDwqlf3afuPyP
QIqCIOfEnu0uaKJriAfMvh+WIEuEn05NB7G1EuKuwsnD/qALN6R5VY4BgSCgDZhl7xJDk8p61YGC
E00RD1bFWLXyEatqnugtXc0SGEwwI+v3ekSMyZyjJKX6bRaXypQSFdoFnzg2QvyBqj4/6iCtRKnC
hC7eqivUsI+rJI2+0ebk7ZYyCozxjcO7pzzjDuhdQS+Et39iShLbihVpm8GMuzH6iczDCt7/WBYT
opY9RoFp4Biux9etSoi1Or2dXf/HRF30aG8y0fXVPc98vGN6KaSWcYB8ir5Fjn3ljBsx+bL0HAGn
dDxdLC3kzLhsLzl/19bpdxqtfrxCrp/72awlMdZRKjRLtmrVROxRYfU1UvrOvV4MPwcXHNWQRoqM
uEV2JJF8FLQcrsPVcW3fTRNk3VCJK9YwyR9/OZNmfgxFnpASuxAik9XofUtUEmcYq9QN01uNVS81
lO50UrsviJdXFc+xb4Wzcx89UkWW7r71VmIOAk7J1BJBJAzTlPDOIOkQfli67+rIWoMoRxAoRC9l
SW9B7qb9xU+u8+soveklRNt1rojMkBv7xdNdOcvPPZ7M2BwPdsbhJsxy+2fHPNZZ7fNqvS1xXiyM
tr/kCNCY6P87g9UkmYiSVCpKhtdH0wA+vAJ22MwjWR39y8qDNc4bDwpXwh8OO0ppOMszArkQYNPX
yMz3mDDiMKkUL0mkh79tpdWI+K4d9lo2ATo6OmJQitdDPN3y1WgsW/ckB9zCQl5L55xbS4ezbgfu
VMt4/ghOo+Qb0MFKfSkcITI6I380WGQk6bAdv95eG/6Do47ugP7bnVyxk0VAnfFxqzJcC/5nZl7U
QIDm8HeWco3ielCNZ/VmTPUtIjfoUQ45TQcZNssaOV4FCZD7ZCg8ZUIlTJWGEqH0wwuJRtujqXJv
87ZScPngGzeJDAmr8idFJ3+ss5e4g7pmU39aOehp5CSDemUXwCH+VwO9MRTVZqJU+o+7zVCOCs6l
sd+kIHnzfZHuQzIHRAX7pru+KKwazBO2impL8Vz7bAD1rQMUehnmqnEznyDsFTvXlSqzqrFQiMYZ
P3ORBurmKdeWaIA7OFHlmaxFWwvANOW4PLH28ksQtSRSBqupuI2Dai0vEfCkvNuBJLWJVQ+VYCTb
BWdTrpgQtuV9qtKSueRS/d2udKG3Mju/9JKLDIMgv4ksKb4D/fqlAg+mixL1/+wkrpipKCShB8mV
jsz2txf6tf12w4/cZHvft0XfukhwHenw21btzra6WforqHXuGEgLrY0G2yI/LijpB80tL0ieHeV3
ARws0hZRODPGCbltz6bBJ0YV2GQck1AR8tM86CkAxnIYoHt9tyT2prG7jtbac+5EQZWOL7/1AfKf
XyIUeJjGvxBh63TJxoA/zng/gHlmasWkei8R9nooG5KeRsnRxfdmEAqrIRb49RBF1BkVR5CHh75R
55KGwqNHZHZIVoUrPwEhh9Q4jz78xKSY7zAGuNp9I/CZ1KqVtMfeThIFhlOeZIrrERy6NRQSiCGx
iRoWuMDXs9UmwIZucnO+BJzyqqvMAy9IP138/1zybTKf4qSmFhc+i9OdPP2z5dbsl4TpyAFyUk0i
R/gSK+Z10kdulWC6V6LTXI+CpYfH/hGa4zqWr1xZoRFL5zQCVm3pOn4/BEbmIgfZ8xuRb0CvztGC
mbfnd24FUJ32ezF2BRjYG4XRa9LJ8mbScGCej9fwxK3IvC1pu+hfyaklYsaEZKvwsYwO+ttK6Ecp
XBq50lh5KFXxOcuewx5VhsNNf/BJcEsqGzgZyWTN9ngJ2wSW0s5WlsXhM7Ggb5cS8cuS6qHVefhd
syZUNTwYKyHrYEkmR13pFrztR3c4zIIktpBO5heqGgu6FH6oTh/7PjD+qPWc8bSd5FSGdxqpasos
OOzTTbHj8JPWRJOcEA5rim5BkhzbeOWlI3Wi6X3Nx4zBPLpvaIfpAI8FfgQVJRGQFz2fxo9V87dh
Um/ekLTFf95B3I7Fb+GxkynPOmbT5fZfotWjOa1T01vAoczyLzDeUrYxgF9v00wunPwdnsUIWZ30
uKn6OBo7o7vwmJ3usVqfyyAQB2CkXPyxffh458ukhYNbShXzUcmRZZ5C/uv/yRcVJyyjyZwGlqSs
Ypm2NRYC0HrgU9u53BOz86TeZurQ+ZRUinW0sqCouR9XOWDDBWwoqUwOdPKcTT6cWUK6F8ibQa8Q
kRldzh1rWxCZGZ4JZ6ezjz8W8eGXdcLv5mN/Eo4pui/HKw/KN/edlWNlKxCjnbPJxf19NEg6gt+y
vh7a3GIZaS0LA7jg2Embao9TNu+bOGaeE6kEN+upwrwUviYVjsdvNFIgYaOJLxeJs9VkYk4IF4pG
Q009FAhkk0sxUXmNX7aT1AAy1kjXqQ4nM8Y9du+3uF6c/0FoaTB9gp5EgRbR/+3d3/EeE7JDKNbj
FfXQdgt7SPaA74jgOcpoVhgDerZyxEEdOW/SIwpu2GazmOGjcOEss+BVL+ssiaALr5Tibj7rP0Us
mv954F7dHOb+Ew4MtJTb5F5Xe7BtBvxWDGsl5ZB0hTGzj+8cd8TmYdzngJUx/dw2vA/oceCXEE8o
aYYlyNaboIlauO5QjAhfLz6XcnBrxkqLEyAs0++gK/uMnbWPvz085fd4Fq6nQdyjIW+/81BNqJTJ
f3L/5boPo5mYw5qr1q3YnOemUwgJ/lLta4voCv7aC4cRJiphw4u5zjffkxbAQ4sb36MQI4cz/WGC
8l9rnOCdOSGCBVh44Ku/qjxzDTmcL/2EFe06TV+CmvNPKQle3Ce6MBJ/g861uqzk3/cDCMEPHXkv
3l5mwnsfpIYn/tcIT7FkKInCJ3kbSMINCo2avZB6P/yR0AzExNhFerbh3DTbBEbVBgMOxanc752m
2ZX51DXT0QEeGDACpV878LdBVYaAocLsQSPs5uxiFdiXawxwQOS6smBjmGq/P3NXpXjyKGZHqIah
zhAUZcpja7x/Pcf9je1v6UmkWr6wUerVYFCnFrmy4o0nqsswWa2XPcAMgUNRE5mAaTcH6V5RGOub
mQ4LWXLY8UPNpTvGi7LIb0XiaYwFjZ2ZRcz8PxZEKiPjeblEyH2RPrkpOf65IMmSyd+XUr3yv1Pc
w9DtQQv6sTTkbQPxFXar1sKqyBzWzcaQi67aXv4dX+RnNPIAe/JOrH3bFXHqzrMZ0G3OFCxc6/NX
Dj+SB4wk/4qHyjtbK7j24APDOVDr7fwN/d7LOJupixs5FglOD9bBAjAkMXH/MjssP4M8w4PBVL8V
IkpDbn9RNgjitizVhiLHb5ub/lu4BtlHZ6T2YWCwat9JgaVMfbOJ7sMBRT4/qLyMtkzjKEAoPC7r
jWN1w5i4vfVL55VhPs1r+GDpyaQ/t3BG1O/bPZhyQ4RtQCPgZsgyVnlos2iDf2xRH152Z9FpFIBr
pqDNJm//HWRX6zThO4z3F+ywc9ZYREtMWs0pzkZncTEPIRaI3wHLvNQabghoMu6Eb+yFtUT/xTJy
xhPXQcLWsY9lgK5hncMVD52dunJoXRhLRY/aEgX5ergF0/u5SiVulGI5nXglOe9OMDKaHuNQ06/y
hnDu0s1N0MyF4oLP0vUV5rskoc5UjiNRIYUvaYSr3Z6QEuqFgU0pC2LaQspOGSTybBVCswKgTh9K
oqEAasgDnTmpsPRgjytTimOg1ekUgSHuI71k9JBQy9Sms7AP5u6ck4kmzNZ7vuJxYlPwb0c7ZSF8
+XwnSaDkzG7i4w8z8nzk/64NLvxIVCsJxILgTjxWMyCfWE48nZj9tjVAUAifzA5+Me/9x1c154td
DjWvWc+TLop/HdjNZxQ9ziQzdeaciFPhWndIyUJEEbO9YgsUwzuAnLqjq6E9Toexv0UuTFJO9O4q
6k4GBqwOtqZzjLy4SC94OgLMHRCKLm0iiEItqvPvedm0OcYwdLpR8UhdNwPnoguwFtbMLoGgbQQq
rs3aXtgtyvmGYyKoQNb/x5EVnc9vYnorL+JfQFhR0crQJEaP+ceMItXGInLv6LMMmaxXPd09NjY9
R49geiepUvn34/FLX90zqS50SI57VJ4/ZvIe4YP/2ciw9NZy15A9mrDaxIXp7tCOK97otONJSd/I
hX9rxOBLsxjFsnTeLDWOEhp0EhRIKHnTexEQQV8wAhiHt6ycaszu8ThiTM2I3g5DoOZsTjL2+aTf
0wzNx2zV5847I4xiJg2tJ6AROpvKa3SpdvGFryLeDIyf7rmRLG1bBFnqYVY80JYPd/rpkfmMbGLB
/Sdpy9B9z1zvsKKx17zW++ABrxvt4lqOBwUqXGtCM8qFqVyw7PJx1paYWKvxm1vpkIpCc6W402nF
JmJLJF93kblmRMEVgVcELIlhPbayyStYa/3XhnbL8rybzv9H9wjkdRJhxVMPQyFJFdddmq/AOFvL
X36jVhKvfqTZle72KqjEiTEhkyAzf+o55za+ZvgMHbQC4PUBV6aiyHZZExpYDkObumqzxyFWQbJf
+n1yW+MdJzdnciN5gw4Amq3TDOE9+9M8QJH8R+UNOOdiR91ivDmg7am5KJUnoInxyoEbhHz5Fzsa
kAX16wqexH5UIddH25wD/m9WNU9shYZKOd5J3R0PVa110D6gOdNQuKxa7uI4kY92kN1DVhfkzeH6
9neIqyznowc7bck2KdWHZMemWWST0zWPXq7FFe5f8J0um9jwhYCvX7VDX6jwV19gnWrwi5J6lnlV
+Fl+itHYKDG5d7TR7d9fdoOMtpeTCyLsrAihzmnsChSm9y02T8MAHlMxTWYRyZ5Pg2bStgWtpY/I
eDQE8NNXXH76UpHgdacANcr7vA+oceM0AqFuDVOPziJRujigpuHNMl4EEl+q89PMmc8/+j3nW0Ey
qJMNLJJEL0BLkftFhMS0ZGoJcbK2gJsA3nFeUMrQ5EX46vG5eoNUPWD8NUCIlSqygQEmscc5pfNr
emIVAjqlfXwRDDz0oKH2rRGIRDjFLtEiDXqDmg6gfLz+VV2ugdqWAhmXm7zxX4thI4LSj91jYk8e
Dab0OhBUFDVhySILOSagg9brXkv4sXuWZWsp4PdmKiDQgF1sujTJHgt+DQz0LOaZ6RRTywN9WLml
JyLo3y9pnlfPacuLnvMHpWimMl+oCYx8BPCy8TxVaaHkCjqngU9kEm6tptr3mwYkEHVlNw2T5Hq0
2/45XTpxC2agq7l6za83os/kXhio62+neSJjbegIHXD1SVxRLC1/8bBZ9rTi68n+hc2BciP8Bw4A
IEIiPI1yESBxDKAnBiVI4LEXhdRN6sGFZL7BlXmQvWw3a0orlQLQaeZzRQJNFTv8eYBZjr+aU8IE
TSZKmSNcvzY7M6Qx9oHEyCOmlnGwLkYmg1Jf8wd1jYuy4aKwE8uENwH02ukZWZZKR/AuWhsfpugl
Ip2lal7elOcPa9V6UAg+MBb+w5FHP1fFvMblhvLrtEKNwqLHXuiibhjQlJYOa/RKl7twzknNOlY1
gjFbR9rkaoRjlYX5wWxIHc7PLy3Mljm7F0BviVztMBSsEmZSRoSMvsqPrMMzQZJQHyJiiEBeu0IN
JldwsweJ+P0TUX3lVKvkEjrHKhqLmJCw08FDoS505Odhu+1a9XTiE9fl97flm2PLMRQbof2Mc36a
RIYwdyDI/D3DOpVsVPALmIyofzB0cq8kSodZouiJ9+GQzQ/25op45zFYdxqJwaB8SgHEvhpFiXJT
clgXIlvtShGI6sO+JMOPb/eNgvc0JpiYnkwYUzZ0HIWTJdMvG7SI7Osl28Lqsw/1wldsER4jn37Q
qiRPXiaf5xiUKh9g1DjY1G9NVEXGLYxf0cXKqvU9ogx2DcSB3VuLDbIsP0nc9ELPDeUiTkRBp+O1
65Ia66Bmc3bllBXy0B4KWMqLvVTpuDzJgy7WGenCfoVGGuNBo592ECa3ncsZD5sTMYAwkwwr/vMB
QAqhjMVENOGT4T0TB/y6rLNOLVY5luDPUBEQX4fg1pEwUdvOFbpMUvv4ZwOa8+C5A/FMdIMj8SiW
4tyttrHfTURWiVEEH+m7rmICC9viw2xHviMjuVRiTEhEr3mbroZLh5Yf7vSep6/5YmsDBVL1vhRk
R2bfoCFqR3FPP021pYuMQx5uG7LQNP+aVWQSVQwZ7qUNfQIDx2QFXzEeuHFJx7MCj8/Jk1LAwVg1
vPK3/csfi92v58tjhUVecmZqRyjawjezWyJ+Ia3C0QZdCFRFVtfkogZeKaWqnsfeaq8HBbTxT/u7
xg6Il6B5l6yqiahc4pdMZlWRuIlgaqJFxUpbZNgi47lWV+W2tZ/j66iPJJjmjZiC/dPdVJmcbf5d
QoBkSJZ9ryoSUPTJT5suSQOGDbeShwRQKSVl356iEW8sjdmlBRu7BPkAsoyDCWMbovkr6gXe1mHf
1aQv9qIco9REhfVNgH+5xuLmEI15ec+WodGKlZGyIs3yo89MNF6erHzHhMLlnRoXZGO4RxGi4b0k
vVPgPqC2aIyX10gxnEURSUOifS5HrrridPDe0BB0tHaSYE0ttrb6JmegoZZ8EKSv89gJAdu3mcR1
0iIDBfRzSSGxGRb0FBR2ul3hAPVxxv2IMH6MtKhvlaZJhDDNMC59P5tkgQnu3riF51/gWCn5Ueuk
QlifpKtK8vv9jt4QUlEKEijpauLCL5X8PQlDyCmpUPA+poLu9QFFL9JSQpc/7ZpidOfOVHTk/u35
IvJ7e0AFF2gwIo+HdXzjFllOAFfOB0jafv74ytJIynlNK4FjNxoXU83VxVWpgQNwxpc3oabDOhyX
2pQRw2+BWE0g+ky8UCjoR6ZjAQOLWJToK8qmnUsTAFW/PwCtLQWK3LFE0HPuQ2oyAvT56+2ibezK
J3A7XVHGehF+7HdPGPFSmAd50u/b7zZunjjp2yDeRX32laESTQfDURLS/JP9+BRliU2kEp0ImooM
4Jr9q3W2bZjpMrMWJ/X5WbZv5u63HhXnqhk3WRnPXQT0T2cEhkAoxMVNAwoY7PzGMuGKuQ829LXo
kwDD+MpGooqdcO50bhbJqE99nAY4Nng/U/aAVOZfuwETJwVy+jRGH76xMW4eveiWymS17o+x85SM
/XboAoawofP4Na5f+uv3+ERrXudMPhBK3vSi5uMqh1lG02wGscbeMGp6sqynfUnv5ugq6+JLAD5Z
OWM57B/UCV3S25O8in/H21QQGJJYRbUkKPGTE47cePbJlE9W92d+Zxc0DBOEtFPet4rKvbax6SSC
Zfiw17mQ65keF6BhLFK2ZINDjTk+yxNKIkeHLOx07ABuumgsycCLCL+9NqP/Ai+3w0FXw1lW4J0v
WeT+zVMHAGObiOqQ9+8ZQ+bI1nNWvgG9v9OobHY3WGfBqRj7dlvt6QYYQSAVn94++p/vxGZs98EA
IGwjEPovDxOuTaBmTAsCQkeSwzXRO/RNbwGlteVo3mRFwPIyofoLCdhJ/hgsdw3HD5N3ylguLYBm
KKCLfPfZKr83G2eGb+Qao9VoJet10q8jUCJvpDiWVJAFGI0n2zzbTwU45xXIhC5i10w5RuHUbQbU
6qWOFmFJ/NH5JkTaRKE3Ac53ghp/fU3ZL0QEflO2XEkayVpEZ/6bcVdlZ2MdMiTn4iHWq67sbzpv
Jq+QqAy1K7go+o5OndxUYpKMwRPRyHAhqz0m43dY6uaeXADkfKz1CdFv4gpfKW7irr5rXAmxC/pe
+DfdAiYL5a1XAAO2Bg3OH1rQlDS+c9T2uH3zQYwMBkkN22VvKIHuEp5CHRxXyUyGh2NpzQD8HqOS
+x/TAZiX1IosrF0CtTDgVzgEdXMy9JE8sknwzjC8DQ3n78CdByp+WlfIT9dk7LoEVkn/y5xzYPiq
NWQaEI5GSdlKsmcFdtg6SFFhcL54CZ8Wri7a7F4kHBU9PS0lIdYOg7oir0+g3NHAmdScHTO2aLWV
pztwLTg/COH2oBzEOTgHaGdVFbkFeJxUeENmUfK8kyvPGtQkfDUKpUX41Da3HR3mUvP9ohAgq538
p/A2hcBl54etYHDPjwGpZFRIMcepPEc4Yh++Z71s5aNIGPvKylcDvRE8qfKN2crXrzu8DGMwAz9u
HzwLf9h1CblN/w0iGnwIykzCReHbz/ayTlDEYiQlRuSHjrt2xynZ4or3Ruj2Miwe7mOOjEEv0ChB
TBuuSy0/6fKwmJ9SezS5JuJalZ3F7bt7Q1tLm15stHdEEGrae7EXeXZlaJG5S1pv67SnfYu/3fjf
4i/9mZ0aEnEji2JNh01/PGchlGqlRZffPyXRS3+o1kJFlX+FPv/GRa+I9hYI9e2FjlPuQnHt11tk
a5YjbJnrWs4hz1jtsWUVZxaGGnjdPvxHgFK3G4vCn5LGFF3g1e/KKRW8iyFFk/4BGcBpkS6jdZy7
ntEkReSlN0OE9Xko/R/MGu9LndkxZLxAHvyxN4srhSZLnVvAIJXJq/J9ObgZ28qf4iMuX+YnE0XX
6WAC+N726qtkPdYy90H0UUHmFzYbPGesS7TpUa9pKI/exXg87LuN9RJyq+U76SC8pSQG5vqjByD+
NN0leDFA1/LoMP19EDP74A5fqV9xVGb6+/e2AFo62gg9QBeRpI6ytNJ/BynpFewTjQnvQKjNeaBb
r2aDevTd/2v0raWHdm6LIWWOmUFZc2nnGvvbMS/Y4A6Uetwylzz3BI5Kz8FbDMAOTpCOb5DVAgVh
VQ4Z8HuXSNPSQbPuet0hmOcJLz8gNsSghrE74LT+lg+B3vxkR6C5iOW8/bz8A+VNPD/aouUP96P3
CiFrESN3uvJpcQFcqZAQVzMk/EM9CgixLqAPVo1Ql4bIfVORl1GMFCV8JDeWCq2x6mWxDvcYD3/4
foZEwmiMf3fYoxY8A5QcXaIemoXLXB4LSQ09xACLgMlW2SX2j4xCUq9NZELGaG4zu963B0e/n7Og
wg0wg6NdS1YI9LWvrR7MC5Z7huo000JMqQpwrQoewo5qU24+1n8wLCLRQa/FdvRPcgv35lpHNB2w
jsH+Hq9N5QAYRseeLeGDq11rVm/4D37B7B9KzmJddpOTcxJdbUNKpsNN7SQy8a5TKD3//LtvKT4A
2z9BlCsOr9Yxb24e8kLMQzlKWHqOmB62fnZfllfV2fklbtALXs8/Y3cdvxWYWsI75jNnYxiPCPD2
RKjF4aaoXeCvzfeJSs23pIBtPUmOktWJCtR803VCdCL1Oe4vJJ8GmMNE/c4asplQEkgn0KckkapG
/lS+/ib7M9icYPSuhve4oiHBxJwtviMIULHeLXFHnKMESJZTdqR8tK0ltUSAnvUJmiWCKWPDsbcx
Ft2cDCW23EVpnDaM/ZWmIrQOF0nQFPrP68cjcRDLfsP2S8DW1P3lqRH2dItRu/H3qTYgderDOkvJ
Go1hkmgsQVNaZBuRdrPp680wdEfiawsUU7S+x9DzfIa4cLVBckdn+832UIPEOYZ/rjHTLpqjsLCL
S1yalPiXYTNw3akCIg0kVUnk9zGeZonWZx6t5JU3613y6f3FoGxc9Ihq3P3dmHLh2HhJbvmErQdm
FSuUCgxR8v0g9p23OJYtNHXPH+rNXaKvI+DHhLTLbh0h22d/vTD2nvdkNUEF8dDCYggq5SmKP8Tj
We62eaLQMDhViMg0UrD2cac3Fhk1o1eSiTwCSZbwmqHRCcUmYiCgHbajNI1gg2cmtgcOBSvxRS9u
b1qvfxEzm4CTfp3hkRv5RjWaErCfAR0+exfFkoKQ2PQnAFnSaH5Uy/fbL7hqRNaOsW4I/w+U1aLi
SIh0vD1SVG5QNWFel5lbl+zvOe/95/iMitznBa5ysphLf1QyoVCvAKfYVUR/zfx15WuxSDbm9Mza
znRgSixj7rrfNF/VG2Zh9dYHhR4TH9YFibNRHtYPRHGzt03TqPT7Rvuq1lLSEIw/BgI41b1/FHQS
0dgM73VLUxoqYxV94tS9BbQmJMhWbGr/KFv+ydDr6chTKFbTk0UYgQvEgZreb2LZGBiAmVBeANkY
ZUc3w7Y9CNceCt7QytY9KokYXq3KGpmjvVbWFLS0v1rhXZ/v+VItKGYTKfXV6DeNd+0ZLjuUOZQy
sKQ2tHrOcIJtDBXndi3IBX4lgHTKkQkeyDPmHhLnlwgdHA0ZutfG9Cey5SCHQaZZnj3R74HjBieG
osOoFK4k9bJArU0ES2ZbgoDGUwPWxXC+1o4wLtloHA4up4WkZGHA1J3tE8JFP6nXkQZK5pwc1bVL
9RFh1XaU86/yO+WwxGNkG0itWZEkdxCnVbr6jhNCKqUO5+1FOpau5aDd+q0VgvbJTb0/4hK8zXxM
ZijahXcbtQBditUuVSDB4NKls6VxlvN3kAaRvxrX0sg2osMsX1qNWhasjF9PxqamGkKnIgL89yAq
QqG5TFwuRQfC9wwIseo9iMyFXGNy7kkYFHFGV5ZlDsaJYWjTRG/BM8cEn6qLa26K6WQxb7eDpuGE
hC9ntMv8uj6XSQs8YiOZodIDblNTrszYxX2aT6hvURHhhRgYR/m8ZiTpnRieqqSgNkOC/Pdn0259
ye7TS+xTrikXT1PAjLnfdKrmmUAYguDrx+OGr4Bf0Ceao4EQTID8CfaIl79+FRIPZBriQgE3byfC
MEyrGxP3IYm8cdQ/A575fGGSGnVBgF5EGIxf1Ax4Rgvsslwav8APFRNcPFsIgldtQ/yQprL+x8kc
rBtAEMQOX8eU2Z93mzJ4gdIxSxnkmn9hOjtG0aErHv3ePS3txuLVJg4HUpkYzOS5sttu+oZtlJ+W
KfpR2yMdD71EOPwR1/ge5RJha1PKaiQ53PkZIpSZpTfLBtqjPMVvr0LlAl43AiuHlcGrdqfapABm
lJDP2Gw1F/0S0L/S3sICh2EBSXPAI0ql2DW1pvMa47zvRq3WmxyMR8MVEESzWN8GaPLqnCS2+D2Z
85R5qWVLsZpQDNFf45W4K+vJ9FMhfWJkOhplMDRiQEAWRhzrA3oJXSmmQlbxKn+gIwWhbAwQ33Xa
x/Cb0Zgg9VkuMZv1d9IFsUs+i85BgRGsUe7qejqXNugy7a2ZhCHSVrFbnMZDNNXoEpLZpwoQDHKW
ZIkjOaw6zLMQ4AUtpOS9P0JaL5byzdRJSm2U7vDSydVQDIF5Kyue7fanq6JaKc9yBPXPbewLqxvb
Of8tw7E0UgyhLfEZiHsu890Gtec0TLTIhgRrRCGxZk8TZrQanXOLn4RGBg17dBzyMgV5m//71iI9
OXrbjqzLYH0sgYeG9lTcbwLM4WG3dgvjxi41LzQkz7uObNQaJbHChsdKpzu9pFob2z3wWduCnFlJ
6f0RIulMbkFBPGk0+umOc0UegmZoEoQ6rgmffm7pqkpnrBUPAp/2450g9Qz2VBBBTly0S9TvBm0C
PBaMq00pRMIPLopUmWgRT8jGH7MY/ZCiIJKonpD8VNoveUNSySkq9SVSLshRhRG7FnsUEmql1qmh
Nbn0NLZvKx01Nkg5Xv85Nb5BZh2XyNEYDvIIoQYNdq2wrlKl+ccvnxOTsxDaE47rnz5234imnM5g
Orsj1MfyF5E9kRCqGufftQsA6f1ZNMi/gGh8gLwBLbBQPrC2dK30T3/9rNhSPQIMjEBEW8zVQh4X
DdFBAqsxfEvAmwJp7GBJ4n2RetCXDsmVoF3BXd6CTJ8p+SHyPVq7wS9Qy/t7Ylkz4EivD/Osdyj6
DUK6n2T5lBD4hKz7GymLM9fZ1Muaz6caiO7qty/1o0QjrxWT0ksmJ1+BPLF+gAiHZyK98YtqiOEM
7Lo6h1jxu5z5It7ctARitlsYzypL2pQ1bSyhuK0uj0K/8xsQunfO4z/ov+TitV1AQovG/gPwWu2T
uxnVGy/KU5/PJTCdVjM/BODVF/iydRdrlTzwg7SdOha8Vq7xngwDOogHMY4M+OqXtxZUsc30jatU
rN+3sLi83mGEIxAMKoFCN5+x3E01xdf1LRayf20/sCcEr7HWFLvEIryirw4A8+TZ4rmOQdAEMaVo
hbF2G0t12Q7LmZm6ywzUXaQv83VI7yQq7IWvscWIVPK+rnDV0dQyI1x025AFmhDib1dONbhkofy0
arxbTmCRia5uPVN/94oK9qExJ8V7atpCFhH8o7lf6XPFBYrEYR1leti5MXbJXMdyUnwW87Qty4jb
rHsAA5WTej2KIDWiNGqgetqJNXCGvnu6GXmp/cqVu66NYEbqnE8RERSBjZpkJNAc7dNlc/yUsV6b
6ODowPxPaHN/c+PKtMVZqr1wH2SUNZfsxwchOYjl+ZLuBZlzZy3KXAs3sa/j8zlSKXSgO/f1aB/7
58fGXLTWZv27LJBk7F+pSrIFAVAJ+j3HkxRNy2dSVgvbLpSLrF0yv+/yPjRI9ZfsIi4UkYsH+u0W
/bV4MtzNkzj6NaXCkAjV0HCXXIlD7+qwqVtUChzU4sPkzBGWzWz9+RNvaJ65HycGKfIY2EJXt7+v
UhjsbSr2HqnSdJHmeHy9Vgy9n1xaKFmKlYiW9zFkF4jYK8okqVOOQMIE24kW847F9vXtymV2ZhFY
c+84OyLbE9rhnKqC+ZaB9zgz8Crt6bRBIQ8BuKuZhbYqhBefVTcUYZWkrdGT1dznG4s4JhkefP2g
pNOV/9ZlwI3BI2OysyEMkabYau6V0jKi6W2fdxpr1TwZ99aNcltPG0JEDGhXQxBtZouiZLGLMXgH
sSrevS+HXR+HUS4ZBg74bUk7UUOlt6YAsHgm1CGKbhbkMgYMwKIYNHKTrrqPxxFH/x7GUI1Os0NV
yS5rOSSjuumVqzXF/f96yEStAU5MV1HBazRtEUPvj51HrhgIYzrnJTNV0HxA6PMAyGIECcFhi0qL
caKscHwtmTTXmlP6DhMEAxxZacJ6CtbPxO6jEZIiG7Unvi34CMx/Y2puMGakISnJiyNW4e7wUoQ3
V90G2d8jGkKDKS9OFjqEOFs8ChktPSgJ6kfePx8Aul+Y7AJ1m/FMnwM0gLq486nxtuF4MCLNVNFV
IUCrxeXYyvn7pWG1349ozhKFA1PxAnet67ZUwRD6b1fumIIPl9jY+qw5IWGl2wlo+quHT+9h3BVu
waF4Fn1y1EXvcz0HCa+t65z+aWivQtgOLpeZCx0wfHjGvVpO7e9/QzVVp/MRT6EyrLQ8ndQaawMe
GbkF6UC/V5mSix6o/JNDQbXcI9pbl8RhGrLymt6UqdphtbxGYGnTvNWvO/4Qk719UENBxCF8zjlx
dbXLxEjicERd8CbER09U2oN0DvQGUiXxUcfxts2vIx+YbCGNMgyxXbmokh6Its9xfX1AthYyBEPX
rhtFIeETJ+F1KDovvgTiriG6rcVoZyXpNtQYMpQEANe734jcn+Q9wFfPJSjOy4yBwiBp6KukdlpQ
/+6wUzLQIw4MzSlPtSEV6HTprwMgSIGHv1j1C3Dybjhs5E9vbWG5Y9SGBPnL4/udZojniqEDlHvo
rJ2jlIxI5iVlR/LKnEsp+StHzbCeHK+xeauag1ctjbByuaexQWfHWVGqmZ90TYpSgPVb/h7r/wX4
VyBxStxA+7O1YacKRvLVkdtoon2WNGQeQePeeDUsOOtkON7hmRSZ7Kx3xIiDZ3p0brZOfffqHEMN
BnDG4Q8YHmz5TTiYOSy4oi5iTHEKCG2XrGExSTsUv/IKPrbChV6ufys5F+vV0GQtmrVyuXaeow3x
VLQ5aGvTSAO35iTaCM1KdgsFGTnQ7jAvpvTQU3nhRCjmYx4yNBqLZVc7gnEsY2WVUz81Zn1/LCDN
Ea4+r4+A7InjK8GNMokaSNUztd1vqWMSG0SbbOPX0Ojj9j8NPMOOR85xw4KiMOz1DZfESoENbi1z
SF7qhez+IjSWEw4qXFH+Xu3gYV6PYieGsngfWf2WABZDEf/hPrVgUxygKaPeVhJyRoT+Cows1qDY
rx2qurGJdQSXRM90APbQM7jyOrsJbQYZoFn/61oUKYmNvFNB05O5izIaRIqF71iLN7Re8DaDR3QO
4pfCihdObpFzEO0rqnFjxD0VEibjWJbnsBCyEPUOvtu1zUDvACg6YomPkjRME+rguMg93yEx0Mh2
+mQckx2PoYDpbODzgF5TWu6vFfqtu0RPb/P3ujIo0d21aONmGaDtK6O2m9MFEo/74SIbebkLr+h/
JU60Di/UJylZ4eQ3DL1q2zXUeHsIs6YSR0H17uxSvn9WVNOcX3j+4YljENh2VYikaFVrbxp9GZqd
jQljk2te28Fs98ATz7xMCWAsWoTQGtetvP7GtrHkMoEEVA3V0KpOz+N77i0+Q6qRVydMMRzeto4k
ajgaMwcsTgv+nXZwj3aC9tldDcEeLf2cqYVpOtJJOxWngoCHQY9icEE8OX3H7OS2j6INUApA49pF
FCIIR3ZyXFDbFj0eC3TQpKKrrICEhOvOjzuV8nHsS2vKXeH85KdtUbi6nOKb35LpTW1IX/uCnzHs
G4ehkdQ2q34xM7uwM8KQvi+WgtmJ4QINz67mH2DReK3EMVA0GKaWtuLYZLGszM27Xsjrh/aN+FF7
4qfGULy4bOMKOAmCwk1FSp+LNoMvHS6sT5bTJo912a5Z3GEGcK+RX1VQnUG1LmU0YreGRJfxs9a+
lYAykNwI93TrUb5L7HuxmzyKf7MgqZqbHzqJ6iFOhJHK7zblyPS3HR6uXTmWAoQy6ANOp4hzeAK5
9gl3iDTtOqidbQyOLz1xV66OCYXX+GpMUu4GQvPJxrzfddJS9u493cG708BISYJpU51Mj97GoMRi
Qfm4WWHa+YNYHbhUtmPxKVkMcEE1xvOdzOLsnlq79yTKQn9JQMxrnR0osprp12I1B+Zk9/4EDksM
1rWx4BCnTAqwK6IJZApIeWia7fWPrCY2z0T/2ffXRzTcb6Gb+Ca9iTSmoaY64zkWHmedAJ5Kk+V3
UC4A3v8QoOh1YAZmFZfyHqxBZWZekJ8hdc9fS62pjHyxbDdbPOAQI8NkS9tru/hGrHCX4m0U9ZRR
Y8nwpSaZ2ABGWC79U21nigMLEyAwEoQfBhG2i8IU7JGyFNZifaPb4tECO3XvLzQcgmCj6zGLgRAX
GN5GUQZCvYgEiD3jX1HzcIkyeNiG2m3zDgnZdnty5ucqb3Eu0n3q08IEYLbwKA+Lja3yIYPjUqpY
x1UQWgqND7DD1Y/oOXKMARYqIZAqjGbPAivlq8Q0p/5qovyacDROjisks8vetzKx5mVgLw4uLkg7
HCGkdCFpmgfJxw3Iq4HMKq+yKcAs5ijLeSkBrz4MdrQZRrv4htofKWWUb2gfRTGpsJytikxtaLGs
XLd9qkzwq1vQ3wftvSVMhF3GnVRApJmv0ShEYJeWYQwCiJ+HDkFMcqpDjxD1YgBQWmrLr7xbwC3x
9dOKkEu8CZvh2SZJL/psFAINBe5LD78w6rqjyvwJpWjvwGysSogViO9iI99PG/8sFKYfNc5551FO
ac288+zYh+82UyqrZHR70jbSvbJpwfa6WM13UCfrERpmnWqNE7eP8btb3Ez59SOgGBpwu6k5KyVL
PzK01c88A7PStsCMSO3apOMUL15YL7I1ZHqCSqV91zLncWTmQ/YXS4d4NajndpxtmfJoWiofBj5m
XEUOcoIFFgM0L9LUeUkpDNlUczoCwyPBMnIui/VbRKDg85se1wwC89VjLCa+51pPg8YKZlYxMfMq
YUwaTLU+/nkxifcpYgsRyVLY0SFG7Q+ocXNjBhBBStTjTv4x1hlyQBRPkPUsEG7cvKEY67AUa6jY
F+4aUJ/472uo79bJEsFzC5TYx+/rd64JZBADBOkLHc28e0TnH52rnyCLs9XBy1rc2ftfVTBswPRO
qR0PT8BJ3/4yFEftbkzhxrjtjwGcRRjB1DuzFJT7VzOdQI3QpYA/nkeE8GNIiZJPIe7mPnQAwQe9
Uu6RYb6BkkKlhwQNDTN3c6gW2ifJXhxv0tNydyVdkbagOgdwf8vcKWDv/zuOx4pPAT5x4XpYiu33
2juiXt34exSNnLh06O1VnfP0FKzq3ROKzlIp7K/q0THCGyxFzd50LleCUgivVdkIbYBs8JzvVCJo
uFLD9mGZ1miZQ3y2a18v6SRtf0H2/6PpPnmf2sqeBz56aGQNfWM7AxtCVH9TSpJV1CF5gFlK5p7e
Lv2ia7gtGf5cPWbd6Tmz7wZAzOw9tuVlPQNZ5YyNV+gZO1s1uREHy3BCG1cCLriCyX0EX5NnQ+Bn
gKhOTIwDBF5Q7UK9oa8CzDbhIZoBZaH2EQr+8Bb+PNLFo6l5OsAZ/kFXSqMDptiLHbS6EKwBji4i
uWOojwfKDcjFF2VoSR87X4RH+kVdW0xu6MmgV2ooZGKVu6HjAAHCiY5Pt+LpX5B4aS2h4fnbg/tr
/yDptGh1tF4etipz+A4cW8oWPV6ESEWvGskrGM2WSmeaerseEfnQ+FVrKxRtObDsvWU7tMik3Hmw
rJhmu9aLSKOHDJOZnH+jnNZVyALQoPius4h8GEgeZ1DgYgopYkdsflYr/0DOI5sujTiVhl+fORG3
dobm8VYFH7Zcfx15PwoJt4keHqmICKPvl3oMLybuXRCTwVmmxM3eOVasSoIH8hD7+m+K6OVBRFbA
IFOUEX39y118Y1wPEPpEa8tqivC8hPdd2PegtJlE2FGIDNRqTw3R4fxOgGg65xm7JTYs11GnzJ29
jkKXGFCGtaVQjdTsCjnN7ysrhqk2Nw5jI+Lse8nzhelifKYBYTtAhlCZTX+IHpcJVOMFVvkCuui5
LUHE/nGq0RXDf0DXWzPOG+QLuYVeZ7jIB4ErQv8ghh2HjL0EHw3t1273JaEobsVN01h3PnTREVNw
OxcNG3+eOeaGBsp7ING+670WGIYfucUw8FgWfj8WZeud93deh2yRnhsapkSY9TIzxmOQkq/S106U
lC6f+pv2PdW2K3wl1+Xila6A3gER00oubpcZfdrKQAoSMhmC9CbEM5ytouLqs4M8DJLyfh6ggsue
MBPSZzGPMdEKLwsmumnu7apcA8snUmDeQa0tT/ng/Z95NFPH0O433EL2jy2DCgSF0Fur7s9rIcFF
HyaxIwJN4E/tyZevUn/mWpdfTNlDX0pUhxEL8KtolvgJi2jDZsCZ5YhHvrGaBd5DlVfd04ruf6C/
Bbp1v5Ufj1vPGWiE5vNBsKmFz/IFExrf5OjHJlncVqUsNqglUMOkEmMelu1L5JgUZGg16cDf48nT
yj1Hrpv0l3uORnjWiSV5J1VxLDpbZxcjA3UPvMwq8pmPFlvoeErBs2KTENtUThwCbHYExSICmu+p
pR8/1JeqBtIq9hqM6MCPz1JZ7Aw2h0Su8uij50hxVaj9SynXpEIasjNg5sjURjvO2QT7aiYtTEXK
6zj1cNwxYSB1S7QHzdyO3cUZ7IocA5F5wIT1Kbo8T7M7cQC2sV662HqKJYq1hhrZ7ZLYU/vloAOr
ku/KQ4nUR3h5agCpGTrsyXkTkGAImg7TLLWIJ5EUHcRGFrq5ICveqQ5oWUHc6O9CNaXtTme0flIs
bQUDcwam1CqwsczjG5qA3URR2aeVG1pfU0zEdtjAzbuA62E6WoLAX0V9hat2kyVjKrlAP21+sm+D
HRTsgsCqDxREi6FT5m4EWj3gkU2SKmtEdGIsCJ2yVr0/jpWoBsl2prZf/lpZe5bQAv9JLwJsymtL
jL1d+ITBH5dTk2FR892aAyflfietO0Y0+SxZgHG9HT2+fuMxPcb4VRylsPIYuMaPTG7d5Kdtm89n
3plTmyjm6Nj7WPR3djaL0JEDatYT6c3Yrjdx67tm+s6vmfcIfQT1cxQp42flCNCbGYpixF18f9hb
jO3y2i7dRzuBDWg48x8xya1DGOc+dUVkIhOspIFCZWpGhSDoeOKyBSRIiC9aqQGwDsmW2viIskJG
hA/RnHwSj4KD4y7leS8HXyj36M8Bi6nB+sXTcIAJ46ePn7NVa3+gx1YYzrvwtY/Ehfbo+eRnqsvj
K3CJrGcTQhvbWqYegFbPq+Gai5Hmuc113zB2JPurgTdoyMUnQ3i/sJkUvle+srNNm3HxapoesPFW
Lecj72ecI3ZpvABFwNJTrC8DV559Xwzgf+8778D7UJ8cv3S8Bs0gAa3nvRuiJfQAzmE+oALDGrXm
XwGhYSY4J9rqqxC8nU1fb9dpAVmqHmTtHH7m6SnalBXW1j+FGbBqRHQVbOyQV5hsVkRTkEY2xMr9
h390Dphb2E2OZIUPRe8qQXb83CRxbvsVUhsNbQKHQJr7HOtgLOYUIFHODTeRlE03Sy6UWK9yy0C+
j79Y23a/ayw8gsemb+h3NPZUTthl4XZdcsd8SU5F3MKRYvwq+o18xN7hPnokVXT64GPIreKG2zrk
LRi/b1zo7vgxUv985y20DV0jcSBzmCNQDRyEuE/+NOyLMol4rb6FumyrnuIQQuNEmkH3Adu1Sq38
uKpjpODtmKPbJYNKFInGb6Ir6A02Tq0Znone6SmCG8/Mj4N8e8BLngHq0IBOGzFO3R4BvXqgMBvG
iJdud0gP/Y7LPTpC7R3E/NUU59/WWcQnA5bP05TRiRioLOFtatT+A8o1h9wvMf94jPdf6hBb02KZ
dNhqgHDWPHA5Xsby0YNNr41Yyg6sJTOwLdnoWpOr8qLNvcGTWQXGM1g70ymr0Xb16DugBgxGSwRL
r1dqpngFE5ZeeaE+OZ0LTcqJpG0UfRQn2+mMIU0lRUlhtNooCwWGFMHylst2ntG3nmAE8K/uagAb
o4VQRD3p+PYq4jpcO/mIDe4QXUYvp51Yw6BDpcgR6xjkYFkBrB0u/7uTe5dB03jtzWHyfsEKA+lQ
Gl3gsIig52rJ4FYhXZXICRCrPXR1NfY29y8DH6uhY+RAalMS/0z9IU/YKx6GXnT3Cew3fBW6cqeb
K6K707RBgd/1/tR3gJbkxKQ5zUvLmhJv7/tmBay7rWtpkKbJCPSBiSjN4LTNOipx2z1QKHBOiyMv
y1l4URyN9w7Am2C/V6RtcQOmlI9NJxClu5ZbPup9ZnOZXOOU5C/1OwNIxfQPMl4VJr+61TNkq/z1
j9wg8fo6HEDIQhrnlAw4IosbMy3MPmwt9hr3uIm7qI2fYoCPoo7iLYIVrC9zKdnY8BtwBLW6ACRC
MOX6jxGxnBA47VbHN6yxCeFBa7hKBT28hMgUynxhbZpovSWw3Y472kRdf8mO+1v/XbSfjIKE+MqC
ZUDCTq8vzGfDv9X2kJ0w2lrHj26Q6jDvlwLI+IjHKzxR38IbsO9+ClPXpw6g59L1TK3cPOxomxt4
xpTeWT43ackIvmKgyp3ia197nX9A1M+oyKvg8cweox02QEvgGZWBNzvfFJln9KLQFGN4ulAiPYp0
K4+bSfq1DSJbgjQitY5X4TU0j9eCZ1Ix7T65aubA2eMqpKWoRfQya2uxxz28/D4vfView3XIB4Xi
+qWGFFXms/1672LSELkbY7RV7cUOSIKXtaFNwjK8rmHq7dygoR65M2ziiTFFLJzozql9ol9aVrmt
f53muY38eiWjiFWVh8cLuP1Fk5gUM2aNjzdh7C5rE51aHt2Ykqkxr5of7nusiTNN1qRGcn0Ci53R
nF4ntSoQ++mHirPrCHcmL4fJiKUjYBN+jUSxMiGGMGWnJI70rFxjhce18OGUUTUsZrxT9KE6x8xQ
pjCd/i8YsmXPswPcGpKdTg+v4BhjgzKU28WmtH+Y5Bnw+bZA3pChN8mT6C7ajq94koqb446bq814
2DB5aY60o7MurcI3IBUFD5fZq7PktEXz1xZrh5YQg0f+Rb9FsfvSN7ni2L4i7h8SDKG1qowIjcgR
+HbuHszZKcK08Ji4EP3ugXNnW3F8aHMKg/Lz47B2+r1Ke9Vb8sruEbtTSZO1Ljkl+Sxa9zk+f7WU
0naiMOR6VY+6tnjBKBME6FToI9bOW/IaKBZ97pJwI7eqcOQZ7BW10unjLQHyC89WKKybJvbtN2U+
Qwt5ckeYbpEwBQIUkbOTZ84He0dHrbMj4/F3zKCJZBIqYSgqESvr5qjTgkvizeYcCpdUAKJ/Xdtn
LO19qqMoOr6mhrLsFksXBg9KobAcBTUZDuS7Kme+5+sryPLXRL7QpIiybNlIjJQ1MShFNnNSr8Uq
3N/ysJUfLwbQPaIifmiMBEpNMsRA8qpWo1O8d/dLFsenTPAyVHVkHE6mbqcI99EhFWQ1FvoctncL
mG0Ao4WoE7FX5UaRKFh5odQuXSy05yGc5Lu6vxoU3DEsCCanfDGLexbTXM3e2Lu9u+1UmrHCH51m
gbqXYOe9YhPmZgkeR9Wz6/p2fEdDJ7NiwmLQgFMlKuZchyzLGC6cHjrLT9oeEZkTYxRlYSDTvhm4
eL1/2DuqaAheVy8psIV/YFDlpjIDTVHyTFcMsmaGOhGJE0v4B31n8LqsV+eTB/C3E2RuyflxXT/C
2VU5pgOAvr33CIkPisvhPeCgjvcgLNC51I9JRVUMR+10uneLPUf5VC8TCt8yAuiYa67RMx/UBXmK
g+5QkA+oRS8OrPaslkX/MbEj2KOQBjaV2rQ0iMJ+xsYsIPzVnZAtJ2GJT2uZ7/a/dMO+5Qe2C1pZ
k3L1e6+tfuAZqU/5PijOh/PjyULYJGEyB66WF6nGz37YC/TUF+K/Trqqm4bJedCXhb7nTq6qPo6I
+SdevaHUun7cPuGJREsG+da1zMltXtaDCwtMcv+2IAL4DcQcF93t2H7GLbPCjnVVgNp0O/cw5gV7
HZj8Byt5XqDYGqZEgLmgfYYzFxJ2Klym5JB3NDdfbgtyULdeFVbN6iWUnBcMCtmWjCkDGrukHzkm
ulbBz61mmMPk3mC0wg5AP/rs0w66clNk1XuCQmcP3OuU+0bEJooREibYnGIJIwamm5Nk/lDBUkwo
vFozzwetU+w++hLozsGvlAs5se3mhIRIOPYZkA38msPfz36eEzmvE4QTOAW7q+s3d/KeX5T6imvL
ey6UPwhJ6pm9buIn9IpG+z8O0e3imtdhevHQmxyXdCxmrDqVi6xbGmkD6d+ZAeYISndCaEj8ieEq
5xKOVQHFzYRnt8MyChn6IklFwGMZfj0LmCnj4JDK0nI6FSly3CzE0sXvxWTTpv8W4FWNiHN/98sf
09kPxselgZSblwFBdGGjBj6hO+h8WvVVBG6qC9Rhgcn+HbToQ5J3lSMi8xTIoaEvI5am9FDv3Pux
i3ocodOWmMC+4PH2XS1zkzPUvDobZRJVgP3daA6nUNF/yVS4znUKIVi35jUU4SxdozYHZ+q7Q2K6
2FP+8OxcTTQb/YX/5goCidwLBZa44mqC2sWevDtpMvp+PZ5Yy6OGTYiyOMbon74XZrYzzL4lruXB
8yWhBbDR0t28bW8fZqGxALdHUL2PcoQH0ousQhdtQ8LrFvzU81f15Tv/J27tfTou1/uuoxxtdkco
KJLOtFhq7miIhYlNhvTj+HMbbeDX8p/1lRs1/h2QMdM3/1Kg1A1b2DFh0Eg/+RNK8Ioybz2BsE3V
a2ghZlbgeWzKDOXVYdVSV4mhgQ8w56w8v8rKk6sAVb7u7aDDJzc2sSwFeXL/lh9LO5Jt9isG+wdl
v+tgKyxBLRAkO/9oMKboGvdaLn+M6JKN7BW/4bvy+H+AJ3qUwbi0mHRmpW0WishbjoqRbmWeRnKc
mtx8uiOgm72ocJzH/v2D4C6/F4hZ6u2TAYUCR9LcSy9xKFhPILW+Av8yXNBF5ugu/8cvyNM5gOtJ
PyWoeekqaTM5gKVOt7pMaCV6zetFqxDPjfdHVI3dD4b4rl1Vpizn3nlsl4o14Fu3wVOTvKbArmHj
3KMQjG/fEopTLH/ne8ton6Tn2YVNetijUh4VDh8o+q6CKfVbXx+o+69bEaqrDCte7bpA3gpk+sDX
Acop5gKmjUOuoAhwNlUM9Hb+teJ+jAb+FP4DBYptBaj++/32+dP/SFShEmkLi2Hvz/KXoTzwJbq3
3FTsGrV1wT2jFTh0uhxAhKpwQvR/u5cX3bqTHwqjanAAbsrV7wbyDk/Pl4u1P739pde8vFp03rlT
eHWN+kdQxOpsa9rnAgGRn4ht6M96+asn8IHhrR+l8j0zW0W7MF+KrJKzkAnZQrWlcIOOpJ4zNK9O
7lmQh7qdTH+2Qnoz4Rh5FdBX/wufwu4E2ourJMKpx10WX5GyqgzHHXScFycF96iBRq5dAp2bAbcP
/ut9QKZ977fFq9YaAdjercW4utkkgBv3MBVGfV7P8boKxmEfzeYWRqilcW64dqYiEVu/JKnbjLGa
Tlm2pEk+Qy3mB047MUGjPkAS1AHlx+0/m3ZfkHbFnOS62O/Ws3atqzKg9RSjcR8hD9SHpLlwE6RP
CP+N+bTbHYdYsFa/EDZlC1fV3qzlJhUZA0qfA2sJ+br9uLj88PZ4nMKb05eSyxQPBWQpYwTnHLGx
cjmMJJG4N0tSTM5B5cAq31LRaW6D/bgeZCn3gFdF44L3sxQPFK9j/YVRYToLtnWtf4TOo6Jhs2jU
6kW3Wtaw3axOKBx9G2xAx2sPtBhAJdn/5Gd47wFSlayNbfbOAEcw53YmudXnAfOSOy/k+Vwyf3MN
gaQkIf/LmAEDqOePNE9MOIrj+SiElJm6k2DBSXYyQzRIXvirFMtLjVX2uO5tfWsghdVQAxQaB+wJ
3NedvJTpte6QbWjglJdC9WKfuMUUCEt3aZSYpmgOsK5tBUelFwsEwy2qHbMbB3g6gfefDKn0QRr2
lf4R2nGX9ozBjqj9g9qffgJdHMaEWor8jIZb51KRXebOtMpnF83cCneQ5uopwDpreySmBz0e4ggi
NLtK4G40GM47P2rn0W+6em/lzWwBB6ZMh6tJAR0XZ0NRaiUDv8aj5bWoGgXXs3kMA5rLXW9J1GgL
2f/32HkZZo7mBYjQ/fYS+DFVREkTB0iQcT6c04yKnE7ICCPRVSnCzXLBefAR7OQHtMX/egIf8U5/
3iQdxisTmhuWPA1qWZp79yhjVHlJot9jyEiHQ6d2nBpmrklrqdmhBSAaaQeruByGjS5hiOlQPbbC
xG3jVYlNVUx27IvOImjuuu+hypWSsKwu7kjOlIJ1oZXhEogGzmZAUjzbCHvVcyfXI4Qojt8jfgU8
CsABbeaXZnLOzKmV7FQ8zTkOHAQ9SdY9lYecTL6ZtpsyDfiCYbWHrxwNTkPD/W+D1o2OCSYFC7M7
ioCM0QnwXtJpCmYqdY7bVEBnmVEiup/p2/E68bfOHDZcudsW7WsKzwOabvsDk03pUsrSTtnucnk5
YH5N0wdEJV4x3nMmsO0kaQS17zrrx5eBqRk9n6pILqExj0+5fcEaDftL53B5c4xostxuL8AatPBu
9D9Z7XfR8mnSMh7n8aAu61i7IXd4fggYh8FWm4eQIVUXhVgAQqMAbZBjPqlcdGVccGZ/YdZ5wuyp
b35OxN2jJDWCYOIQAhYGuL0sPAT1ffyS6MLvx38FTFXDhoSdlkymw7MeLkxF6F0tFb+kiMYNgixu
Zuzcd7kQ1od52KEFqeodlhwa/TqeVmCTJgOLVm4LWGzKJ+k5u+3uXpqJbzB6bvU3sXznZREPGZCR
ezxGmMHCFc2n3Ewfb2nKsQ3+k6OAqIi/KBFBSxXwQysAu7he/Pf3NtwxF9wVnwp9QNiSL6i+wJYl
W58eWktrZUC20YwEl5eJk41WNg61fMYyyZ1aJ5QLl/yUS5Jyz9GzVrNeqISAbogWVmvbmPbi8WyE
QJwthqa8b+SzOTW8cTLHx+5VhN65wGJOMyU7QUHOUDe91ww5gqpwkyYJKPimKR4AOiuKemgOg97F
Mi4syzfycLOkDmwPBZh2WHsfCxgsVPFRx4lNXasJt+GH1Tph6w3gA8uxT5xZ4q8c61UBE2KCWVtk
W9XrSIbPK/uRY/K3F/yHxdu3sDbVKEX1QGn8GHqv0mGbzKgu2Ust+i2hTxRcqt8iXTkrqUCUtL0M
tuEaEy/T9Yr85VxJxVYSkm57eTLKqiAE7BaTV1R8hc5cbGvlqFdQksje+rgZsmunjq7pUmNa2mb8
QckuwhUPiiAsRNUWtSVIbqESvtnMPWvtIL3+P3mSlV7RxBHq3SbyDsbkqaN8yTMFz2eMwFENU/cX
a3+hBK94mfROiVk2jTvPBw6wahMVtI8c9bhbCsKnzgMq3aarPTiOM+XpLVj14wpjO5NaUnYJ++l+
c/L0JZ+lCWezHHjQhTF+3+yJ/9nPgFonOmFkyJTkPoFQAtaAMMkup6Wsy9738xKrUhZAvNVKnO7r
T2CcHHP7uVgajzylZZ58pr3CHvx74+B6M5Sl4zX8jqm/1e2KH/xvWKFrDsYVzumo3gmp30gbpjqi
4W1dT05N9/6eawCDb/9/LWZj+5Nw77MPGpgk+LG9tML0FDNxIOLoyYnxNI5UOoMh7NLhgPlwmB3r
4Csgfh5iVoRzwGqjfdLFXMXNb/fJoGkpGS4Ly3EsWVH9SDWnIqb7CLOMyh+mT7uOXfALH2K5+/vf
D3+Ozd8TUhxciP1wnQ2BQokKQ87o6GfVy+bqB3v4Vj8yD56sl+0bqv45aoWb+cWM/r4zbG+XZx5h
HkhsxEZz7Svf20eMxpQUsORpCXjEOiRdIwuM0E/oa1YTZoRSTM02G08Y7k5416uGxx+7IA6Bz+j9
HNuluzU8r7pq/URf6p7nJJYv1vgMLjaT9s1ku6tOi7/VDUnGpJK2t1WWQym39uFX1dV15u5oLHPz
oAz96rRgSk9QEbDZdgEuHoJZkOf2rR/+PTSEO/Bc86tAJjTq0ksZViiwt7B6ViWy7F9JEX6ZGq9h
s/goTjUHvm1ZG2c/43Q6iGHXWlUQi81MmUlQyJnhY8+wCzeIEc+VACPj5yJ7ZJMvRG61Rywv+PMI
vx7nsdRDsZzx09o5eHDA7CnVcA9BLBl73aW/1IBr0JizMjwFColbYagVscRSrSK/MXeylSkzbw0K
p1URHJC5avbzOdEC49rEBgxzjzXzC5BhM0WUc9khg20Jcvkaiy3WgX99X/64XitfN5vonULz9wG3
KRiWY+AmcQ9K4sHZfFqNpQ5zx66VTGnKe+7gszpU3P0DNSq3CGVSPnchYneCXrYTLrLWfplvLyoy
nWIzng/XvhkC3SxRlscm0lS5uMEbgRakACodTP7pCjIhJoSHAkAdqZWBmGv4PYEdLOIK9WvzvvHX
0tp5PJvuWhTdtAUno9mfI/IwHYkao7AO8h70+yv4Xq65ZG0o9NszgatMBjQznpE2AOCMfnleK21y
KV8z5d49XBvMcZ3hig6BQluZmBQ3gd9Uov/qBLD6pYBHYzs+Csa4uu3nWbNfXZDxtMxPMy+IlCZX
Cuo/ZMuKa1GCZ6j9OILAyKEX3KNYoScOnu5rf5UWKb5lAOo1hJQjDcqykOX0pTdI+tc/uu+2ismS
69bjAvv8xzKgRi1/QUdIaZku9Ca/sXU++7NRWcZLgDg6eLAW3vNc8p9fe4xNU+WFg/wFvJbwYTNI
/QI3fFQoGSp4llk3AxTw9aj12YAx1nZ5yKOu91MJjcEgxh5mpLZs0xB8/1+2nsO3yG1t+bFjKKVC
sJRMzvd0ne5z+eNQoUpxi62RpoD40nMo6xuuiYncpSm6HWHp/R9x4YPvZF2VNTKDF2eZ3k4TO9Zd
5aB5iftM8HCYQzd3TFQCQt6QdSL5fIYWzUnaZN6gnVPWxVG0hXQUc13/saoJ1gsqwhRRrEPgNciv
XasHVPQCVi43em/+EaiEkv8Fyptq2EkcWjD06NjZFwWKHu0JZQhotVU8waOLmsImEgLERWiCYe76
P+XIS7Wkzrz7FGH/1O0am96NEYDEXllUL8xedhOBDb3JWJnF/W/4WyTfdMKuYnGTHmhox83Jtx47
aiYCd7OQmdX/eJmE2y9vaZtK7AVA6kRCYZPugCsp79xIC2gOYlmPBxSt67bLt7KwtVYGfBs65sIf
G2EULC71+vv08tFSpnqzPDoQJaKuQq27ydWOTMEDzm4XXT8mthp+kmFjeLQDNC4DOqgnevJrTlvR
nwxSG4THV8f04r+OhUYegg9LzT19xZohgPqJpuvMXUEMBcTfUb3ELXjEn0utZuGDVT7g87T7CCwq
iUsOyOgzI/KmusoMsKt3EV1+SjOddzfeHgQnPBn3VPSjYy9i8HbfTaP6zFZnRZV8o/6pU9kQzqV1
j1LuapK7G8aIutgYu22uC6boqrz+jHA3PP35NtsstPoQ+f8ef0cpbhxq5hQSmzkmAJeSz4OVCdIE
f2kPaB3/B2l7xQXPsasKLPeGCdg2fOB+8DNHwehOuLI5SlR68pYL4zbpZAVDyrgXgwrazgUq663v
/VjFejZnHEkuMcMJBcVHzpQfZ7qScnED12zJaP4Q4tg3jGwI7nieb5BgUNjVUsNJy85wLOVpSu+t
eHYGTVoCFxzdY7w7vArlHoMy5K6xOJ0rNKn1LWJhg5qfovhcjp1V3Jk/q9UjZUf9ipUqHcydKJxr
yu50Y8/cUkKGr6JRzNVWn1s0qSkOXVsPSdJh0/2P3hQCah0A1RnMcRT+uB7Q2lJPScNvKsenpV8I
ZXVmfp8iRmEZI3txDdNxqoTvmAGDu871lbLoixyAQrzTc+SisCf/YEUwwB0Dqf0Z64QLgwRD+U4B
YAmByal5cR04inWayudbZFvTuHqhYIEeoXwjehXHsU8MSK3f3q36BPjJchdLOlsKvbsQDeHlUcdJ
PmNCSe1M4lP5m8A6TcqVBFCvo3GARBZpxLJrxezO8anOjc/NgZUmZ0YpxLINPZQS+RPKWGfyf4GK
L7+wQZW7SHwnNqTnwpvq4SAxJgdJ1fxHCSzj9Rj3mLZv07ofczoybkYgRqg6AlmkhpA/q16dSbKq
5c/Yn08QuB60hzLy1KDYTTx1RLR6I0VBsKjc+PG2K1DgjOQQzkv9DctdxFIAkoo2BOKd5/llrf84
LBClTx31/zujX+jbniksNvwtmoozwK/j+tYO9tGAxbFpZ7O5UYcTDIagOq+n9KM1UbHHVs+7FuaE
TIW4i9K7A5pB4Xyr7xNwtjDlIntD0c54yS9fb1ZkuZ57FtgNmAMJzXrYUsAepGS6VTpvlsGNK6/x
IHr1pZclGMh0qhPNOVE80tSoYHPr4NVd6Qgi1iiZQ5plTtNbZtRNp1uVZtMhka0/2KN82uVFmNkb
0gHt+Bb3z9LqEMgDXUQB5hibLZfpJiW1rBXnyuCSkDXkVfLB7/Y9Rgt/RxWiZ3odrf9n35g3fWYz
PmbBLlqTBiehg19vTyLjj3snQAM9edDFOmJ848tUaSmPNxVDAqDE/3AG/CmDtBvB8keyB6vLLTEu
NBPfLmJb/Xm41XP2kHhpMPmWXod9aPbONGhDQwJQ9exjlVV++Oe6mV8IGprkjiJlyXhB6NIU9rVD
czB5ep/YbGzitg0urYRCwuB/ZXXU4xqCb4hgv1cqbutg+sUrk7o6nStc1IztOBnze+BpOiXJ4b5f
BFfxHPYE7sI8+kJa7dSS2gTE12QW7lvgg4e/jPHGqg95kn6/zS8HmIX4fMAEQ1HCu8FfoWVv4aSt
2oZ+7VP2xXL67vLGpooaIjRsPyACrzwi6HD3HyE0+J9UTiEfVj1mrYPs1viUtPgmOhcVwPYU/JpL
de4RoywwMkdtDCcaJE09uVCYPd7WL1GHpNbrjGhIjFeK9gmH3cmlkP5JGXQ9YgtExf/rwytb/pGz
4sFkADqigEvAh8rpWp0n8rpP2THxmqJBU03mASblW/QF+fhd5TX6DwHQh6L9EFutdi2whD+2XSyK
NljT9S+kKW2WdG3w9x2gkuf79eUKJRbOWkZYOzw5ay9BPPcAdBTmSYpwbd7EKh7ZKUsF+JSFw86o
jYmRTk6qqAI0/Bx4vuYwfknnDOQK+5qMwFKwA2jrGKIlvde8rHGdAJdwZCTv+RmuJrJUw1dA34/z
uFIKYWZbB5TCIlPYZiwzRWfPz1uIlCILpD2ZUj0xcmQOE/Svi+xfrDzwbcogOku4h+EMZoproIVI
V1CRupQTgvtEvhWm5fTytXd+Tn+Y6sfF65rq4eWcXp4tpUSEF1gmlojwUdS8mIpxmJUdrVPY1lIJ
mDlko8vbD+jXNo6spaqvbl/bfJ0sfyQXQIqBzQczK6haUaJgWwnK2RC7igVQR4flKin/7u6a0cjA
RyOlUohsUhzu5ScF+R7mJ0akId3T0EJ3XvWVPYOVlLnHLb6HTlA0WgUQqgbgYUitRbmI5V44Nadm
BzForGPGf/hiniIJLRPTzbKiqaXZi1gS9AX3uCUgv9xIz+ewdHTzAia2Qdecx5BoZEGCME9UHv87
eHIo9ewP8CUjOYmQEBZ7QBkE4kdp1OPbhgCRipHJyU7Fdq8sUdZtE9gq0GUM+80UkLW6jLXdXYq2
iSmIyQj/mL1Ll3CDsYvXtHcaz25PeN5JRo0goU5irwPN5mQ//qG5850zqzj4jwrBkuLsewM/TQl9
7/8mHuaMCyfBiYBE7PNRHov4p91GzrAEBJaDZShXKDUi1OUpqkP5ikdmp/OMebvhvoxbMO41KURc
vrwWFWCHZMuAhnoNdd63vryai3aBS+u9f52z2o8fl+WswaBkHHzkX6v1hJcCAmqXVcdKAOvcWQUP
MrXwAbNdNPde4ipMaPByRvGo75MNA/++2zMHXEmsxYMmcg3XdNUVSIEUrukDCvX/oSyn7678beMu
uhV4r91MZoR2NVjdjxqUqPb4V1B5OoXueN+wfIlgEmWXyKxJIvmp5CpsVqWPiExo2/runRJIog1g
YGMZ6RAQYTwowoC+zD5oYXCHlZ4UQlmJFEZZSdDCuDA1HzNgq3X7rzGnJAWewcEToGM00F3OMT7Y
lp4DKD+K5BJbHZzjZZQqcFeUzznecqCfB9hVjkX8sUBDYDAoKobN5z/KzsngvjuRrnYTWiSmYyap
wpCNkGMplHhg9Z5sM9hqDtM5ZEAZJ0xSk0VJwoBzL4GAeK8pI2LKEVbs79knRj6VXUjTIZdevk9V
ubthCKpKHCJyzwlSYYbzhw4/zcFE497/g2DniLk4l+7CwNzTGJ/e2V//E26WQUDo7MR2OEnxcF3u
nXy5ML6hSHJxamjkBz84fdhWHAUJ2oxhVrGa6inKPH/XYkY7ecVlZvHfDPGkUXMfXBAt/2Py2dfW
knhM9/cQhku72nacn2aQruOHsRxdX3WiGMf3Y9so5TZx3DfPseMc6JUkL66b1/Synrik0GVW5RjK
UQnnScsFRRhLB7o5yvNMavzzriLmuYvwY5R7ww01xtUHfvJ9NpCItvmceFNKkaAe9RHWjUMLjWe9
+zUmcrEMgFkP3G5UHZG6RYNI9eSha3+tB8iHZBsmYlah+fah7GTn/C1NOI76bBqo21h3iZM6ii82
BnOjVftGRbJDU7TUPq1xxE2DBUutMbq5WpvwxRLgmuZPOtDRXX7l7uh1ogQ4RkwBRzwGjqKrE67v
LHdoWaK40AT/rp6jVW0dtmW0MioFWG/iDI1/FSys6Wh+uzmseZH0hgRNSV+uhXWAF+DuHLCYhSSC
Ez0VP9Cgar5h91KQsU0X1OPOsBXMmByU47LQINYIgaBn51HtCeOHKY6yAI58fh1/3GzbxHAzbFSQ
Xd9VP9teF/bkI7jIHIrWY085DpSCyLPforoZWSq4FmN0gHkYqRlfq307q1UG0qAcUnc2J/6Yn/ou
alWdsaelx26XYjoKiS0R1RVMhAJ0z8P88vxkGCqu+iuuk1uTLgKenzzR6xP3S7T8NyO9F8bbuL70
uRvmnh2a25b7NKoQxxJG0hEVIYzGSPHrZvKkDrCKs8V8wqa0LNSsBzF0CMW4g6SuqGiR/wo7P5zY
Xc9r0bjcQmeSQsA7GYUOLmo0mM8sLhIlRDTPeHsLVI6AKkVi7Dk6YrSOcIv2trFA3+lD9xqP858p
WV7riPPOZGN2c/vT/hoGfJm4Gu/G+fLTnh5FhammEfwW9gUECmlannRHl0qiva4wARloZhdRASLv
gl2HBInQbOfuzS+Zgn6De+HTS1EYuMLXGkFP7QAIgAS0mBZZxAJ+65UZYUQFjYoGusYK+9GMlf++
DvtXkI5X6gynJH7Fw4Rmp3Lc4NH+EpigSz/t5zkaOX2Cbc7iWR6GtErTUHrEuTuf9VCw/m8671wN
snMUD2b9hTSmEoUsXIZxuBA4hbmh4eFfYQyPi4AFB6Zq/2pGx0nY/OY5w+CqvefwBfFkb/MY8laM
LpJuqEDT8TRAC9w6+XItCT0ZNS+KkAQx9eWkoyfP8ZkKV20EU8s5JOXAMdturR7kMNNoG2DlzrXM
HTAGX+QIMqMt8RA0nsvB620elZLAO1uL1TTA7oh8BPxIKfWT0BXVGArQD8BD4pGh5wny898Q4J++
tfR7xn6W303rJz8mCyVpAUl93fIJz3VbrSbMCIKX1APD3v1ToHd/eTVECOZjyEkAjqgHKWZbPx5O
7FEaRh8SEcMiHHONeH7yOjQK1Ob8Lc3LrMLf/qOND8hmOfpMLuDGSVPumoRr97utbgovXIugfiIY
ITwS+JadgipGusVRicTXRsLo6QO/tlthx5KAbA7SMUoWKhRu4DAkVzd9LvC7Ect1Rd4s20czfTAt
t/mvS6flihfj8rmgpi0CjW0x7X+JVle739GcKGeetWRtl2RmGR6GCSInPxbB/E14orHmZuGF9T1m
CI7ziSJOuyTUByYo67pyT0H9l/BiXyQjpK7Bf3JhzxkSP2JtQuX6EM7vxf4LUaIcUu/3fVq8tk3i
wSCqhh8rUTe/oKaZLntuj83QSGb15/VymVjlDL3sl9eodX8f+mxzkl5eyy1RU+xdW3+RKDDhnBfe
IhaspOweJ0d+6EKLmD6A5Wn+O5ZcRaERfkciA2lJd5hIcZPxXJBdwm9+oDDVmAL3Wlg3Kn71laxB
pCf2f8ucVW2lDM8tA11D6sNKH4SFP7LfCIQUMrXmVTo+wT1mM7h9or22JB1ua3shv2Wa5bmqvxJm
/L92qZLXKH/Ue9730IczQoCyntD5ZEC/e4LgC5SGqJVFldqjNLe8a8Sgb7Sr9+9WMmYwrtHbRJZH
guccfLTcJumIbSBWHtHuTMeswTTT5mXLjgcs5+BJcfcjx4IkFyYDK01HgyBuOJkxGUCe2mgeqQp4
0T8u3QQVv5WIYZmDJxjS+AtsjEHMqn95vXEZQLIe9EZgg2/Znh9IBL3Y/kUOJmo/gy9UersiXcEO
H9YqVoZqob9wSGvgajLOal9GN6yJ6uhuMONmDZLu8nnWKogoOKwb2bJPZPkuC5pppYZtTtSufr04
zXih86nv8HJoHwFmuTqt+xWi9Z6Y154NpGoZ7FhTCm1sMc3VuH89N+npCiud529EX6UW6iwLh5Re
g1yYpDqdwFxKKHsNY4f17JGQEWBaTVPT/i2PTKw9kEAFAUwnyXp55L5FzpQE9a6kcUgHn2csBOiI
/t9Sl2uAv0P+dsIYCcVloQx8UmC9Vj5Vg4b1yJyfMpgBHCIRuwjhb+J8MJgZT7CoxO2HFSoVJ+Cd
sRDb/E/KtwquF0xvVePUb25DGzuT7L8+e2H2HtsR6IqO7W+hCLLDwiTd2j+4k/uAIGxmQTxEQbTl
/+Cz5/f7rEYxjEGP6pcQxWvh3cIGZSlCydiF25n64m0Pz7lyckat6Agf6vZEqB2sInm6oR6wQrW9
TzC/XSf9ZeKBXvNNDeYWuqPE5sFbjsVhaD1Vff4+O7klmtchEtru2XMtw9Vnmlv5C89mjYXUr09u
YGB174qC7ml898nkXDSBMj1FElB/tdhU+/qqfvE+V9HCrFOFtZup9WvoQk5XL6cPQ2dZcJPJbvA3
GYpFK1db7lu2dMpRZkeU9owcbGtIxhQ6DacPxxVFAOJaICaiCaAlgu49QfKGuD0PDCkmkh/yNyGm
JkIwzl+YblSatP2PQGfwDlOM9N5PG2IZVzFBbl846+eHF83syAUq9RuVQ/DNBWY/YDZt6pyicgZS
89+EOTykMo2bcPyUsr1koEVEdv6E7/+fjqE0zV0ZahYJoJiJ8X4NPOqMiuwIV1WOX4woV1QeZLCP
y6Hze1vNBWtRDodOzh1d71dn/LRLXFTf7Q+0XEDW14d1SZ64EtTlH5XJGQh886ddXnrCclOADxkK
YFRIbobQNgSPp6z8yUyC9fQeolCKaYHmedisilRDZDPdM275IBCK9TyuKYbyDUU+hYIblRIVsUZM
74q0pcQOpQ9H3e09ddoUMbZ4IDFgGy0KD41TaUs4CzdvpIqreQW5ChBKssauV+kmLnJG51HzRLBG
ZTcNdk9BpsrU4UTT0YnspL3BERIg2u65N/BQU/VnQBddN6Igm6RaUJ9HXtx1VqbkBdCcKyBoL5NB
1uLOV9R41+esFdyClcTuFTkSFwa+xSjCOTIGsbEptW4KGlC6PlnGNzE2wbKLqPT8absPlE47kfst
yOMjQG8XJdX4h+hLg6GPJm8v4ksR9HZjg1PmIiEk6tRgM6Dy9RnHA2iDoiOrjB1pn9u6/LOXSMsX
eOC9niF6BMkY2JZt2ZnvqLh9s1n1sHkg1ZieWT01eUpWbHdu3FLN0pj+d9lBhsl9EULGJonO/Fnw
rI7IfGvkZCoaHg8NF5/BaMLhg3eV90fMZqjYmm5qbfxt0YhtFVnEqXmW1PO77535007OFJA04e6H
ppt/2ZGeyY65VlN0EX2pRelNQnZveO5BiopvoNLdF4/DpFxvLEBecGqQBjvP2DdSFxWEBkU2dZxX
clX7X5CagqNVk0xptIrQpgwMYC5o6wWuH1AUweIQsheBrxV9P69XQ378+Vw9QgCOL9roiS7kcmwI
L+YNxFmzbj95FlgyFxAoyV4nlP7XEowoTVVrKNJiS87yKu/yst3WKBghziPZeiuL8EiXJMIGKBpd
lp2bYc1WTSw/JEzhqigO96GhKlviwna2FVSBrRyKuW3NhE6aR/BHiBIKiv0/lwn93gBAcWdggYrM
zjHgCPtFEuw92e6lIlkNvkqFeRVHjuxO277YgBtJ3LCzxgsYFYiVJY8E3cXD+7gZQTRmg4C5wxms
pCbxRB3CJZfzaK3CP9+7h0W20ZDk0uJiX0ZjiHakxMffgmqf8SWaFxbXA9i8BPqW9bWvaqRCXlte
SwsjkSkNQTpL9FB+eyRhvmfB5IZk0cBB6StmRfFdCa6TcEbILemJYXKP5imQQOanpyv47+8+nj9Q
vzKxHrWuybQY41J9KQOsK63zz/hGGby+XNfqKGh/Aac9Zzp/iCG6FveeFj1spoe1ok+dzDXXgaGx
T4oM1EQ5bFcI20CKB3B99u76N/U0GD10TqJf9Z0RdD82I4VsXDJdmrARgRj7om1x3pCLUzaBuqNm
6aiuEhx/RSA+6ngg7LkKhZ2vMlJq6UIJJ/BwRYSKhvswmI8/k2Co/Gt7Q7QXu3UAmRNwphx/7o/o
Wkc2MwySIlHKC+tOcG43XDb4Xm9ZzlO5IehtykTY+TEmqgfqDBQ+xM2EDkPBbUrpmRp7UG1JVyvB
/oIEtHsMK7pLpNXckoj8CP/Lzqkakpcq2XikZD40CAIEZQgQPHpgJkkKMmuAOqdXmPKQsFjLhzgD
HFJmohjux6l7Sztyk+6fKnCI6fHCVazeCQhvdWWN+eOSYMFNFdEtTwbxjjcteJSKdGF3qh9ifMN0
QKj9eO8THfwqZKl8NH7+p795e+PnvZdLPU/qBM7+5JqmhWK//XDF71LUqRVBiTboHv2k87bthlwz
S0JMhGIqmjYuFycR++pyzNVZftHBSIvsR7Q1zJv7tNi6SMZ9aCLOe8Is7k6cS11c3rs3VOIlMiDV
MO0Y1FcASC6ZOMmSsFA6xflYUj8TkM4U5zphsGKXd/hh8ZFNl4r+6OzPHaF/lLeoII1rrcMnUUVW
LaGT815A8TgTTA7N72DfCvk8b0/zpgpcGsnPvVyhQDxMgG7AeS8D9OW+9rM5cQTEnoXZdVKJnDYP
CNRsh4rKjUla09+GDRw6ue8IkvOSNy+psoZI4loW3JC21YtxBbYPc2i3d9/lB6ME5P8pzpxuUq6q
IkBlvKFixBxSxG2SzWgDlXjbHeNOSl4QUOHVivqYnIO2klQy4bPA4nznt+kej0QxhFT7oPg6pafN
hvOZM72xTz8B5lhJtB/ZAScErSXFPer4msfWYe3KZd+Kq+ej+c6Bk2lz0lVx73YIiIQmMS1l4tnM
dd5pc+4fjeHcCm5hsDOt0yY/cdacZUQs+Rk8lhwVhrEcvm8xOtzGB5rLG61rV1PID4LuV05xxyJ8
V9ef7o6Hk2lgzgTY3BhrJdhPmHwSoDDURGGPPbLusp+CC5cwdEDK933vK0GYqeehcV9M5J/94txp
Rkkr/sahz64Ef5XLpyBXW1OlUZq/kpTPSHhex1GQqxVPf20P4U44O9Lt/GpKZ+m6UzuJnHfOtSxI
F2SG6/IOfSdeEZjmak0pXRpxMpfa3N7EMCWLrBViqCjKxGqBV9aLtNUL1c/MTdjyewjUUmUS1uIj
ILOfPSQnkFUTQT+zzDJAq66UvjlNh4GwmzCqdT4WPJ/0Ogm2BC/55lPIRK4NSKMprzdWH8oFtb+s
PVY1YawZVesMYk2gqaZEIyILMTljIljoCXyOl3gkmjQzAQsXdGQo58nmcaV5Nky/3WBcRZhgNbz9
bcTm6SAj9mu9vEi3KpXrF+md555NDm9gee8r1BenJAc3UsPVARrVg37VzJtH1QVxEKQ61/0oEtYD
cdZcCUf+IfWlJy/bDvu4k6t1pywvtWZl/cpsyZxzzOaVpA8ifHTkoEvIDuGpe3hDqh7nkj5ur+cY
QF4cJE1U06mpDTMRwA+YSGjOa6XDMgju6/7+zetV3qB6BvwrCpyIeIcrQkadeZj9rQm9e/T1tdtS
tV06PKU5UbDaMJBYSSChiNJBzsuYQUf7t+KWp8qibOF7LrysxjAwVlFdBYKvcnclspkW9ptxZZCZ
svx8V0Qhxq6ecZd2Xqefy1cinuNoNOOYrhUUYahKqouXTRn6/EKX2LgC/Rm+pOuDtKoF/dRufehL
YFSO9rPOThOpEEQMHPtG2PgLCfFU2FEYGfswQfBVh2r1fJBHwwEmJn2gIMl7VP8JuxoE39T+F1gR
L2xLkyfzN9fBpU0iLy4bKyrta+0+nda7d5gBX4i0abKaxi91oHvppPeEFWUscCIJz6mSU3TjUehH
OlH4XYktzKbU8e9nbPt3Py//uVOgXQZWFMaeuImyL8s1C+PIHmYj4+PNyf1sxN7nGJuse3YI0849
ujPR4QLOpN9sLZG6v98+c8VEY5qCe1gcqCRNZoyJJ6X/VlIf6HZd1t8lLsHd5Ymuc5QXjy5E3XKq
X9Muhg9VvPbkfIr4umqn/mV+22vwtZ1zXFvMEFtWI4tnD2ueYr3OHEl4J6wgG5YLsVIZTYVUxTxb
Rv3Zv9ke7uHng5jrbfUSq6m7Pysq7mKr9eJq0gC0zToKTWR4WQzGshoHOQhmaOuXtj5V8UgFuIBL
dOKwCsSNknJ1zzAoaXLgz9tckFj6bXXUTZjKI43mEnqezkOoPYeUrE1oBbi4R6Omi/1fEo8uCeYo
FvOqJvjolbnd01QM18eh4kDRWNvHOwgNoZ6114C4CRXx00rTDUFgjYq3rz1cDuey+h9RRNRKiW/Y
il/Sc0W5Cvm09ckj8bcKdE0Z+TLfZWcYCn0jHvob7U6eWd2qh3nM53pp4i3pBBI0bL4yMpLJBdkk
Vc/h4CI5E3RBBmyKJnvgWaGrKRSjltDiDFpaGQsStGEXA8aVaumn834qdYnk1+11Dz3xvWgf5W6z
lPGhUkj+f4YB/p83h7aBHPoXx9oBG4t8A7B/ifzrYFf2yIRLWBPRDOFuF237Xdym+ykMV+xSE8wQ
EFnQmtmp9gmEcgP5HAX3ZHIqsv/Cbq6a0BTlNc8kHEavrlNjb60pdtzDAaDrwT0d1OGQeibg6iK4
j+5Qfv0wpAay8QJILb6AAUiHCaSuXeeqBRfFHr6CFAc4wjxmq4pQISp9jVLCtkENAXYlxLx9DIGn
kXrvV2vUpI8yfn0LKFbo5sgANOJZXjTOXBYHp3GrWNn+2MFtaVn/DJfrzrQ3F840+Hh9xmKZuZk+
tBuEppu8gW8+uSMR3NpL/5pl+oDGYk75ANm6Y1BbnMCQ6wEh4tS8GgD9VtASy8bbrUINX1zcZt53
YhSte/tBs2cdZwWNdVbExxF8SQjXgsMwY99ishqdXRYoFf4WyuZ/vg6SXxKehUypItE7xQ8iWmLj
vOwTHFhKySTLRUbLJy26iBSpfWcI5W42a+v2DX7ew2nao4kZmbP2d3zTUaYRS++1tLG25+laAHCR
SwqL8gpqOp2QfBalr2M3gTBjAH1dukij9Wx0hbQPvv0ks5N/KwTNhBJWEoJO+8+rBigNBMyb0iWb
mFhf+CPhcWx8CI7FBdPn2DjFB2kv3EPKUOIubEQv0M6YC7CrCbJFuq58UynIEUyVjUm3+8b5b/6P
clFQmTbkalWu2HrwJgfyuReuzUIWnVbjsH2J7GLFwtHBM5WUbjV/NViSDyh5FO8Wkdr173rflJ89
tctnAVHsIyliLtUpM6CghXND/eu9YFLcKicJsXelC/XiB6NjjWFM9ntjmhvIGyCL+NQEBu0HVpKK
mn9dCb5v9Aaw/GO6SAzPsVJRCqcvlAXJtY61ZyQs1mvJjXAJ6WnLZXouxGbDIyL2Q+FDBBBz5/C8
yZZdii5MsjPefGFkUYjGkhbJfCxYMPyL9YGUyyTsIzbtx+rdX/nfqtc9hKOSUi51r357aeEN3BJG
kBV6ehcxHemmXzsLyE8JWov51Zy+imGQScmyL+aLf3qTD1D1r4PBI67oykph/GK5uLkxj2yrYKSs
NZFVPJx/G73iSD64cO1ah/D+0jUdHH5ewF9/BUBynEVdeM4coW5sul9wmNr4I48yt4KV1ed6Xb/G
fTCxUHEIa+Go4p3zw9i2bHsKph/wJhxo2+l+GmbfzsP/o4fWNDlYz/PvLFLKGN3u+P5HY6IJJNBd
m1A+ZtO7E30MMNjQ/IZ4k7VbUwcRmaIoRd9spRwCq5pFKIuPL9CBuiMJUN0ccqk+bX2Bn3DPeulo
6BQ3O3XzILQu20+ivakO/mLX6byYODSgeNQeoP+9+/MZ3o/x1YUUftiaNnff3m0WN5F5i1xk2ObU
KcIIX2WtSwLw6Fp1DiSmXGfaKW710EpMML8445KT5z2nrk03JvWyH4iTw/MORWQjF4ErMuTDxVW3
bWbV4X/YtYY/+CwEjLQBWc0RxHg9XxNOBaPWFIbtipZ57EiJjERPyYkcX6aFbRs/np24G6PyEbur
CdeBq2OcO1BmA9H2lroq796A95oP1wanJt0r8nq/bOzH2PMNIPSJz+9sqjZG63xKgbvAKsg7lDeZ
JWWtv4P5yvizAqrrKaFDMWMQYRLgNVOf1hvF8ucJkYMR1tUzFzSVrFW+N8cHKMzqsT6f9l9ve7Dz
fBvMZ278EEA/yrz4j2/YyWTT9D64F7z9WZk14q0IdvHo6Q+xRWYWuRrDlaITAzGpFJNupF8mErW7
5W+jDoUoPj9+ZU0vz35zRroqU7I3GvR5IzHH3tSnATT2OHqGkKTiOrdbWJB2XzujUoKJXfeQoFMw
l2gfTLIsIjSUcS7aCNmqJxOSnJwKGBzJYv9ZJpYf5ydoiz5dYJbKsNAPFsnTtcFBmojoDvUx1XOl
RRSIY/J1vllXq9FCydz1xGakyy923OHCLSJa2EdGLpUY6tPqne8rCM7dhVX4Agkz91stuWicaryZ
t64C1zKKMMmG+JO4/NLuiK1+zLGMr4DQaDXwQLEDA5qshPhsNo0yNlo2JHPHEkWEsJ/XZ7h7fyNw
PHBHP3slAIpWzAizHiECS2SchFejkYLUY6oF3h3XJlHacl4bpHNu0VYJhHen9L56tuvzDWmKM+33
+yCtHRyYqDJSL+SW1lVupD9xqTMmtecoKxYDEBFKmq9m+7uPYA8hEeIDKoFtGDYzj4o8W6Za7Al3
W2u5Yg+biQDW6/qfGMbR23ekpKAO/66fNhgi1p1xvK6aR9ya6TgKWzGdxMn3RJqaaqM/m8LZS4zU
BmFLHh2kMkcwNWiiWzVFkqzm9uuv5K5LW8KRSb8W08pf01I29X/QJuExRLMvyVaExyWqzx3a6Hkp
qdn8mwNzSEYPTtIEkUog8qXgTRDPULROLx68+ztytQlogWh+4E6kx/+sTzAkm1RcuJsLUe83Mifs
88exUamBKSwwudd1u4HwiAISWBhA7SuDkkjRqfhZ93P7YjD+8lNPkLwxwYTQt+LjN0kp73/AFjp+
EzQ2NTgZn1ve99IGzPvdVnOlnhc8iRQrmHnfQecCbF8WI2tOVkh6oVGp4WhZr4CHNpkTP2KgeRPY
l/mB3TCxJg/s1JYgkz7+/qtLK8qLiDm1Zr4+vSPAO6blhGKMJHXSwAyrgC5bc9E9uScMGLdmRGSr
zBkO26wNGAbnjh3HfpGhJBNLz2PAvu4wkIenFZNPvA3aT00RXrN37ob9embmIcEY8GcWeC+O35QT
ZjT1YfAfC8Q/hQNctRjUU9tJWlxIkPCmqBxEFNS7csNIE+1pnHI4QsK9vXXoI8CKra57GpKdwY33
rL1QyreSMBBqAQ8AuamNG6qMvX/ZceHg6Rfswj9cnt1yWhhbe+QLe34P1EKehIb8DBLuUh02T+Ty
97myCw2Zpd5xwo4EP/10GHxIVNFERc/i0/2lEzx0FhnE6oOQ7jArd5g0OCClNQI5K0fNaFweYLmE
AVrNZWhfbKeXIT0qCxK1nco9B8M2PBXl2O73tUgBLtEw359Hez9o2x4+YWYThOrFFgcwlxn7TT1m
6v5sgBc4VPMILhC8JWLeaDecCX7Y4jV1gmN78Fagac9RedhCLtQ8X1v9dKSa5gGG3dJ6+Tg+oY2a
nral1Oro3Fdyq0W3vccM0ndxssiNHbvbm868meS0Z/cf8L/msxAi2FZ+PHiCKoxhqnJXsEB1CuQl
36lAZ5dFpNlxY60AjEZKkA6IyP9BsOdaBziKoomsNaD1YIYZwExQnUfjdzNvB2hgdMMBorG3Ij2s
2aFoS1YywkdzOzewBwQ/8gTnzVwPyUX2IiPS1T8ANYERCSmc+nd0s+gd52dbsSziWbkxdGsUrLXX
SuWpxyuULDlkFXSDvn3qpYf4szgtelhbjnmL9OsNAIpCRFKOAJ3onAnMOSaKaGqKAtYC07rbSazr
kIAV0ntTICbbqdBYxMKF5KE2WnXiAPntxtW6gVUsU9L/mqw4WstiIxLsjH/CXyMqhbMIXR/mOcwG
aTICwdg9vf2fPO6CTeTbSBAsLWX97JmCPDgYDXijc4cNFG3nrjE3LFkTnIOFQSs5sUfhUdlkaUiS
dCj9g3G3ZO7rLX0Nq70xu+hIHufcM+AXDD5H8F3G+uNwdIAH5CWo1aQJ5NOzHymrfpr44BuEAPo4
+zX1QJeL+AKSxmYqC35dPzH+MWM+HTYlm34XyDy+P4z1aT/1La0b4Vy6OGlyMyYAYTMG/fcZUeDe
86MfCQkX/R7zopx3EVvtek9pXPQ3/JRsCW15U3brgBAPsJfAzlnqODUwpGy/y7A0d2H4HJfxrUVf
CNTIa4jQBVA5PXtTEzZQu/UBMJcmDf+UGlCzuwrdDS23v6Q7iTGWhjZd2FhK32fge6j4h5kkC/q9
YI5LTFOAzRbh8w2cyJy/0xtRkzEpEr713Dc/K+kgFJljv44eyv3QHJnIIF23DmgYU9oZg0LvOIof
x0jmls/UMmNeNRheWrozjbGOGttANNAMi9Q7/jZCxmFQQrlqLzzZ1dot+2l0NzxKiKjgjKWHbL3b
RdLt0tNIwFdbAxs5/Lyd9DQY8WkEdJtOKIiw1z8/xyCMOHT/32MRBqu9w7ODVV5L/H7Llb9Nc8LN
k0e2iqov3Sat9zX5OVv514XFsncCAWm+tBEvQmj/CViogo7v8ekCGUtWaBl8EQkTj67WppNYEgnH
3BFsIbkGrgQS6Iw3PA+5dyGmcSwl0TZzWvy1oajqb/rz8cv0341ET+LZMKQEcOLkD4AVMtQWglNT
vAb4TXBitdjbDZWuSNTT7xqziJNuWHRnevaSK0TIKluL1NGg2GIvz1Kxo8yO+apIPE8fXRiGhA2t
GWYaYHAo9U3INPK/2enT+8YCngujwMsXZOp1YbZB0l4tHEcj5I+Ld5lnMRv/uIG7A/rKj0sPdgP/
gEBIYmSIS3pbv1/ueexDBIw5EnkIRb5fXxITUIEtXA8yX7AszYuHcX3Q2SJJL66VwPGAhd8tdq2Z
dvIH35y9lrZtcJpj5wBXHB6DhkJyWp37DUyq/L4+D74Ik5eNFxjONDvvzs2m2O+9qBM3EwgkDg1t
7St7otKts6lmLcF2FWeu2x2Qs0v05Jz6Du8cp8AkcNsg++DZ2VPtqBtZFP7hqeZNdWdOdh/8VBdg
9U2HBC6CD7MdDa+T+OJDLa50Y1FuscoiJrIGwuFIDcvGvX/lvXYxlPyRlJdypO6nyfwXVoRIObrr
nMYoXsGw0scoQX1x3LopEv/mTmpuUlvAJ1ty+NsjZ7lkUTYZJlF/+TGlb0IRYs1PtqWQOl5xADsH
RQDf1xNMxsVhM0UjdcVmT205gy2Tbc13/5EacnE2zWmic9hqvbGX8K6kNBGC6cCggJM5yN8Wyw94
lFOqDib14FYJDxWpfpD6gza6IE29qm3U5Co7WFSbBaFLsxKAhRCxM0AnqiOFqtfKprlJpy6UWC/A
Knh9G+fOD25O6kNK8NCz7mSnPcWn7o+rHclBq6QjBXRteiHQIPEf/q+MBPjcn00pU0nWiASd0P7i
WUQcWQ1vyrqp2lahMYtgHcIKYbfplhd/XrcCA34+X13tcIhTUekgSpbM4yQIG5szlMK49TgTOX+t
YURdLDqKsrWZgXw+0rsc414ev84BjMmDu1c6evKkvIN2H+lv55ld+67/CzofjyeB38koGWFc7uA1
Uoq6t3WI2ORMvP+yNlNVrRKd9spMtyouOZC7vPOPu9hsvf+DG2SN2Zeun8inl4MrNBbBmmXLHP1h
85MusB7P6HCmYphkJKxshkbS9rMfa4wI6J/jx8Qie4GguHXLjKfSkwrf/ABhQS6I47+ioQ9PST/a
T7rj1Q4WqtWWPNTQu4HwR6xyltsMTZBQ7Ph2THcJWC6v5JtRhMH8x6HbukRkeq/DO6ZAZDCFfVU4
qb//a6AQCnfjTYVmc796MMjSNAvl12Feje0F5pQg6rPqv9ChNdl5yveHIMTpTt3zuBN1PXbXf9uM
oX+W1arYaiz+P8Rf1qluXiVJwiwNoaS3GkqIbwZxmQmlD60EvkpdKLoS7K/uJMZ7imV3pZvWgAnx
+Tp4wMvokaxk696PMMuHG9jKVg9aBz2wiOKvz7zcEh9Gec14izsQHyVuzwdzIneoT3nsTkM7FEG8
mnSC6pfGFNgHInSZEBQQX3mrUE244oOKxI/FOPQ26vskOsQgcoTe7cM61IlJ27N+CBsH52pP/boA
syPiSc6mzMlBnFH9oBh7xeR9S8rluBmN6oTtUgYr2x8QGZnG/AXCTg4HO1wYCHHwNblMaack/3pm
6zry41sveAPZfDyCgwOolhWKGdSECsp99y4Y1gox2V1SVVkfjIdrYxjGnsY04nK3L4ynUL1YemGB
OhBy8AIBmzQv9cPew4hhv+2p/0hWs8SpZyQgfr4CmST8TkCfj2btOXPgDKwewSZa8gP5QDN+6rSj
/IUkYQyNmCKMIunoOd7aAn7V7SF8aNbXfcoDKmnj/T0MdB3eKhF2W5R+s8lmpr9S8ywiYkkZw8ab
27NIf2cgqH87b0a1fLAgg5udyhO9884pduBnL4PwXAT6bJaq1Y3BtZXsZHOkOKpIw/16+8rW8OZu
S2axqZOP29ziWV0SkP260cbkqSJw5EKOSB6C4ZMxSojAyKCMnmTMTvZvOiV80jZ/5x8HjKIGabzT
sc7MlzEuS0sjL9SgRr9AU6QjvOCKWdJyQ+lJ26aMgDNVzjgPMU3i93SOvcs7OSqk32ut+OOl79te
qufKIBsdxRJ+0GJAJ2yAqKnN80vBjMUBwft+jWwxLho+IYXB8dfc18LrlEd/DdsM9s0M5lK4U/gp
ddSSBxJbD+6BNv00wr228YjIx2+0Ve6pAQht4p97b/snVlvlIO97MxXHGGHF+kocrSuRQgF0r1AO
UntZ9cw6pW44ZLHGrpKVIwB8tMGejnYX+aK3P80gUmJEpHRK3ItTacQagbJqBs598YrV1tRvB8Md
DRVSY9/kd/6yUMkOn2uZUKdMAxxsmIbvglmCcoLGE4ur+qKQFDuXPvTSSA86TcQW3k7q+E4dJW9N
ud0bVLgJAlolXjEntQk4wym77dI6m682nxJYDg9T3fRjjOvyp7kkoASuNP3JRDa+45oTKvHKZ34B
cmThzhUiD58E2us/aa3aHqB6t+EnjfzHAoi3QT2e139vBFbRfz7REgrPR/QTLDYDLYUK5fyIAGo2
YRSTMqjc6WjsxV1+NmV7e1Adav7gZ7n9PgvXfF/O7UMHPdxs4UQrTX4T5NqeDthyRr0H4PUXBBaf
yQmn/7zKvwsxdRCKp4NevIov5qCp8TFxRUuZoHFI8HZVS7Zm4f1Kn2lZqEBUqIwJnU68QpUgvine
ZM0D168nOW/Pt8Kg2a5e89bC/0HgQCX6thjFEITIUdk82jm18kVoRiUiA/GNxQIvxLNhbzkPvMW6
wMUYo8x5ewrHKeALHMzQxYtz5Nmqxyh1NjA8g1D54/85TO6YSFML7kae/8k/r4HDnd7kD9BZhOCZ
rEBgVBnyI8A5L9NyPBXamGne1kp++JIgf4+x8Eq8gvNGemZbgSWGyprJC4HH3mTHDrM32WdPFthS
Ez97ZHkCjrIoMuanKL+bednhs7iCcDl561gHk09LlepgJoMrfnJIdsRrRjKzlTwWZ6JbthFqrNN5
AvOlSUqN4nRelCHmRuNg9+rgEpoyr/umdPN8c4Fytvf2BvQvzvWgoTldIjAwyhgxXGVWbmYoW7RR
yRT3pekt9V+JaE3E/G62csSUD4HvqFig76b6pQ2nUGZZt1xjq651JYG5sDoZfUhOcgdscWJeM1he
By+GpyljBhZqX4EjKGpzurKDuJAgLhYlcRqoUGpTa0asunwE4scFT6aiVMki8m11eGsobqzY0uLD
EPG2lqJ+76ZYaaTZNdX/Oa2AbSTF+r1JRD8zflHOVLeW7nSxEmaUz+Bro3vrpqwV/eE/vglIe4he
IO+EoWDFtt6meIbkvHWVDm2Sn+DPVFVlPhG2SGXIisITur7HT8uAGRaEcqOXwxMyMw2qO/U3dVGO
wUT7DcZW76XeLJTumEYfKqWmmUGgWe3UyUkjzLni8lGvOFtYWOZ4m+SWUGZAaXyuZA8sarawjEoG
j6dze+O/2W721VaoNB1Wz1tG34W/MWo44HAmAv7xJaJoIGUAT5MdbYrOb6e0MwOOyM6fsUo8ipAO
BbErJn3MSPSrnAQ3Si8tKJT56Nrvwl8Oh+v89pwsqZk7IodLl3GKkYpN+fD0u2U0ONVaGlUAAY62
bPyxNRDVmMK7V+mLBNCAQWTxvbQlTjmThSlZlfU2gA94ksvITj0P+YhrVv19H+tnHrriCz4YpXMV
w14oGOSTFEDnP3OFIMqXprQSSFMSorSlvtm2732saZqBIuu45xcXtLlJ4KuoKDrBHF7kvgT/m4eG
Zw7qAX3helW58XE4cES+3ZYc63B3chKF5odwKcUrMlSxXuU2PhYUF25VDghoKsWFwENrQB7envxM
0tRCdhBchR554XBfNHTJeYzYIs/u/ST1ghBfFix9fIyUzoiqzKxum5Wt+TbZwtOz3NOBxRXzYvii
D57MKxQUvKspxv/GTtbD9ugaJ7Cp+b0lwYWlQkF0rnYDhI6HgDPBsoef/urOu9BBFT4KFBVe74nt
jx5L0LqRGj2v6HT7aDV3ospoyrlktFyhmHxgTDmEGFI/RpZkROjpGIF/Je18miCUpxokaeoqY6cr
4g4qt1BiquyuuXH4joO5iChY31LTeqQsVb3xXHp3yf4CmGs1Yi2KCEo1YZmBBMfQOTd3NM64dpxI
q0lbcgr8OxdxavaOdWUawwIZYJXeWSHtxc1W/mak/n5n5oag7VvMiCNTj/QWqXhUJY/VYO5ycChT
FLYcRvpaUv2pFUxfxODiFzLF+dFmtB0+DFOInyTVcUIqSC/fz2AoogfPCNshBDwK60i0u42J056v
RJj8J5fUNy2aZODYUkH1equXr1J2Is95NjfyJwkXo++vxQ2EGzUpvHG/Cu03XGuboAA3HGd2idfZ
Bf607HvcfReoFSrFBKwSdgn97WAAH5sgP4NI11IXcvFoFrzBfjcpg1u2u34xVVQ0FTZ4/O5gtE9w
hQBfbVW9XIUsgt9loWKcKh+Un3sCDjs6bioASQrBok8E80CqXew9WIM6z2tdF09LYjEfWeky2sE4
UE2YFYngMAOruKdItUX0c2+qv4J1nuEWdDVO3ab8mtDtANxEGZE3jNaoBUMPKtshPQ0iOYJZVY+k
8OQr9p6vNrimnnNLJJvYgEM6PWfMfUUTd8czIeOz8YNwJk8lBiZdISL83nOSH5jk+MooxkOxrpLO
kLLGAwUdCIOt0bMzgYGIfZhpq7IMlQQfs772Ki0Eg5Sej8kldR8366oyq6Y6NElrWIx8vsZMcvOB
SbQ7CHbei6kExEve1zVPU/fVQgmkytiwb5UEhTin5m4IxlfJH9GIhFi7gWFz+jhxT2A2sR6SiZJB
ZHxqT2oJ8lQtHgeXJp3btlVfLFnNrCff45PsK2rEZwEDmKef9hioiDhyYT+A0Q7k/4Xf7fCBzn7P
TfXcBHMm4D/gjtkzN4t+kQ4j29IW2kXxJHQRqCUEyWUK5EG5OIGsHCOczX6gdlKiakq6PXrqpzM0
k8As5Iubv3acnE1ILv4pDQrMNOHG4fU7VNCCEP0w859c8xPbimLSZnoXF+ttjkX1jrtDltgVY4kE
xBX7eOEoqyLUqC0xXnIBe4YdLFwUqKKMSOAS4oZ5Rh0hV58uvNn4lLaa+a/Kxam955v8BQf8Cd2k
vnfykR9dVMtndj6lBWi6b5elsRtezCl+MUUK1w2pz7HinLLI/7SJjiwtU+KXShqVjZ04PviP3u1q
/vqnBKtOgGWhL1/SGeFZrerFS4Z41pAids9HlJHyotC50BknmkZOwhFgZBKe9fKrOjm7pNb7A4dd
xznqyJk98FzU5dWk3nMASlkXehj+AzFFLKVKz3WJmFKrHqkyDZu77WRvhp8CSKKOFMooLCRNOPI1
s+PzbBYlGnDpWT2mGCQzwTkz/w850dZVqdHYlNQZVAM/cu/w9MqbcA8Kwd6ewQpvns0sS2igD1iM
iVMNbTYDXqeNPRKt9yJs9yawrLDkqTNXWVrvHiRpESw3PfkW5LW58AWP81ZsJb/UOATNn7SVMrJM
H4O0wOTLZmU9JF2OqeeCxwYCwP9wSuPWMOcqz2WC9bNOteQNoFWBvCFQsR9Lukp2ufpi6OiV5+ZN
TO7hC80Ez+jGnYWfAluSzga+vPc44GOF2Ned4+7NZG9GzDjn+w0DD092CMCGJCvKM/v3IH5WfC2m
apmWoIUu49rTA1wk0TqXcddo8ZHq04lc/cUvv8HYeHbDHCmconYz85Njr/bBFcpIafCJ6JfQ7C/0
lMW1pDXj1WeVKwJ1pa6uZb5pYVpNx0OoBv7hUXce1EI1AdMT4S/hRntDYURNY2B/L8rGXcEIugrY
ipiPupwJ/SL0nUcdwpWE9V+G6U6jKPHhyWCdfPvQ34lUA3Qee7r4tlUzr1NoWS0Ux58OK+FkKEuK
G/5UP5mWDQRCHyFG9Kjnil3mwqYDjTqpzDClEUrQ1BajNPTSf8o5MUlRIzOL8+ncNzdQnjqdQlnj
RLgvAqJy0/FM7CzdbRN5rUl94vvb9KNjOdRqdbXHaRTXaxiOQP4jUF1lQlov0Bo0eO+odZMCcSzT
UHpZBvxKKgkEuLrtKO+3GtM7oFQWbKCBHtX3RFjzAC1QgaLggz1crt86hMa5MBvksj+V6gIx2PUj
c/fmAWhtj/ordOrOZZXifkdO4bop2bHOtktOPMaV13N+gsaH2I8u1K2CX3+YtyAPoO7pv8TdEsWp
/zzhaYwqtDV8/L8QgyPouv/okMGAmpRD8KZbua5DwhwnTepo8U/kNnoC4s+KBMpW6YE83erCZsaN
ccBlTuK49GRKz5aqTuEy7BwuAce/r3tUXIrCAGQBrRSYQpf1PoArAKqPnmyp5m3Xw0LGoSPTFjbB
jJ0r0CwTDYMOnYf0Rcd60as1Bp3cWnWNbQVEhlAaEm5O1ZDrwRiJLgIImj1uRR6cDXNLyXm2LPGe
UfdbWhPi0PeloVWKfhQWfhKke2x/raoA6Uxj851jydY+3smuUNUuZg25jmUuhda3OzgPB6itxQag
jeyLtNIXs/DV3rMBwMiAo9B34kmtUlNRsj5c/KpJ4lIJN/+EPSh6JCbbXUfGrwbLL9d6HYIl5Psm
yfu4QRkVGbXJ/YAvqZEzwVDB1fGh4h2hykCeLGkQ15VLT9KONlBG5xzpl26u0itx7k4o7jy61laq
orcckTscMckZ5Q13X/6QV/DsFltYGGb1P+hkdy19VRSnvocwktdDHuTn2MCCerZrOfScGJdQFN++
OloNP7kftT7jlS/XasFdXldMLCJzP8K5LgEHRVySAjYFC9xZTnjavzQE6hasGucAxUjPP1b/RZEl
cjd9P7mFShM2h/uWOelzCjF39B4cfsb6KiFok8Z3PAknnEuc91K4hlobIOSTCFf3OqzoNauDh6LV
vMrFQ0V7Ds1FjTrcN5ARQZc3Z4mInH83XcYTAbSDlIFXhhGonTeUQR9NlX4BIPDGi4pkN8LAoL9M
Tw1siyXqb2ly69Q7FL5ZCNzsF6v6MbdBPHy8IhLuer616reYR1sCGDzDgfB4GOtci2XAgjua2ZZ9
k1eYcLeTTqz21PVXDzMomMeB+TkA93sB/38fNZebi/A4etMzow+9nsAa3c5gXV1E9DNRjCvQGsNJ
UdB/hiqPyWHJZ1/aHInFjHbYg4uNOlUf6FqrjNUuPlJkAIkwLwd03x51O0YZWHNe6lnuCS7vJPXA
ndumxNA0dAE1vWupeJRSBRb0HZ9aV9rgEEQlTankhSoEJfk8R/H/6bHGzteJDsbs21JFhJDmfj6O
8ldnqERQ8GwK7KITMHJ2+NbbJy9NjkOjAWnXWEHoqtMfSOF3TV6HLf5uhHZgwKatb7uf3UXtWvI7
XF4gBm1eq8ms7XPczlYcJzVRDyEfKakQtvx1fmGS5y7uFVOc+jQUIAWi+U2ocYlwX4GdwZX191rz
X31wXeXKHue9e5a1NFlmSyHAHXvHlFNT0XaLEYBv8Rpj8akXBP/eUMmzukDJJWyQPdmotjo3CgqJ
zk1hLsLV0CEhUUTNlpwxsxinPGebmRmLFo0OD9D6khp2OjclfPTE3hJrAHnXQlDDQybfvBfXpvhG
CA/csw16D+MzeZGP9qEDsyXehKA1BpSIZjUxRf5WKKWDNPby3dlsH3DIBxcTwBtRga/DDXp6seCr
LZzzeMPmwOY64XLlJwywwGTF/rlpYPTt75Kfo+iotUBI5GemcHASx7k281O1UaclrGArRUwrUlRv
yz/kc4S4zuQW68u5xs3cBZdTEmlppkW8R1tqwk2ZvjGtsx18OcT5qkoz2GnI6C9tHxTqWz60Q4nl
rdgpnd9ZZWSBu9yl++84P6cgML3K/UTsgOTh6jm6t0YzRf6Ys0Tsf0VYm36XqVzBA7TIQTOXkoaA
qbqji3ZbaPO8EfhZNSHIzBe4srEDzRDGuTEeaR/b+Ag91WX5RTXORKLri2ELskInCgTgZ6tDxdle
a64Da+Vdd0nHqPck77e9LGapHa0Uh3tIf9mXjyeTqas8W87LhJcsdNj537H/sDKSRhgr/2qzUxMr
yG6KRzgafH+Qrct1EWqCEhMMvbQC7fhDjyGEwprtadLRWhlYE9YF8IU5/CS7JmZ/bFHv1VMsKJaU
BESlWW2FTs/0HXVhnrtcHqINWGBKRMf6NINli3HnCLjwE2BO9yuUKrT6k8JgglsqzSVtR9pZ2xRX
L6LF0uC9n69RTPMaUqYhUSxTpfgJFao+bU0ZpASz78NxkT8np4Roh9rHtptb6rbwfcIfBRh71rVK
ORD6J6dF8nyQVsFMnc4qnDUkST43DOC5QJkBvB9jAhn3ko0QQrEKCt4eZPSmFESrCLFAdCZisrfS
HquPuiF8PCLLXLgt48pGfOPySyUdX0zjCNr+uoy5B0xwyIan3jQUOg8PZQxmWZ1Ev2Vw9cUBGVLt
F+MHB5kivTdSOL08+uPp7ruPCCBuZXL6/v3ZQPPn1uRNUMLtZDvqkj4FDHaHGVq0wabLzQxGSOgX
CRDoJIaJjH19sCxQ/wR4VgsUYpZ6VcN3QoE8WjbRyo9GQvrERCv//TDJcEdaseq/A+Go4rgrwC6G
cfHvJpPpqG0Ujx3ItXM0CkU0VVFdHzQNeL9wPI1Jhv8erClgH32YkYt1fq5sFKdUzbq2bN4T396u
o8m9PNdOIk6xMdxcAOWN+cJz1mNnIfDtzrV3Gh7xHF1cLhaJuJ6bWUNwUMNJ0AiSn56z1TGRFpl9
CjB/1YpgrqQq0cXlelZ69504VtdwcpmdvIQw+Ty403wyIAOwCGVIxUH6nRVtZHx2+DwFbLg7p4Mm
dFMM+xiK/0nFtEkt1CuRjosxELVjmAdxSDnQqHtu1O6gLx06y87Dya9lJi1+C5IdD7kDIMOZ2c3F
n6/du61w9ebjx0fA8dVzSF09co0BWs4ZwVOVmhXWxg1Y44Xylh2YNGX9uhoGHtPx8QMDHTW9GB+/
QDaPfJNA6J4YFb6kaCjo+tGHWgJKMSuq55kUfn/0sBEae+czvv7fZAGTCDClLJp016KDeO9iN6vM
+ZfLa7ntTc/sZ5tRcEwYszCCvR3JtKrH+DM/Dn0faedQNc0XjKKlUp9ZtZTb9oH4c6xwuVt10FFE
ERt5Oe715SD2QPlg+Z9+HUKNZVdzM6yCC0PaXdHWRt4RqTQxLpUjLXkLE7sr5m/Yf3+yUcIt4zMQ
9tO3jor317dZMSDAa30EEEJXUhPx3Z9m7+6KAsrH/wqNVVjpvv1hzr6maVbZDv33DcIZL0j8tvMl
zrIUDzCTP3a0tLPCq5QsgDQXzPDQyru2p1yfzeoWkwj+vr3fIj5R1XT+sgYTabYdmNF0n1r1r+np
+uIUZceaJ5uzG1pavshIGOqkwPmdSfQHkNUHO7Z4OC9eLf+0kUsSHuVKK58UFKCd41+nPimUHR65
FBIAX7aOktNL+5Qopu9mtn0+uWX4WMAt77HVYEAEwUCg+Fu/cKa3ncHeOL7AyLu+hU/H5Ucp1+I+
oDe4nKCCBZdlbblMjhfmPU8kw4YvS726aAhHcJ5j7WUxlLhI0LwDCMXLpSqOsXFywA9z6KCSQaJ9
MIkb+aTm3nce34IiJKC5/I61be/oiq+u7Yax1jT4TPjPDSNoSf5+TF+NGE/vqgpkXB3LTY+D5Qp0
jZWMTPdBpHAI7XQUbggjJZdSfhukENjhVPV5fx9DtW3fJyDgcFrDiNLzmuyrh+GckB92jS1YeTaY
1JCaL58Tv3i5lIffYLiwCX1LB2U1HYHt8RJb02dffJOWN3OhK7yuXPMYKp5a32NDXnxVwoyrjJ4B
3k2JTJlxFIMHIxe/5R6kwX0D8DObm6EAwDXtMeXdgpdIh7unTQMf2OkvfgxIYkJpDMYw2VCWz1il
3SiND7L5U3Nv/wTeuejqXwJT6M76tviu254nEfyPBazLwhkcd+8avb3jtrAiLPJEoEeLEA7/icPp
zFLrjl2Wkrk//rvz6WLShU5UOUfV4XV9kSmJNyPGWwW3/s6TJXXxU6V+RFT8tRQBhLM1JBUnmV6o
SV1SXbMboCOlqsEzKZl13DkFXHW5SSO8I9EOJx+XDEa8VspRwS59pHUeRrmyyV3U5R5OeKA8yHZm
EVJar+OoLj0+CON6yLjfLXSAJzj5Y9hzGRPsbdL4Jo7vMh1bRQkfBXeOMHFp8FZnBDWKhaHoDR44
bwal3yFTuNqWCo99qxlfOeCsLSS/dhZLOndKVGDkZnY/J6q95K0MR2lUHiC0uLWuq4z85MvCp0rV
1rZEXSk8/wmbptwWg7MqhV0uEgUVBOJYTW15W5qA3v4jgVV9/TVXUC6+BWDD3d7M0UrMOt1cP9y5
NtM1u5o0PBtfLA+LlzaIjS0VjyJi/BbNN+23sJzxhBVixSYTF/DIZLx1kflZQq72ANPucKwYbN9s
dxVLufrO4vfRmFj5IsW4fsMwYttW3HNQoDb9xJujK1SRD92dc1wlgHjIlsBmnx1B00hzhJa9qNsi
i8iYZwjhshMCo5akaVzUzFaYXtz7BuaLazAsjnjXl+CiydnErDUtrOgPIwH3ghJrDT7M18FmitwB
qsT7lNPo0nni6xy9TXDvRjqLRlVWkBzrD1PjAJj+MtwL5UqYoLF3gDGAT+w0YiWLqklK+CwdVjl/
IyeDYq9d88u9hHfLMSTrdvkkY9WGagxtKCBHr6bv+cGGoSxaDvP48zhVE3nT3K/RjneM0avPJxdy
V32hGR/KEN+ugWVFbcLbV55XB01aR1NOUH52TuPSrIpdJsGZDRbglhn+/D0X9aNM3cM+3GaPplOw
+sGX8mzOG2Lc/lHAuOl/ypNqEECAw8rCp/LAxe9CpicUq/JB0643w6X8HoaVvJ14je+6TC8WmJje
3vzpmCsrbjxIwMVYZY8FIDChbRvav44DZ0aU1fog/0iPVnU/2iDeq6RSqNueqEWvCXydjy8MRDjW
fd9tQK95n2FfjGYv02bCVEZRgkXY3hxcCZcTFL245vYvDD7FJje3qoz9wACeGL7bv5AcblwA/FB2
FJvCXUdJUkL/pVcCx6D4I5SfoQtW6Xw9Oto7gpBWqqlyDFwnRDLusfoF/7h5msKJSpWAV0F4haSW
cZrVJfMSz+riRW9TH+JZOYR6uEECBVSF1jusr5/BRoUT4oEhlSfjvlv4Q6dnWdA6peus8FpwKM1B
FVfMAJdr2x6hEyx1htFEBHf2kMI827NFASXtabhum+2q5lAJGKuiwE75U5f+q70EvfsvgpmDQEGg
HlDNcfWcTgv+XtH9NZajaYATdW04OxSLC775/wTG3+ElZj0ZmSWqj/wA/aTtuiKVR+ngi63s5j8I
z17ZOs8Dm5Yfp7fdDCP03QqSkleyf8qRkIVf/3ndcLEPr1KzJZJ2DILqeaXFMmAW4DWFr1DG0yI9
2pRurmQBvUCYup32fOd6rKxikL3ysKzF0OZpo21pHR+AlwPlQW1wmZx57nI/LgSn0HJd1m/TkPm0
vQ40/GLlaVecmBZxuMuFQvYlR2wr1KyqUOOJCAcfup4ero0rOCSTITIYKa3Vu5Lh+igYk/dzEbyZ
i37tQTzxRGQEKhWoC0eufsqgON/f4sKqIqkHebKhTEO249XECP1MItxWPMMNzHQmrX2+3jQwgh7k
mWc4U6WdxDBI26Bjs4bEXekxvZ0OvxqS6BNaWlBbdhAmskz3u3OotFJPMZOWvlKzAOD2+0bG5OCC
yp7KYWT4E7l9zEOirTYM1N/JNYJfDTNlHcsVs1ox8aGBt2A70JeEj0KxTkNnM9wYh3JqYw1+Xj+q
RA4TdKA1Q9NuSVtw+pg2t1DnMg9+C2A6fN3rw3RJttw52zDpSWq2Ip21D8e+LJOIwi7/PGqtWtQ7
L6NO6j+nrJg+Bw0hs++YS4TCnijObbQq4aDcDXzmCYzlsMzCDIA9sxHCWFwyzXNOfxhzeTpFzJbo
xOoubj5i9Lj3fGHc+3aAfZ+6C5TZ5bt1h8tac8ncmg0J2o4qWq7Ym8ndvM//Fid9v/oTVeNXLzC8
7UriaiOAnj4SGR49dC2v2EZSzX/3HnQkIkTQfjvdYDC+TS5ZUgtZGLrPbQg/kgejIXAhn+EPSpbL
NKEavhT5wX/czutAWu4qDovkcQnIbDf+ujUnau65u3EjkWMxoO8MdgdWQuvZ5cY3C42EgpIBQF/E
hOywQ6teHbodTfinla+2dybOzIjCvGFuGBTK3VBjzUre50cQ6t5uHzjGwuyhfXPNLSfYQwjxOWPH
wNTGTZPcYJY3T+eWEISJ+UWlaPLSs29odUm+d7JAFc5j92nofrsBQuH6ideRVfi+c/7MjyNRoPZU
7bYg1CLXCaqCDArhdcKTToOA0Sulig442/t9feLsbLq8+4ATWdMijaDQt5cU+DB+tVzPFX6vvNxC
fJlSQ9PjP/RDle+6Z56yPwUCtiTzfZg/y4LHevRTUqQEotGNrsaU/lntPy9OpIbOo20IQmVoI5j3
57FaSNlLwmoGFq8uuGeC8CI1AibyiAVZ5mDch5QdPDRUqCc84t0lIZL2zrwwQwAedj5v4lW0tSur
kDIJWCu6dWeoqBCwe678tzab+cU4mgM6voKco4+cY9zSIBR++1EL9DqFi+RhFWBqB+NEOuBIpF55
E8h1K4iAF2q3HfnnFZlUvMX4PSQ1n4lE1d8jh6jK0tNWaWA1XMH01yn4IL2UH/tKoVzDCu8Q8G3+
q57XmZWDuXNEl6/E70KTIk2ZPAULSvQxq/yU2RlqG5+kzPV5NPu+tSDagjfX3AAUlOZQyKYfsQRr
5NjqgWnTRDoLqtmu2ChaiHgnux0JhzxWjzzYS+AIwWACQh7dtT97sC0knR2QPyu3CxElgT+BFkd/
eOG65TkFa8jAiow6T9dcCZNXfvJyq84sOe6LC9mFXjN8x3Ny9qjt1McydAlOPCYCDIUE9cTwJNW4
vZRYXM9u9IncVsV7MJaMqQGrX9jbxfLDmJOVhCp7V7xPauVncHLNQH0gglOuegmLPQkTKkTRC4U2
u6T/y7G122b+PJV9JpYOI7YD//Rgwh5M2Ha+OCXGhJ1CMG/M7Iv4EFJnAqjyW/z7AdXXDttt7TSK
MuAFj1vy3BkBtJNMMnbx2mVOQ6C9a0ct0KkljOWy7IIatfWfUY3RNBXdZjfjjU8632/pTEMV8dkd
oiJEjoKSXpekk07nVZNJKuV7vrWkljpOQ+3imORnn5vI1Lhslzs/MeS8wz88fTVXv9aGR6N/J8YE
xpgIEs13uwKYWFcLQBQLcUdpACJtAVzwmLz91EmmN2LmyOGmzqea4lU9zfPYLk8Ohomra2DOyzHI
fAV6dTO28DWVYdsxZbNnDhFYXRwoL3B0XwJjMTs6TnxOPreGMYmRXz1XKEYHZFHuOPLTwuZkD1nx
GAkIsnV35YuQEQ0db/dkLyS6vBpdG9fvQ8y2HBegt6bXBUP+8H7tF+gE6XYt7SRO5qkL7T118wCy
XYX+tJLcFf8bLTZI/r9JoXJTCF2SxOJG3AkrD5vfBkBHkE4TYgPDa8U0cv1oZa4kjatd/pZECjF9
3tD127daSF9GLy0Vxezfcx3s74gPkitOgciIoyqtYR+49m7b/ZjpLSdQNfvWEnAZe0XJgseigyGC
1tjWN+Zc6gmIZvRWZBzT1EoKKLKiShhYpZAPDS2iKhGoC1RNzAWxYA88DaIDmZ+kk5Gitpelgp4I
D4TzXXJTWnb+gZBsrkkKvKSk8nMoWqDnWFKEfBLHLa0ouo8KfMV1hxya9aQkLM6znz7DGQooKd+X
oME5AHNiuFaiIdogOkFp/CJVBY6CflhlmMYSdhWSUJ0/BqYPJuY1lPLKjGCe6xYtYIHGe0vHM2tY
aL0aMlmWifl4TB1326sL4r3FVzr6Px7SHzbQZtmJ8oLyjjmvuhxZZRlPmfmK2mfwJW0KKa1YBLaZ
61+feVR5MVoVepV9g3RAKZ7ltvp27A10OigQf6pNEdUZYwoExMl6i+WTZ2YS8OJSuti1QG2bUGG5
qCNcKgXNB+2vHRP2H3vLquCqphNOLak4hTlbCAhLqMLAuYdtKg6K+rrKUzR4886Xiaoq7CSN2YUJ
SzVt7VwVhUSRcyZ9DuQxtTVKJnBLTEOGRPy4y4FaOKOD2GY8as8KrdQ03OF051vPgPFHIErvXl1g
7Z2a+LOf5Ztb/LvlOwbNrXdUst3Q7uU4oQIvl23DLtLYEh4j50hEOaqB15RwOMQu9l5Gi/DV6c1c
dr1Nu+/RJwxMhGIaRJDt5wKAb2rOcr+FcWEbeNQmdMnIq9yVxm7GR61TcfKO8dwvUg4ySWcbBmif
1J6T4JYhwSg9H/BHHjkcFQ4IeibA6p7DkDPH5lTd0eIAxqM3nsW/ZwTOgihxT7gsqujFys7tqhvM
myHvXEfs2RFt5qG89ilWTBaq4yoZv+IaODw8twBSrBBf2NDes869xN+GfC7RSLVyxCQVDJejgtdn
hdXdsLp/2QTuAiLig5JAlBqrWZzF2t2zKVkn1qsc6eirOcscdI0lMpjkXIhzGcW2xtQmlPlgzlLE
ZioyImU3YU0Ru/QQUYiwLOVe6V8Wky1m+UlLlJsvnCm068gPnrA6ISiFHDGxZ2Z+ues620qLm1ou
V4uUaYoweoQPQkYkwCBF3tuZoaAXuWCRciscF2TpigTQ/xryiDd0caADx8QezOa3Zf9EqVD5u+vl
+kuokv76nqGqJ+NPc+kD7YQXrQZObg8RYEF+AHK229lAhfgHkUp2KqEnPAq5S7luxdqKHvCZll3h
P1511Dc+b7gKa+2RApHo5fRfloxmCpuuJKjRyY1ggrWiiZHGDcXUpI/6/uzOtT5sDWN0inK2FV3J
VYVEPScqFPu1fuosi+JMItYPeYKW+raRZU2FEjfA3/aHTemYjxHGfzdZ6hsR1wANA9nF4wnFAz+m
Le1XDH4kQMV9Lk7lD5caxA9Ll+7c7D1PF/0JwpJG5OVqhnHF5/gYd0Px848ljOJGU4EeqQ3O9zEt
MK70pMdAirzdLd7zgx0ajz/Vf5e+x0K+mhu+WHYWpiKE9M3QwjWw8vi+1uqckfEFbi9D08ZS5rj+
5/TaxpA/E9/KVR39CH+WY5eLBwTCmO80ibL6fX9HgyV6VzbDT2uFrgH/2ZCzrZ0USc1VMz9iRirU
VLXbtJVQKo0PoSK3RquICmvJlF5YfFRTdekPonpr16oQs9YGg/WCm4IAr1+rTRAOSJMElBxBmLgy
ejNvvo+cB8zGsMUAUMkkK8KiNG+qkU9yX9CwcQIV35Q8ubeMrQYIIU1qvZn3kQegC1X6ANGz/KRu
8jYFTpHR5cQuzzs74yU+cB25QeS+mbmN4SFURV4FbW80fYS17egAMCL3fvO3H7Jm7ilj2Avj2nA+
umpXbWjxqhCgKN7wHPf89kqw8/sViP32qaZq24VRnNf097ERMZD0B7ltQzMbpq6wIqBuYSD7ZEI+
DFAC6BV6q3rv1Z28XzO3hnEZ9GND/CCFP16DSo8W3e6y8oqUbOcyLfSv7Kek5KXl8SE399BWn85n
++X2AhRp8SFlRD9erDkecRAjHtHJyWyQH7WCpEcKrUUnXNhjic49YFI4pNTnfRb+2N5N6Fm/lhum
ti62d0BoeB5cdtp4akAIAB1Rp2M2dmXOUN0G74An9rM2IpI6+cNwNPhbmhD50nBESCeifbnCUhqM
BeeOwF7DL6L6uLbtgsfRZK4YrK5ngB1vr6qmvbSWgg43tlG+wiH2spAMoNJpYs/wdlFEmyg7sPtv
UtQDql0qGlwerUQrR2jMC70b8S3/YtLeOLZQzdRc4BFFJuvik30M/w6GcmB4RyOcsAjGbufkNp/z
SrKwK31A4a2acYntbxyDpwHMtPvok0W0/qUM7X8As0SVuVYpv3YRYhnjIrYuASLDDQHiRvqBM+em
HTOL2Nz3shu/u3mIai40ABTwBO4QO1IEbKuTKImkJT05OtJ/tKumKICMsy+D7TWeLxlAG2PZRaR6
Zq/jDfn0hVMCd188HVJX6w0vx3WDAS2EFXWyBEGgx6aoqDuOaHX9iDynu0dA9X9VS0GGgNoEGU7+
r8SxjxgnDyRApjW/OSJIt0Io9B+HC1wZExhSvE8CImwpXjNEvLhy8z+SGLg6Msbdm9f3DwCc2t+a
YG2QgtQVtC3aDQtvVmF8y4PLpFTIzyt8W8Gyz/DVX0emrrnOg3u894KBY+dJHFpJJeMNu4/rMQd3
61ZQSnR08MLYoN9gKXqhBZc7JgFDu5Bw/4UJ/rDCxD+16qZt/iKgAASxLhQjx1udCmsOg/pslRFM
XCuPesBO+KLrlsuKyOZ2c3fQe5HZqDoQ8eoQvFZ/GlwLRTd0CiiPR7EapDK4gpLXw5BLtR6UD2i9
PynEizd39DbPQTLFpYxjbEkxQaldYgbUqANZdIqtSdFFBHZWvTmeRTCbTwHkfBEBGMoFaeRWlLIL
/oTXZXp82rm+gRXBNr4+MZA5Bbj3xfYyiwIjWbs5D922mOY7nsmKXoYxICh9rB5HC2FU7Ei5tLNf
t464dvCNwC5KDlxOCmDLTbM/JYh9mUMn9kiY0Faew6YBQ07P11y/fzNrAqyKEo2mqTjDCCA9bi2d
jZlFxnv15ggZiBP53S1HKgEPjA8DT5eKEcuwywD91PAqAl6rQ+OIQae0Nl4hCwoTQjkNHjue6+4E
Up6v7emEcLvAVY1PPske3tDij0sKCYFm1oQ6S6rIVQSoVY2KWREnYZnVowEboQ2LOM3Ax9IxXiDJ
XA61uJhFt+nNLGeOIshgsZxyekvmU44kB5bKcNyF3k6kCEBjOYVHpBTp7MsUPTqBMc7sL3VJzHYz
kP/2wki36sxTPP1mgtAbfrILnoRqGoCPbMCuKSR4EVS9OCjY/J5yWBKXDenjEaE7v5Ik++IHAGZP
vEx3KM/5LnrIZnTTgdqXkY2wIA+9eu8ffw5sObTuFlXj9vdUfe+5NHdXmxJYuWRYDVwwNGvku1n+
GlY2YbQUHkLgYonRBc6e0d5tQENqwqVGRnCqzkAy3oHfXMS2TFKmFUg7x6cGdsJc/9m1kk+NWrYB
xQvixsxkpVUbTGK/2agF+V79pPWkqB8TsgMHckdW2YLocccizKtkdgFYkc0aPNyPNddhMKM9MLyr
XIoFSgMM4H9K1/zh0BaE6Ow00t40N5T5N5dWfC7gPkMpEVFz60CM6GtdFn1uZosHN6N6HDJvBQkd
L8FjD2IHW6D3fGRcdIkqlup9Bd6YTDo+9t91+38Hk+IwtD4z5EC70NxixrABhwqzthY0rquU2c4u
5yEnql1iES27c9aV/y1YMZYDOwC+yXXvg2w3aQNX58u+QoQcg1zS8IVxfrqK5TS7rfGIX+6yupHM
yM4dKe8zscSoduWfc1oamm2VU8WfkR3QsEYwaQpMJGChOQGxr8dLRtUeFZOlhCNkpLYkTf+ulv10
0lXlncpAbVhHiWSDGwmqYy0akOwKvyRETVRjTcxyhYThbWA0L2+3N33Lb6BazxCJhL8dP6r9Do6F
M3HchZEeVRGJO6kNKsU9uVnwWM8of/TnEHzP3hohYONa3UnzsH6EnmJnXM3Ee/MRPmYtWCZrOjn/
KMHTaKAqoQQw5Ydu5RpjSNBgt4RTtojtYuzjIjM0BOt2NPqo3O0U0DIraX/jEN4ogJ5pYhOSU0uf
b9hfLbtiwWb1jar02gHCcX9Pnx1J8cMvJbeqQDUoSEO4AlRg7NPCl7a6Bblgu4gajGrx1FvMSPvX
DGiDwfoXeIbZdzxN0WQbUvdzBlYpXGcwNE+Nec5Zr9aSS19SOhagMEzhpc2924PbIwZjbBG7osUg
3fRgLHVkaE4mJBTznBPHNL5hN7f5ef/bHhkAbXrUdQsHDGjltiyCXbNp38Ta75BR2U23htm3k/D9
GG+Ns/YpOVWkbNfII7+NeRhvPCAO5rYsAeULZEvmse5oI2A3SXUlhGDlMbeUBsSMIg+xU/6nt5kg
1gRXqo4DpadRFeRvc2II0ZFQWoQrEHHW8daVVREb/KjlQ04wePTHJPIFkCgvzNA1e4wsJ7YwN4Sx
GS7s3wDJQ1nUIt1tcH1WK/GibATObnZD8Ui24O3gFNfyxfhadNgVV4LKS8KWDw61SN1fau769EPn
IBas28CQqDhg8lBR4n04WlyE+0vHUzmORkdSqzG2MNlQ2X27fU7QRxlQDj3eA0x0AjOZt+TkhoTH
kfemxYMe77WSl/FyOkIzaNtC2G1mNtCtpiGTSeOxHoX4Rk4Jks6MBWr+1dT2yqH2oZyn4GNio7vs
adVfWJKy3EaF68YohbLZabjaKixlyMxbYn8rCKrl64Hxx6IokptD44oodZzMnly5ie1OdShQgrv9
SQMfsR5cJiYo6c0A4M4Y7t1QXZG5UEnqTOX/EuxB3EbyyMXx2RRqPiZ15gAxkffUxvY+AOOm4A9k
PbBLIr7nAD2qhJVSCqlMWyIyymJ1x1im75ZeIafpQurWHeJTn+lrKoXgUKNOJ7/pI66PBIQmfa0g
dM0GnU1NyiY+sl6vGEgHdlGGQnCntykRVsHUi+P2r5cMGfhxQyffYA2HQ53lusiUmop3/fjf7Onf
MQF7N8TYTHv+kYb5yHM7Snax56NDtZ9a6ai8FNTEVEf0PLuf/4OJ7fAYu3K5M6q4y7F+U8tk0Gnj
c9I/M3rC3HLBXoXgc/gXxJIdha1jlXdSMTdBLDTaqb7gzAzJTzAwasUaXiGrFP8X9YmODhiJKNik
w903M0WP6I91mP9aR8GphZiXTPE4Q/jFInbssAK4et8gC9DBsbYaYu/r5pChnmSoaYVb7ndzLkMy
WMFxiWDh4Tag41wn0RnKnqViVl1d7fgNnfAVL3AjkRalVU3v4jqyZjEIMG7dXW52yTjpHxqgfu8j
LZDE3tpsYmIT/YoQAZuGySEeDjttGM95M4PrR01iEsNVB91WVmcT66TaOkWWwimHwfOFvVI6UnAA
LY3XLPYv0DvX0+oQyDO24847yqCrsWO2jWPyP6AUO0MgmTHUpFsXDH3HhKmggAI/ao9PEwY3e5Kl
Qmi/SGAgnOeRW92VhNWnAbYwipSsY1x3yOocJ6cTt9qhoMd1plELPOICAIhkdSlMMpLFZ7XgOWan
ruhqfER5+HLrdGepdMIx7fbDVRRTGgalrSyAWTd2e/MbH5qL7mOMCqHymGQA+IYk8t3mkdIuiWZP
tyMroE6ZSsz0KqtP6LVOWYxopSFuLfbJkXtgKqzANTaEHFDc1awoH6A3ZOBhTPxAVCG++5jO1Agi
E7BD8qx69yCbDe4APCWUhZP23yHguApEtoCd2RKM3sdzuiUSFWLXre4HFN1sqHKAdlrpZwFYA7wH
r+4WLVufL/EUiluiW3WNJ0dkWthGt+PuzgJ1mCVfaYMqhfuGGNZW3vXAYWUrjtDzBZHbkG76FkfI
AjReKZDdfCifpdPNbrRroWOYDonodKSGQRXo5prJkUnoy4Xt8RkzOv/Sm3ffcIoYcLj96d7CuBOQ
Kq+dicfPwCR+JQLllpPmiGBVmrHWZ+Jj3aGUxGuhmuqMkuh+ZtDVD/mTGdSJURcKrDLE34IcMWE3
do6vRZ4W26Ue7AgMr2DE8x4ZwHSzTzcai+ZY6InXSO3IWVLMgbiUwgDwokMMxaWgkOrmjPfYDhOF
zmBsgwVEldNC1i/6n420+Yyol2cXqtaBxrUqnfGpYsXVZsujNy/LenoI4PlvWVmJZgyZTlQtuCoU
yAJBJQallysQuq3yGkTiLhiWwQTWTsQz5nOb84IQtcqQSL87Xdqd1oO063B7IYBTPYoa/ZxzzgAP
HsmD6kob65HXStZjfGL2mq+eG2cuE5XUJ4hvK+Nra35k6jTs2px6zpz9K9nphM7Jh39GmUdDhQJU
qFUoRHfjSaskj2UgNFqkde0xb+rLYh8ZyiBPoy8qyQtjKepJNR8ksN+0UJ266BjX8tK8SE9/gqcO
f4bryaBL5gb0zh9rmx2QLlCEmGOHn6l0HRBldzpQgEGFwLnG5TC99x6GUQYCzFyc/zves5fXrF0z
aqeLZq0u9R6gDi+bymRXFZOZ5X2amqBS68IuwNHO/ZmE3gu9jOxftpiMWj/JoK4GEcRvgC1OMWOr
QHFdlkOkXG7DScZIWpf7etpdBECyl2a6zIU8rqTuNdgofbBjBcBrpS3OwBkXy4SbaPRAMtXtGN7A
GAqGhwBcxIMWbSxofsPFlSZKZmxKUUVcJSqLTzMnHBv5WwHyOOfW4+5KP7DexIhekgmPLskKmcrJ
eVoYgDOy/b33tTUFVovxjPNEGdThRa7giqjLrIdaQ4KYB5fXuFrCpoLqsWww7rkREkrPkQk8lVq9
zpPtHgsa0/6UnYRPq2IfTv4Q0l5OB6DVxzSq/AhBLZoc2dh/j18R2A4LUek8s/k/y67tJPcdeuyZ
WDlaiEyCqBRCY/t9EBJBHQqmYYj6s0JYqM+ZqCtpqQz12tSv4u75HDoRkuKlU3AoVbhorU/FJ3x/
EfTr9wH5iJxbyD1cazZDOiSp6VYpUqJMrXPvkOaWqw1zIzPikOtG3yXwXBrvp9OOI6wwn4EU4Tgg
21rhnrg2OsPdPnVmIP7ktfcTu0iomn1PvMQ29V8FwfySBLNXLLnuERjQggQw20s+mn1ZM1R0OePZ
hVm9rK2x2Q1dYa0uODh62/xyMSaaP7TYRErU5jqSHdypN7A4woXeUCKwflrIXE4Tr6Rw/RqoKnxb
pEB31EATqPzYKtjR1v9wuZbYdvt8CR0EbGXGAnYZhqU/IuezZWhGHmdbLegR3x7AlfKwP5MAv8Bk
VD83CoWZFHW8mHSBXK4DlUliE+GXykXBFAHvN7adXW76sS3sHpRB6GDmrIbXkD8qbKTjuPN/jFzY
EJiFmG3S8NVuR44q/N4qKHkDOkjVZQm3nyD9Gh++3E2avAQOvNuC5Iui/z4S67RrjQf7RDbXXUko
ZjpzSVubB+SKqvBaRMJ8ZcYZHLuqg85C774Y87pUFMMJSk87COmEs38JrvUJZWOmS+YG/w8elAfW
qhf5b5esgQKdfq8ihUaHLoxCz7MDUtTE6YKQ1DnM0rJ2B+HSzzRZq0h8Rpw5ARI8dcJQgRWH5O/U
3PJp5g0Ls4gPsArH2yRucauN/bm6UrVzBcbchx86gfsGgOiAa+ytmVbwDSZwYY98jETRH87oskxC
AxniB7FtQD6jEvgDCnq8WysjrAPU4Dnq2h1jTZP9DpK/M+O1/dpNklMsntIBiXmjh8bZ9yPoRhH3
HelLB7T7jdiYV1X41+zoVKOmMc8w0WWQwi0kRpe3fAqjHsTqDpsjofN2Yajg9EITqZPXHDSgI0e5
btAOX+JxcpdoAVo5c+z+yMLJpN4BVtCEU8w/5fXqgNpbi6NQxDVBHuz8exVGUKIfiYCk0LEg0CbK
zim7jN3NevTLabFaQa4g2CC36dIOOrKpETJ+bHrVxajVYTUMpSA44x2iDLPwYp7vAIceCKZuSRsu
OHVnTHXSxsF4O3JVPGCvX4UCAQ9M0XRe9qiwgViUXxBewvdeQsnLFsdAHLrODC10wmbJxsfj71bx
fNRUySDNen2asPB58tNnyvSktDM09MX1j3vpBj1jeTZFooLh2UnbLKACWISavVEZaDwG7p/HuiHA
cJBWl3I2CxLEDEP0ifMcWNfznoRRknxylIe8X2UXMGLOZACXTAFevMwAqwUdNUbvC+5qSI1EinW3
naC9x2ZHtRCh/jtu2UPCA7NWBkswYzNt2rImRUNGv/pARObcIQqOHCd7H0FjODgZ3e8QNBwXcUcj
bufGQd6/kwGDgwDdQHTXHu4ZWycIIfq1GnJuaR6lJlSvw+gHGIArkR39mcQuo15kaH1gbduXeRzf
4c06WqIVCY16BAUhszj0jcuS/yvmy2jlZrGOYGYGSFEOHrUR9S9VExr0MuPaWaYKh3Y0e5uHtl+Q
FpnUpvtB3FehLqRhyPxd6ZABy5eInWnIb61iiLLulnCd/Q/6FntZIolU3pQWqdYCDE1H734ImFAG
rqgAysec+Ni0Mj7K7CtVQTy/3IcDX74fAlhRg1FWq2Errmvs28zNDGKGApfpiBa+sXQlB+9eZ0mX
sU91LvSQJcbv7T8sGdce99lSLJWavsonfur+BNEhbS832g5M3wIVQR8h2OfPTI5DrNW7orZeGEXQ
HssprpuYDEy9omOUnsGQcmi+vhi4Ay4lK59YCgt9yEVLvhGfRXe3NMRngv193jyOKv+4tmdSMoN3
PKelAMElhlsiwSRVM9X5jDlLIilWvU8dHr8rYRC/IuP1aQv5FLpvbkiJfHA8busrz2zNAaU+iLDa
Apjhv/c9Osdxo97EBvNOosjAH+724p+O+tyGZcWiHVvYwCtBw+hS0ZJPBbvfr5L+ydCTYP9uswLw
D1V7BgMZz0oZ4LQ/NKfNHMSzL6QN9ehNs2NE+KsV2AFi2cyF8Sp+E5eEoBRu7uWYN70idBcAlKXH
0CBSb7EUug9BckLiWclYiRpkVC3SEqT23s8d2ngN6UM+TnV5avmbr9SgJllw6/eERY0aDXfBYoTf
Vy7gMjjxZ8odVCZzRJML/qpqwYLL4aKwh/p3x4wxcynfHLhL06k7aFjArjhnNdYS9rBLtdbrGUY0
DsM2mRYKaRzniVluOjOFNZ4H+HzmApyAcuhNmmqYYUsvLq826nKDUv/pJpA+9e/t+lSIu7fmRc12
dCb/UHcTIhU0eUiaFAPTufHnJd7fXX2DvmYz+OVEHF/Nz8jpfubiDlqxMmdhTsNoFynVcMljb/sf
1z2dSdDiT+rb3MvjUv63km83aPrX1NJ2X6eaoJXNeJklixq3PrS0uK64KmmckB3HH1/Mn8ybAOjf
1mOaebdeWHunEu82+sTyU+MZDjJxYZeryKZqhApqFHJ0nrbVJX+gDzDRqJCwgoUbwoC+1sI892H1
RerOcDJp5Igbj0NClNkZoK0JXElm1olc8dyhg6RDpnKvvzkPbUqBMAXZJ3GyA8CpUfxm2utSU4+o
NeLIfGG+F/wmONla+z/Iny+sKs8FjJztnpdoGccLooG63LVNaFcvYRRhTent2a9ievMbYDQoaHem
WDuI8jILeUaQMJH9FQLNXL8zJtNLzyEKyuQSi42AC1N6mDKEHxUmZ+02CfQLpR2qCgg02gV0lx/3
WtJPKUXEn5subYmLq5LazaqqeIRQeekn6suymn9PVYTbEfH65UrAediRd634SG0GgKLbpY4hAGBx
rb7CBkAjkXeN4+vvyxLUpADD7wkAMNb4dUR2f7iiWhIIS5mZxWRVRxsUJ0Cozd8UwEbBnFE23o9c
h9UGGE8zBU2kawxHBl8zCnqvttE8PZDzNiObMYTM8knFGuyqdRyM/OtZfjxqoDqh9hcEvBGubqpQ
dqGDzXYeQQ+4ZVlWhC5Kg7p/pc9xHOS9cpTC3brap8XkqaWDZVmjL5fjZvDqt9NEZPC0mK81Alhr
kUJdGnNHkts+XXAI4bw1n0gSbLWPE39HEklXE8j0T61ChPkiOtEqiTKzpaFzbbTBUdK1o4aIWnh4
/6Yt/uTIyUVlYazXLwNNPhHml26A8XzEWiXD7ezyxJB+if6MHhwF8sEaGVW6Ez2XQSMpT4UdUWGu
TmkbMJbcL72IpM6tbwNPmYj/yEwdUJjeO8ySuQ2a+qHzmJ/PHv8nNWpH4bTrmYA7Vg0BfUhhZWL4
JKLiJiB9Yn9X2dJcZNZW9tQUg9YFHu14b5eee3RjLOQWIE8SC8DUcJ+JWjZohB2BKbA4nituGXei
utZtDyOb4CEhcN7HSZZaIoC3oP1bhGODqJQ4o3sobnxGgC/a7eRqEwX9oDrJiNUCRda57hSPC7UO
Sqpv3Ms3m6HLm5tLR9LAS5SD52JG9Q2HfuIIiuwH7MBrbhN5uKZUJd/w8XNolin7r25Yx780xLUs
ppJac6+zgV8MoU6ryFvboDQraLb94Cb3zCtltVanazykjtPKyW7L8FHzDBD8WhfutBb221jc3zgt
4VFU6yWQVtx+kUx8IGIewqvaMPX4ra5J/JaexDKuxEk7j2GhNA9qJdym1Ns5TFCat8lmbyrAewZ2
dgmJZUTNk6vR2xP/V6RC99pg9/kBU4grkKFDlfXwlU0Ls1htk2VLcbxtNemH2+8kzlqSTzZkkZ99
kfbTRVBn3cyY58c9rw1Kd4MP1CnzObd5W+CkT4ixt5hZRIWvS7X9n4dP4SuTpPlGetqfOG7RdmnG
aPNDapSs8C0WzHB38+EHOZ585VZ58wbo6e3sF7KszgqsuCqL2BXrmq1tOGXCOKDa7hanxQ/yqXf3
G1paeUqIERmd6JaxvDSF3XafEgAG9CX1m2pABeLrG9UE090+z3by2eKoURR3UhFKK30IWVci5za9
z4Ri2KfdziVBgawBPgiK3aWJQjRJxca8ybkX7S8A8iieHZhjEp9I2kWJMWvf8MtjbAAYt3YtO9XZ
G521Sa/lEYXATpMC3cstPplxZXI+Dojk6mPWKb0WsaG/QQPmshFayjIdrEqI2nqoSbBOv9bF8YfB
rm/2ONZyIQHCeX2K/T+U3Mhc4SmXMcet/Lr7SlCaqA7NaXdxeMZF/mFcS9PfnKhihzauUNXfCxWe
zExbzr6HTF69MIEGFyF05sIJaeZ031dg1kYGqNOiAln6DUqireqxywJTEJTlkxFsGlpNI5Y09Y1D
Q8wmujdi3l4REaqUk2z3l3GMwgAzLuulc9Ifo1gyqejMUPgSSiaH65tL0NxSy8j3fHO/jHcauQnj
shSMJOM6jTUZkNiJi1Ya8Hnpv64Z75AwW69waJYrWuKLPkCVBz6xAAhoSslBCh6ep+IT0MfEGrji
hAfzyPxcO/IJ1TjpPrP9rjJWuaHw5jWeKFoR4Bs2QS0Xv8M5PvQ0hN46ub0gncWScCReztWmXgq0
J9oVs4dUWq+a64UkL/MbEhwCuHgPu9iOqxicedBGZzNSlut48FJwhGMtO8OOpMyv59i1E1Aera+B
eYhIs2K+KHZo0NSJqudK1gQ4X4tDyKBToPPzRMDYQfZow3KAud9BRF/DVcWd6EziiB8oe/4SskxW
jQvW4CwhHq1Jnzrhj5n/D84KkZcFyVs0oliUsYgkrGIlLN152IFFMfv5F3obRyaUX0zBtthkcUGJ
JOioKkGnbFbWjRbfC20IaHjJJAADLQ1zuJZN024x2cczTFJlOh20uGNpDWvvhbKYl4t3EnSEbD5z
G7uspvq5KcPDLY1Noha8qwyWUBkwzNJY671kRiKZXKiboJUkioUK0JmisQVODQQVCYB5yUSsHJJ8
Sgs0XPOarvjSbzJexljmOMpsq0rQ1RdxWUcyTj3EAySkTmRQOf0JKLQFS4FYy1Q6l+uRNSzMUUOo
CZMQe6HvS85sTqOr52DF8Bs8ifCRrPC5J02Dj4hcF0qR8g+0ida/xbSnbu4xs96rr9KPMc9+De61
lbcIVDscaV1xwdsPfpVuyIfIUaDH4cTcJtAZTGSikBmW/+acxGQ3j2xfM7C94CFbFZSO7qqkdXwq
65XmSnh46QPUrKmWdCMreL6PnnYiH9n+5Yf/s4BltKa0Er2Uo9VW91tOPCWl0OtNT/l/KaIFNkQs
6MmuGoos9OA1TSsE7Iozkwshc0hwUbWE3cPDPdQA1Pjtj7sfLqglzlAnTzcsuVo05g14yBc8yBai
axAXXUZWewn8su7ki7TmeMtTVzhWqX/Bcei67FA/cBLjYYqGnYt02Y1L1/7E5MSK2Yukn6zlaHYy
yNogZhs1zQB1ABwU0FbtGD6SasvjhBIqeWmorgylsFj/dbwu0BQPFUMhI7B9IKUlTCu9wnvXUM1J
67gCfbhRKP8AVRiXyPYtak/xEl+FnPS5eNXQCCSHaL1lkT262Gv+KhOlTyI7UXGYW1vVXniecflq
lkaa5Sg1e5JU+NmXS8JwJ6gA0xAN8Eg9p1WiUmEeEq0lKv+MPANBsW1fePqkrq0xhJsLsgRyGtz2
Gj2WjIst03neQlj7DBCFzDoCupZd/LzTVZ2hy6WQaSFXIA3xVUJxzM2PwG9U4E4NbNS+4sFRKdG5
h0AarH60XX9XoRTnonWD5BM2nYaXss6gkybviWMyuWed/Z0Y0kR82+MZw+wGxb8pwA7oUTMWqLRD
xuIBv+GmH2n3wpUpoGeHeIlaE5nJVM4Otw4oGTzhokNPFirbtht8wnSYyAonWSe2h8dPUMeHIIqP
yP9Axe2czlTU9IhjJIU0joYDfMC94GUj0UVwp1UKZ3D2sxgDvxv/nsss5nJoPb2mFv8hwSbxayQs
avt2TK++HcHNZArbfOmfjnyNJ0/Wo+0P26CrK9SEedRUoBUS0PHhfnK1F8sHwg3Jjp1GsERqJcAJ
7WLJDUg7AX+FKlQ7Yd7hHOFZUn2zkOSqvHUcWGeFGlLqqVaiTI9+VjlGtn+Kcn+zdpZiCIyyKk7q
Hjqv4pAWpprELc2Rk4o1SsJ7aQUO8Ty5IdddLhQn32dob+yKrAU1qeQcNMP8YcXBs6Mwwyto8Tj5
Mpz3TPvEIS098N5kqqJimB01aTGzIuIupm2cZLOESFpCNimkTF01mjZd4gstp1fpkhNxYp7B0CVB
Iz0xedAEjheOShnb9jhNSfGHhW+R7duovZkCG4cjmMpKmEk3joc5D5rXnCLJFVVR9//DhGDiDcWX
g5xH5E2JE3BVdxFnsGzGyXefDaPQEUbOM0pGZREGhbfh9CUnDQTvPFE0ji7IzQwkgLBzrJas1yZC
W0woxz35vcvS+PCSx/8w7Z6bc2LAyz6e4gtEeumNK6X8RaoTW1BttOQsNNkz4gcVlzjGeedL9ogR
tVdMsLlSnVJ1JUsfHr1p1IBYc7fqlnJYfMCJQDuMRZfpk0BSTLYXkJk7cC+0xcjvDv+Kt9k0IYOa
9nUx1KxRhvGXez6LJBdLjFJ0u1pidFrcD7AR3r2HLqPdgIotbHZQXuZVZ/hEPVdDQETb5EFZbFBn
nCvSL8gVV+NO3mDOhgFFHB/PnohX+Q03o9OMvrM60LkwyJ3tIHyxiwPtCJAbGrkR7LQz3HpHyx6f
V2gOhRI3roQgy6BkhMEBP2NcWiBUwyqh8U2wYH4TEAMXgGEjR7rbLxrUFUi5tVgv7H+qw8Zg7jV1
pqgQaC1CJ2Z1ijjPWfFSkywJLyvtZc5oplEm6i58qxBk43SPSs4I9zIYQeQ3K5Lygao7fKcMjTwL
j7b8LscR5MWyEG5y7aZQB8fP6HN/c0Yj21PpyfbDEB4OUvuQRrGslDtlfZtpG3ckFwLO+prYl6w2
yDI7c/hA+Hs2NCaqlwkeHfoMofEBRE/iAAH0t9lT0U7M4MJJH+3A9PWg9mczn4CqAK+q0Kno/u+W
flN+QPV19D7jbQKnUupf+J3lvh/5lg4DnkWHX7N1YTue7KJ7auGYn39j1PM4S9ia48mS1sjKX/tv
qe3TkzppS9oqpzMf4Nx1huLTEJ8ppu6zwNH2iuFTkLpc4jksVzp0cHNFMxv7LK16vdNVuYWU3Fyg
pxKOU7LlppaoA7Q64f4pMij4ySPIHZXT5VGMZh9mGu5m3f1Tez60Kz+S5j6WdTBfImw8OBjzQjaX
fywVQSM5zcIe9qf5KmLhNBTasbF3KLSKyEvLLIJlgGKddrmLAX6Ggt/0PJ0ox9DU1MoebtRwhVRz
gh3uWnn8t8419FObD3Np2q51hnSJ7IzepDJTdcuNrxd38wuXkG77EHv94YsH79vMtsrvmwpTrsbj
QcHd3AwynHQ2qBCYc8X7UDJ2BdN/b74/4zWNO0Rwo1K8x8tz+5j2rMMnIPqqx4tvnSFQm8fa8pPv
JpYEtSlIjh+o4YvMxRdfH5F+8q7nLA1H+pyVflUJwyS1o7FZbZuPlSgaO/OGeCrE7HMxFy1tOWUF
HqZuakABi4JGToR1PyXyxemQy6038ANTmF/XJAGYzwpOQLHJdnK3JGdvGVplB3xGzqiDVRJVhhrm
7nBn8XxTLfLE9jNOrJdux4Y8Xh8pDx97pKWCUMhF7WqgZNtIOjIYSCmHm9khE8IXuDq/yoMgKr1D
MIgL4pYXwNb9D6/PHV3x1EQ1LufZBlRfoW6nOdNF6fNEbcbcGElTv8x9X7nu8Abr9WrDHq4c9Rpg
5lTXjFVK9k+0G3fw5xKpnttANWqp6IrEVUoCf/844fPKL+nFe4fx60lqMcju1lgDFGWYce7beXqd
VLJK+fG+rn7jSG6lpmYNVSvutDFC4LK1ZdikTzpEFFL2YAQ9PNYWTaVBPIzuN7yUgwBkWqTOoqxq
cCg8A68ssWAjH1ZykocaeQcUg2DtH8utkoLgYpHNdHFklfglxB6jI/OqW3V3ux+hEvnb6G0o/o64
l7svC5aC8lv7QFqD0aukAbe8JmexUnx5g4J6iyG71dTBAmiTJna2s+fzAPSnZ/SrsjpwJ84oLNvM
NSvqSrp+VIzvxtln6NMo3ttc+xPlErs3WWMvLtL5lRysE7ZpCAHciHTHgRY9lr6iYu9Qa2qHkmFr
xRudG2L30rPqPpMtu4Kgijc4jVCTFRd6vLY6YSt9EQzh/UKLuE70hVPFc5ezBpDfdLXXPAzmDZUl
p0JKpfGk/By78ZCSY/bBO4LlBkJjLKx2D1+pRGanRKkAvtDxB2kVm5MsmQEjp0H2N/bvsjE5jBT6
yt4rjw+5CjnsxlVs/EMpoIyeyv2q2SABptOzIxh1NWziBbL9xck1w7ehJENOLNXgcIMIkpd35LqI
I2CrgaOQ7vkjGP9GcD3YjFcZfnsKdYVTo8Av0kd6SmHmvP24OvRSZomGlXZkdYINmfW6+QO9XPXf
7RZBt7VussNYXNpF3CbIge8ZkwlBmW0+TqkKife4FkkhARyJ2lvs4sfaNUAhURSyhJOAoEyCmVIy
dhZgWtwQi+rFHIrtMYwTa75VyH1ltfCUOhV2WqfA2JSOYSzLLDjDfLwhEuV7/zFG5OTbhpciAHs4
XspbIBtanmakbWml1V0qA5u+9UhTh043b4MSD3Nsuo6S9zR9bY5x71O7eExiNuTMpuFSwq1R8tkO
gBTAMLlI2YF98Pzgi3UiH2RRUj6u9DupVACCQfsxLhwRNv9cayjlQsoEW9zUOmG85ciNrCP9S7s2
a1UikezuCEO3cBlkqLEzvaODPuEdIC4muCjlmfURGGmeGsnRCvP43CXilc69Wp7sHccNPTT/JkX2
2WjpJe94ow3b7KRJ0pMeEc8LNAwErIZ1OYflkTBntZFJdnsx9LtJZLOXkWg04G5jhq9nJtsjYnQr
rlV4Pku+EGKG02ekDrJn3/qcLKb0J65SkLLaksgUa2w7OyZLBVyFGBnEu1anHQ0qIfY255NLTX0L
UW3gCADo2VsIS89pO+dMc65WkYUGjkNcBrArPp1Ir94Crlma6caZEQDkqttinTWSkK1wNuwT5aiI
SJ9n2zpedD2rCrDjah2/n/Aj0uxbNlI3I/wKAU1+vryio/SWws7drkfhUH32dK4cP6yIub+cbLdT
k3XptPJicT7sF0pA2JDjc7sJsK1DMFu2bVqOhST9sVVxLsZfy/9i2jqcWh/APYBUOOvV5vLKqte9
ZWG0nCTKllo6w9/mfbFPIEH52DLv/axSAnx9tj9A/XFYHc68Ztxd1xG1yyoB1p+stH/NtcpHtp6Q
KGPbyedAf7oGiQPHAdjAUOsXTVy04AOBN2YeSCSmoGLXe0L9HDRm/0wt2OBJbnWVwac3VuyB3mCg
rYH4LfT3vpfCjoESY6WdWJUjNiTYvpWzzVuYQN3wwQacMl90ioSzCuqiTNlg21NkOSgLfMdFay/g
TwfOBOGH7UZguYJ1JvdDqtiZKXlqNOBkXCd9vEKeOrbu0tS+LhJXC/iMTqsIGX+o02PPOx+EQ9vW
KG75eMQURS39x1w0O8m0BNWvWagrB2Z8IrDKIFNSyC+1gHr80eW/4zqknFlWd1ABor8c0/A5/ja6
82FGaWDWZ2u5346YF1jyjCFpMTgdOul4vhhiEzSv8FLaql6xkEb95dilinFUYekclvpxzV82hHTt
d3AnDKUHAkZXy6JvgqALZ+z5t86vznOEJIgd4rtlWYEdfOyhABrY3sT0UxqUHIvENYjc5xWBu+aq
NX2tHduOjCJHIxrLdBj7xPs62zzH1xzvgWzbP49AaS8t+k5SADc1meUH4JHFGwG/mPulUiwXuvdu
639U97jL9Xt1lfUrXMDt6jjqv+x/Tlcq+uchuF3tqujZ97gDBY5H8ZhqXqVsw9tUEoGOyBtFRgoB
2QthG6larfl/OSEVodfaZ7y/L7TOYEHmODqof7dZ5sRTpqbvgJAA769k6YVKSlP+C4AzZSucuMdC
mlPmFisTZD4u2db8rqc/tZleZiDIyWS8P5b2E+LtwxYsP+922RAJccGA2umagNhRnwmQWkJffk4Y
HXJLMAluDbncBlobS4UMfN353X7OMLC5sTzOuNM7bLyQasB9nOYITRYxhHMWObNCdycAvKNN00Iu
w0bqdq7b0AUCCY01EefzKsURl16hb0uyS4lt3rzNvMlqfjcG1dBSTZrqbbfRxgcS8K74PMI0f9Vq
pHSfQI9v2sYvdGo7qec4LxEbw2e/mJEEFx662or1tr7Hl65rtZkM5Gj+7r0BceGc+1F/BvNECIT9
OxhHSCuZoFL9szMSkkfOytp/Hc1gXd71uKewBWbMuewF/djNDja5nKj+aa+wVAN2TYwEElQTR3Zs
aZhntWkcVEPQjZcj5P+trKPeeMpWwlzbZa7+A20o1RTFCD6FSXlEwBvhrKRlrZru84UGFttAJgko
ZQnmE/9PzrxQpfaSDwEGKtOvJK6woI5x0Ct84oLjl2XsKgddQtwTX85Dv1QZlw7OYW3cuiv+4uhi
l0ARKFytwc07Mcr+cjevKy07rnYbmaakvW7d/YGOFUIULuz8tSwJ+TRkcu+WQrW8LVFq/sd8UQKP
n6iFUPBS1Ii0o9Bu+Wamqb5IYL6a9ZJl8pWFYOh/3lau1bT4T/3ZvVf6MLSYDz4bLuoMxe7GE6I/
tEZHCdTEBhNpzdtc0SdDEe23yRAnkl6HS9rM80kHiB53oGbRN5G9c6iR1zM3HYqQhOIWwQojQ8MD
NDcz2cKJth4+veLnKnL1jQYXnDtsEM+UfzgJ+Iuwl2sPZmEPiUjqb019Q/35sKUdQQBN+Etdv7Qp
ho7wCmZsWVjVDLS6CGeYIsE/fY0d1E67fVg4pBvBhkWvLkID603kZl2ZqMH1w87FBtzgl90+pVAl
ZLDjsPjRFQAIYvTLfMfHuibb9l8VJWM9RMTFX8vr15NuM+0fzQPsmbPpU6HxTqk/ItTNmCSb1p3/
8nDBwi84ww6oM8rSCLBeKXNnqQYBBUmjyLMzXGehTvjfcqHncYwML6j1moynzSdcWEs1rcCfyh6g
IchPndypB7zxOBpM21ZSY7GT6Q0cBsGyIRMekseKbGXBxvSYfWMxE/vTaWG/7A123RN+/C6KJum2
JRTMpbtTAF24ZwlvHkNPQyHIHW1pTd3ox/f78LjF5O5HLEdohJSWMk6XKrFCaCHLwmHR68u93DML
bMwCho63VcB91eEFu3VelMRKK8G+wGISP1smEJv2ToWzdcknSeXbrtThyvHm2oQu1BbadvC7zBSw
bofL/Xj++bhSyiWeaBYC2DrXXLFp4djMh6m7ZFTMx/CG52on4vdbD7iyZuOlOC6iayzxJ0ELv9Kt
XJlHI9jBhjLzo5dLd3rAOtcZCZHgvpZ/yD8Z8CL9yk5LpGbxx1XbkzKbcO8acFoh5bmbVrTKcZFD
zJLACu5PCItjudMJO0vRCoK+Osfg/+R/sjbyP8/E4fqoWBUIiOQknbqR2jvFnnoqlhnmA1R90OtU
zuViKnQ3E2c0isdPWjJpvTxZdWnfPcxuYjj0DbhoRZLfg1FSrzmZoatwMHHOwcL6KXErRz0YGkB/
qGnFH6hDlPzKSf4TL7sVU1ujNQjUgddClDJwqd6ACViTCiz8ntl5Itn5T203RgXmaa+MA8M9RKx+
897y5iU9tXWfNoFU7qVvN9ivqsHVObDINKqnuyKd8THU09tmQkNtkOMA8zxUfAGhOSQeSxTIfxev
qTfDI4BEN9k5ZsKHrRQx8mizf3MDYD6CxihQQcORuy1CISEtcrtXWIXan1C7yDrY1LbmWUSCRsnn
j59peh0/g468pjOXVWsc8cwX3Ch6IgCXCyKewCakTiBwjuyMm7cUXRB7GT0CYA666UtkFiIJ3Gff
YlBOGTaZRjDs04YYEaF0OGdYrDFGsTN6BexhZ3Iv9YHpDdwR9RVHeBI3zos5YiAE+paAwi5yqVWx
PK5IqwAuu/5y+6yrnrbwRGbWVMmY6wpQRLWrS7Xt8AJ6yakHzbt9J8enZItffAQaoWizl6C22nTg
wRI/1tKntKxQYiDzSkVvSS8JUU7j/OR3/JxaV8aOeUUtQcvbzE4/3rXNy1wINc/WVco699+JOwq/
RfbKlVqg9RroSe88t+ZaUXhb8HPDQjo38WEvpQ6ez3z5BI4NvKjFc7M3o8kf/9WFfeOI8Ps5CD/i
OH+zuVCLmt05Non6dGeUb+tqF0HvcsjyBMr1VXMsNQl7F7qgswiPEMsE+iBwIXHg56X9iw/Uo+B6
5ax/YMq5C6lBk0AHTmPdSAALg8RBAMjfMZQKHdc4zFOjBIiIK4FEjvH4C6GtqqpW1VFInKAwwD3v
ADoUMJxFbzBgcxoSVnViH4HJ1OWI6UA9HmQrW/2E+XmU4sBN3He/IdQAy5DDLfn9W0VlaTMmBs/G
eXuQd+rRyBkIezD+Mfww0CfEHQMVjI44qKBH4Mjp6Q2dX8MKvY+dVf2w3Z/aw5v2CHnekILF99+k
3f51Ikx2Y5xBKSQZeWNX9A0Q74+PlsY38K0q7arSe0ffJ8I4YlubkflOUAiFT1voHRCH1okuE3fH
++Ivysn6TEBCFFEBggcLVXVl2nfs/gpd8lOhmDnggER5lBHql3XeoQX5hPLAi+QXClxwVwMEod/G
kYNed2KczUCmI3lDGOq/FfMmqE0MXr4dC2aWBeJG5BADgj8njjQvksYpMwpofA7+TN7aSZa0oOoF
W+jUwTyiFbruDhXHVOFs7Pg0v5BcOL8CuCZ/FjTc50w7WrmHmC3RNJJUYn7zzG18IYOMyRl9CbMv
QsT8wYilA01yEXAVh69qii/MEYRq0QtvYGzspx4+TJIjr83sVtcjnFrtA2y2ux5SgP35W/UZPP7z
1kyi1Em8ZOpwhJKk33tWmywVH1KUH6dRUDSJQbhl03cErCbMFlBsTB72xAIcd+0ePVccQT71jABy
/xH84nP9vakg4YIb0G5a7+yRBbA4sqVJRgbmTPYAM2xWFp5R6eF5D+YT2Iqz6vYq5/IAvigW6r6X
WlnTUDiWHT8DN0HhLN5ueyy5NkGpL7mHxNVs+LAUbWo9K2d9FzxfmNsDmAm8mjumdlIpZlAiqBu8
nnVdw49l+A/GFF/x+PKU2DZFQpUF90bwlnKYcZFg4HZmaV978rny9SHQwr4tBazD0d6Al8HOAWjZ
XEd4H2fWdKifdpdijUYYcaWS7996MYu1P+Vi2yjZ655O8Par+Tx4AG3g2Pb+ZtwnFK3Mlb+tp/jV
+lMxGEBAuQtj0GzQAqZE75hOhRTUcK4scgaCCennUnBqUXN9JtVLWobNYr+U7CWX5emy2XER2YGo
PfIu4bEkDVHC+K/YpE23yZDI85fctvmZ7GnQKOs//tzTKdEg2lSZamdJCrBx3D9LSlWz/4EltiNN
NkjDHpJEML5ZRuF/wrkVahrPSOzOJdCs8lQdiIN7qoyeYisEW4QnGZ1GFIVHbRAajbyWe5Z5R3ET
t+AWD0v1UE0LOELVv/JF5/d0Cuco+JvU/xqXutM8zYioJ/1TuvzOzGlyEHCvkBqynDqpyHJb7ZM+
ycena1KskO1I1YjtdC7jLWcE7UOB7DU8VyK3SKD4v5ZoT9s9ARemMwkoHTdNp/wfBCPg6A6GxXfH
nddAFNz1OUayLKDcO34Dfspm9L7TaLTrY9KZ5Xtwkfu6PYRceOd4G3f18k6SN2FPAEGDatUkB402
8bMr2zX+k2wBjg5qrP9hUbfXsqFKnN16hfs/5Vkdilerj+m58G4xADh3ni9nOXjKJsUYpxe8zGyH
Gq34yL3mlnQzIz9PP4FzbtuDU8AREv8wM4Kr8YOLoiJlEzhbvsPq9lLgsldaXUxVHuBbysmvE21O
Z7ViPnMHbiEKzDnv/qoh+h2tfdIv2KgHQejax029VnazrfoEZEIFk3PUUmCpMv+7TJI8gDbnMlQR
TUBTp2MyPz5eVU9Qd3xVUOsVKkpv40HUcZa2IToIuwb08OGAL48CShozD+7Nrag5N8u+BG5nIuPR
MLF1Jxeury06uT7IRlG3pyItE+H9pViHCzrj9ZJqH5lKtzf9iCpbpbf7PzwvzEtlpaN04cbaizTx
Ni08qYPrl4Ao/Z7jeJ7nIOandCGnsBLo5zjbDV2tu7zyq08Xd20YQ7PkihQgw0dVnB7m8n3aXm/5
SwENeiG7ov2dvyvj1+BxiMuBNsc2+fO7QfXprB7QHDOLePvoiGNgEifS1Xwt0QKGk6gFwSv0bf96
LflO4OsOLUasnnGo0Iv44Ch5bh4/R2NMQuJDmC2PPO+Xko2rL7IN+JqbdXjBOFfX/NP4KQSaLa9o
OuKJpgVEZ7nQhImvQ2k6LlgcDDCJ2tPaaHPiAly2Qyo3Rve3Ka1eihLYpcCs0LdCTSlYfUAR7lnM
o4wqsU+0cKBQf4Y7F/tgT/2uUBX6FbEvH/sMx2U271PE7fxuwSo56KhI1z3sJyuSpP/TotRRQy/6
K6qxH9ewGnpT3URHEnmCd53KCDwelIt1GG6ruon0sLUUvAWwJtVtwrEtb6SXkQAx5x4gnsdSpkdy
Gz8AKt9qdf1vd4gwtDIP0w/WNjS7Unins9s4b/mWrsQXlhMcvJcQNDDrYJ3cHrLh9/+9k+vHTS2z
O56o4TJHG4dST3+szC4h6LBByprA4F8o/0ryWq5XY20OVR+gGSieLQAiibfFuHrlI5a/1vk28rGF
1/OvEbD8mIxcQZj6XlOgvhNSbCY1G1liC2tCfq+IaJ0wVn+rZ+E+1dTlzrpiQ9YyIxqqZnEQiwLC
FIidp3jyWODsf0iUPrzmCG7m89tfbSI+R/8oiDFtCnQqa0SatimceA9h5vXz6xfVa2h20i+1vw9Q
Gu8Wz/99xG+xb2kat7W37N8wARomQMUA9BA4l7dq5f6lZm/vIv2jG3rj54ZZwvkSTkSgI6LbZLEV
LzsJsMIphWWlKAJXCnpTug4xzsWdCMMn5fQRr3zijcwqaUcjQzoKR1UDjWmfYXuTKLE3fBaHEO1v
Ry4SSVSusuXk5P9PlWC1PcsGTkw+NjooelYVYslAjHrmrp7cG8pgBlEiwh0ix8tpzvEEdSXb1Is9
Qz28E+keT6ZCxU0PRioUAwPdSYX9b8iqGOLzRdMp9QZe+gFEExyiGpa3VVwKRGlYMDVc6W0rnYGJ
6zr83TVf+hBO1Qk/NgcMGsHa1CFUuVVl7SV+Wg9M9sYyqiqPqW7CdUAQb+g6KpQQQrkOgg81X31W
mS9clizngfNHJj591X/UF7lr4Uwq842yi2PjjMzoqMZ+GoNNVnmSjNsO+ENS6dK5zp/5CftpuyTM
OV55E9izfC5DyXkUOl6ihHmAcIQMEHDGl2WcQVdgDcCNXSaVss7MQlrO5obSU91n6OXxMIK9A8/j
hRNp8IwbiMFqlVQiV8O7PQStRy7rLb7Xrzl3GUqoYtu8+1DKUjtC/77aO7Mny/S0hSRorxI5IaYv
STJSf8qmIhUZMCnUTOmgqa4x1j7wt+8NEm29FxAQ+zUPlFtgG0LPRW/DgauaugJXeWc7cf739s0b
c0HlllN8ptV7QW+D3OQStZb8FI6vn5nfyPaAhJ8ycxyT1iHloHW41gDPX2KcTsudmIlXnJquTYVt
fz6aPzLGSXH1h98HMBVLJC32zNbtaLRZidEGzlhMgNVQsqj+lfz+aCgVWO90m1kuNYcbo6hUC7vj
pTNxOjTZe3vhx3kX8Nb9nHOpmgCjCM5dh/p5aiNXgihujF5LxlaJVsPmjU47yNVvv2CYd++f2BVh
Ryh9+/zVqUZV5JXXM3OWeHuXGf7un7laYk1BXqf9bcPOk5tu18DWby5sjCFrBFs2i0dfC1pzexOr
8h8TjWeQiVTO0e00r1wNbVNvJrpTGh6+SL1x2JoVpO2SRaGA8z/gHaGB4l8ITa4RjcN5KuYGfHw+
NV7qF1JYvgzYy2JFIlCGC67lDstLMfS/ZhNR3s5+mYZfxpyebYAlwsPsAHPSMVKPeoI9JCnf+z/Q
U36TpO9L04br+VuqouqEY8ra9FtgLMlL9vmbhylP3cyhSGro7QSk8+PrQ2F4SocCf77Ormwl+4mu
Qabq3b9FUwE21iWysdRoBz2Cd8MTSThpqDXzMEEpYwLgmEJHCJ5UGkliOTFpAjPlzM99f7ehM7oD
oxI0v/Au0+iNAPlcFEYTfQkDXuFM48NGBHMMDiZojf82WcqnOrCaEqp3hwpannWJ4YUgwK96DgZj
eoPeulaH7JT7QN7CxXkqa75QRm3976X45uq5bnCx7lXoUiPjlxPBOwh4eKShKfm2RJuKaga0ImEp
3jopVrfwCMa0IqAl7Dq+ZgnMfWoETtdBQXsOh0VJCiU1+0JcgdbHgJ6OtMY4FtBJrKJeqVL1/7hm
flGVd9ivYCyRXfZy4IwYpxVnolaS/8uFB2vH2g6cNc6naKIhqIx89ryR8XQZT8qVUGAW9T/epbGu
BWJyk1mmS6XFHDMrr8dt2cR9erjWZ+7l3W+atZ27Vt/F13cdnMZKeaxtAfwNcR8DjjjjoJBxvOmv
q5ZoxdBM5JuN/pt9aM4xbTFQHHSNbx8Qt16egArjc0yFhmUnYCW/zTiCVTduADuhJB4R/WWMYeoX
6LXf/zET2x49EfJwi+A4tciD/9JMkRcPWIToQkE2D22tZHAaaOSWKoVOImystAmiIn69DuhrTdZK
uWZNnqXT2bNNsvhAsGctDRa27tkPLRYYjvwxJt3Ayre9XL04ZbRHHoDyO6OyI52aGZkm3WRe6Hma
x5H89G8IW8V10KB9AYuEyueE1dyMbWdg1KK/a52dI5UBeG2Q4sryZn4Wm/V0YzgBAqga4mWssYPc
U/Ju7NqVptbgL578tnPruC3mdnrvs9Qw0p0p8D0p4927foruCR1apIHnEXCtpNvvrRaxSXKvVf2c
TU/mE/M3PWbhOjs3cIDRyhAtwvmB1ikSkh5fCO3DLFv70o4kB1irbGlyH2/2DgZ0a0wFUDSKdVgu
oxaZIHZfZic3I0LI2PBcKdi1izsCRcOFUMRtjpBmt2akCVHtlKl9ZaO/Ys4b+UuWLCqN8h/9sOy1
YLNrpTG7asliU/GHJ1Mb+tBI2vypvPbuoSau6TqlaYpcSAPAo1m6MUFSbdrrV3XYpSxTCWKgmUk1
NDo4QFFEHUmyuPO2+d2708g102bI8l33m6UmkKTod+Aw2r1eEuDtPXBRiyoCWlm5IhEzyYykwUTn
RQjNFt238Y2YNIz2nPH26s3wprGVK40lVM0Mbwh6RoE6PaMGj9yIj1n/7x6Lt08aS2rlJLZ/AIKG
960ssxErUOknPlOLi9DLQqAll6ZIbuXDYu2VHEsy9q+uldVUI64QZEXNdS1IEz4laarEDQmpBjoL
YtmvQ1AZoexHgHvcGAIwbv3gPlMcoXCC1sfOTvYngOIBGD0n1vwlBd3DtIIo7FUvp0yS6JBVTebX
4m3WkUbKr1EoavR7n6hk4aTee4Lwpo9C3qYXVexqtneveLnmcmRX/MWyQs/IaT3DJDd7WGXGpyjd
sJhzvwhtsoTlVb1bw21tlX4W49eM1n6yxOifxJd1KGrbt/JuiyWcqJL2TsOjPXZz8/EYGQ3zEvHL
puvqQkg6korJCbW0JtoJO56r5m01KIFfJALYZzx6Kwwyk4LHRmBJRXRhr5Ps022C0yEP9DxTzZhk
LPeyTKkGFjYLkCsBI9FRoyritXHITAwez2+J+ihO4ZL949PQK6WQgsKwaDHIK2lIJyuXZIMW2Lp1
ykUIJp1iFI/RE9hyRAtNh8yE81JyYpO1U6mgx/JuKeSogU5OPK/3lZ6mprr3RF6RPtGaRyVwGRYy
dEJL8YNKGb/a+ptrVAymko3dO7P3lermMf00+Df1TgLPdtV4SdfJSZzGC3yAAJ7Xhjpfbxd1LfRj
vE6pnGRN+/VM4jnHSyNToIzrx9FRVx+1829C0v2gjg9Uy70IqA+eUMnhzPBpYqNm/+xy99zPNpaM
mk/q6tqzOQKf1J5WomdVX7YQry9TYx3Z1fuHLOY4BBA1Z6NKw8AwHYk8un0VMDvenots7iL+Jh9T
dKAKeeq0lzTcuZHsW8kmi1ImixTkN4MEFX23I8r6ETi0u18Jx0TZEfl2p6etNLiwkTugeiwDVfXv
ijlSjWkFppJn3KMhaZOpQiewW2+Turr11QNLeCgNF/eekcuGsasFfubxieLTMJw6eaf/1dyF6D7d
f/qgCWuZJZQiT9SgF/Y/DgGh6yT6LAEPiQMQtDuBxdE8JVAksZQT2Zf9XDJNr9HnKngGVyTNxsPd
eQYi8Qqa6t50H1CVSp7dLtSeaVJKrlxEf1NBnUcUuuyH1g3cX08tH2YxPxwyjHj4ZlDA0HczCpOq
aEwLqSCWbfyAf7zoASFx+VtdDSKMSQHl6jXVmyvSoXARvBZLYAQ/ZvDzRGxWyLVrvPixU9U7jrqe
TitTQUpk1XXt1qlQpNdNGDe6CjbD7tr9sn6PfWYVN7ssKarq0207sLBm3FnIFrItG0V15r/H/WuO
E+atzbZENZazYmNVAR6YMBFFJNX/3LMEM5PHAjH1dOuFaU26jLegOgooMPBEj5mahr+TrUyoi7cn
8ql32noE/rPU1UfItXL76fnbKb++rFTkrs3yCCS8ji1ct2AlMKQKnwOgLw724jwSowCgDSQ1L0Ek
kzu9T3mALlP8anGs/tbOGNdStS4ZslGbpVL7LPLoZWT0cH5bKqrG9b//7lZLI7JeEkIPEgLqlqdb
q6AEm2LTK3kAv5OAW0ds4upz5nAePhUBImg3b2z6zs1Aq4bkSlsW45xxq71r2BRdc5V22Rb+bRMQ
CZojkWwDuWGoO0bZ/E86kR4ODQHEoM1FzLXJ15o+755jVG9tYH+YFxDngL6/rJaPO/l0ZDU8tat0
GzyI76FiB1rznesKAwdJH0uUF7FHdSOKtacqmPF1rNSnIvLxshZFhTUJSoGy/+ekk1lBADbaYrof
LrkdKn+vtoA9AW3Z9SgVvnUggxL/4hp4hy+2TCfG16lomFjAPNCY4ZFyDORYXC4CAgSRfHw5kvN0
D5zUX1lcYaHKzdSyqiFuWB4Sb62hvo9v794fTNF41fH1U+IThsWVgn85dMrTpqpIduh+JGqm5HHv
o0VeK+5GJkkZCNICx3Txtzp3RvLzzbrPpktbTAMB3HAQgZTxW2rFx7MjE+wBE5T+QqBMIIbwhfIQ
+nhbxi3s4+O4oU9xE6lYvm1eG1w1f2lBw3Z9+T5auwFzeRyCp0U+lE0vEAX/Vy7UvQHl6GfqUGFA
KOzLNtJ6N8xDni7NkfgT6HCBDd5LRYBvaMy4o7neqjHbvqsTO3h8kfYSbaXNJwAriR9SqDLbDN9U
l2zAMtXMmMq7yimTQmCUDIVEBNgvgTaw7KFMY8b1x461wl2frJ+5FigNuhm5tbkfz9FVjRqaw5sG
rZIlSjY8ogiz2ap9iW4XNLGfxxeQad57HZjS+nP4esvaH9JNUb5QAwqTPj00xkLuRVsAO8FtSdy8
LlkNvDnbQ6RMkDDmn3nj5XPddB2EG5i3ZDfun7dJaswoz9FKvRLv/VuWz+fxAW5ZBmQpnp+FWpTN
p+zqlo0/mFIu21IdudupXGFYmKZMKxBxy1mF5xL1W+xvCmTejFq4RmiE5cyLxy5DYn8/3mw9/F3v
zM+5WSbf8TeqbETqi5w4UBqJpOZ0RBaWfXYZhjaB0cu2lQPbqxHaa/BGaprJ/E5Q7M3KWuVNOSLK
GfkHaINJcVtC8NXG5BDyWeNRR/Vs0M/5wUEmIsAidHQ4/RBwGKp13gnMsc4Iy2f67V10ggALoYMZ
IoNSPs4lbdMmVu/Fw4ikZyn5JsE7jVx4eufO/e7Dl7MK/7J6QW7kqk7xmmbfeAS9aat06ZcqitQy
KCAcXhnqsb2Nk+nDYFkuVO/S8/PDHuV6LMPJyIXqTct9XrllJ+E8QbHHodS1QhJ9pueLIpLncbY0
yVgzC7XyG82utSa7euYEZ2GnYTsq7AHFNPA0stjRuv6N0OYSBx9H4mkRhrs7iNsHGt5SnNtAV+wo
dC0vP+FYN3/pksuMmfiYaYVtJQdF/P7mTITo4jkBXbrhSS4twfrsfk8SB7KTlwutEU1TCY8PjrKl
BaWa6Pdf1Uh8B7XOh6UcPVlIrxTagmcnfk/DOlJOYtgY3eDszLRgYsuhoYJ9iswGF+QjFnmDnImX
zYPqRdrRpVS6wvFPe2NOr+UTtcOJ5rvK/+U+Y/it0SF4FRaAEJVz4If8fQAWWbu1iIENahyEuO5F
3wmbnIvCV/25DvLNek/QueRM7lewWwesK7HvKYVH+LrXzbv0tJyDjWHPQu0WwjPxmsgSUS258Trw
d8ZfkEU22KDF0P9uaW1GIEDFzIXKQnYweS2HWmXR6QHrY+RBOTWPS+45/ENfj8AV8QsUj2YI2M3c
NBx52UARMPtZ4cY6mv+WQkq0eJgim9rLxD3r97EZQEXkkohYjjangnVitJz97GkfHKkm+5pekpsC
W8upc35DU0Il6t4w4WWxKyhNVEu21GRUJpIxbVS03Y8JpEf16+WAC7enVoJI03q+nsRMJRXqVI4A
2g4YAdvKfLelsnUnxF7WXLeIfqi5vQHpeIWhfzXX6w0eDzyWHGsNuJFgN03QcTduK0zVwy1/ZjoS
uuVmo90mRqYSidpefKv9T6UIswc4EceJU7bXtVUJ25kQVWF8BcQsdQuvInuZW2CNyYxwPx6k6ax1
ByUuHchSUuTBlyTkuSafWPR7Iczstda7nmX5NYppEg9ZRl2rY9gRnXKGN9W/mI20ylJFOSZIV0P3
VkSn3PVylonKH5/xiqE2kPtfMghoQtl/u7xzmnZjzel/K8Arj8scaOAnPDVAkxPREYwNUm+okKg7
cBF5Pm6OXL08F3Iwd62o8WIYZD3vtwc4kUMtwg7o7UwWSjbx8XXSSKecyPhE43UWYhbb59pDsmnn
9EAi/QqrhsnN1kHulXx6o7pginmvjpY5VPQu8V/8qQUtZXmhz+rbIv76D23NeCjuEBuuOQie2yUv
fNFT94iP7Q8MlVm7NS+Lyl08PtsaLpVIQ91CVtgfFWDBdOJvq9NPSoTlg6m+PWTF0i/E5cOP17GU
s/msJ+lj4SRc1RmnQfJGd3v5PZ88RXRZAU+syTgGql2hwXD6pLY/7O9czzk03s00lNqmyH4UnPQC
NpMFVxQp6BzTpi0NJ+AAP7RLKbsNSucYjpshr52jCGxfkcoRgzgBM/3B6NV4yTVvCzzzF9QPSNFH
YxO0x104D25FyOTzmG9qV4Zy1/3NB/SXJAMJhqZ7sk+bpMipq5wWLHMUKEkMXk0WKGbUFzgZw4ZA
2tZQqadTvXd1ZqX7g7JP7s2Epz5P9xjzKBZJ2NbNri2VgNWPXuOtmpIvO40Rlsf9w29KeucFZG5P
z4BGp9feY7c8BjXBdoynmVr5cS1zj9cMhOlH2Au3O0Jn9Hq70dK7DkO5srfmCOOo09Cga+5DpaIA
WrSUwy66Im7+NUVcLvI8HvC8zrbsPEvaHsUbfEQAg45fVeSuSSbrNO2U6J82AiOw9O9HkOEleA8N
LcOToqtcsbb8meu8931ZBJEndKza9VAWP65ul5jPsBZRSuz8F4yxjGnn+zxK9nCFlJPKi/g2+m6V
OA8HmBUvRIzVr8mGX+G2Do+0PuRdPqib9veKpE9w+oqg6G+ydk9q1uzKCvC22rH6BTMxTeTSuPp6
F3YBOj2jLBfenFt7vwItKIMbRG48cD0299L/qgodBjt7zflFrKWBOAItxbP/+6zB25VWXvUL8S/U
U/cMxLGzM8bmyinpPh+uHArwL3zwYMc4dOXQU3VDn40tqjdfIknskJ2yC18cgAEjSRFgVH8mVRBV
fo8UNZz1+vZxwccn8WDyKlN7yKLIHVs/L8tfQxrY73Q2sPylP3nZ0lMgDE4Hon2z/IIXAC67UfL0
sxhFoKD6Od70o2TdkS2kiAeCDLvQ5cN43l65/tOKOP+A0xLgVZD+YL4fC0CQJGLqds0quHbTpmBE
lgz0rg8qGdIND0lhHP+HCsclzpzewbXh7rHmGieB+bLVschpLE9ikB/pbNulBOBcmFfgV5/zvPkx
sD7C3cI5ypgunVDoS2C1Xci4fUA9Zi+7bDoToQAspp6+TBvC0MV0PYnzOIuLHmYOV3pYnrkvD30Z
M+/VYXYThteQ0gZlc5GNwCxeeumwxO1Jki6hncjv2DTi9jyguJQ9dCXDhNxmZ3Azcj7ceuARVVZC
b46tlWNW8EbQ2QDdAAEMyZP2ElyxsPTu6/tboWb3CRLFY/iiRBxqQ0r3cKkvWcbQaKP4L2PD80N/
ZRM4Vz06YiCgAoYIb6y4aJryeF9GXU8QGVA63VCyJpDrz5fK05nXsmFe2oHCc9r5//9wZBIznOLn
MWwxdoz9CdQC3mzKt3yihftnr7ca9niwDYe1nRabHxqPaHm/BXv+uNRogN2HszA6AJGMUVhkgtjh
4l3SLBxkG6JEEp2NaVjsYHCIPLEDJmVICYqnNDb90fxFWonEyCFNA5V4uGZ6s3PGWf1Cez7S6wHw
/Pfc2vHDwDgTB5tin6+gra7Q1G69/ilYV02lyT10FFR44JozkI8MjWWWrCKz/k/t+JZeULkFs8X5
ENf1Oa12pQvQBsv6SWvmz0urQXDFXkFxJrZWopAHnIkDHIecUVIfs4ID9sLwun10bRkhSCe/IJxI
QzB1kRc4pCq2S3mlsAcibfSNwGLRocVaW4GvGUripmmw5Hi0dPq11fRd3gDmjeiqavZC7jyg/W/6
6Rr8gCQVK61zZrC8LHn5vDb+RRcdUOBdgVM4zH6K5G/XeZXKlgve0UNb1lUCiGe7WgXF8unLOSAS
EimEe3vsJoTettx3Y13vmlbX3tr3f7zTZJIlK059BlPgn1UT898ryuYXbp/padtJoTq9jEL4vaSo
SqfDxJ+eV0KP4h/3WbQj7JdGJi44YF5UaNvZ6mHf32hRwrpdgVOG8+XL3vGgHmfiDv4Mi7Xnv4nz
CR7dJ1GchnLSSrz3cfnc7DPvux/1UIAX7wlW3AV6QYH6IqXyzbu8hjMDfaEHCpS87O+QKWBACD7Y
jKjG+cXe3T94MANlqPHSqH91F/h7O4X15fXSvVG2bUN4aYAjQdMVO1Sc32HpC8HV/eP1ZQvlWOP6
Y6xrNpz2qkZoOyP+UijkX/25aTNxCKL+veVflKtfsfoEmn5y8vSACi9Hh7g0HzRVfm0wgtfIH5pz
T2JM/zyC5dMt27IabCw8o328BIvu58S3mk0VH0xcpcujOdo4yhBUSsp3s9O2merwfaLvm43GW943
XiFUcQz+EWGiyw55UAwQF4OOZo6/f7VbRU7hyOPh88UMBI2KkqHthEM+IigOscL5TZOxFduCWyEu
bDLC+8zusi7I827GlpPZ1BXrEgtPItcLIHbZBvfI6HbCSjNvoS6OsCMi5nG7WqaWzV9/8Stdit14
DqudkbTBptJj+JmGBItYc4yGv2Z0wGwTVmzR2tYsNnUf+PxogP3D5cYKbTlQgJrQ8oxRqb3yHIwR
RMJbt5IduUF38iWE2evWoY+cKJG3Jxr/5FwHDULlqmOr9Bbnp1mjw92mlgWoXTzSgy3JHnxuaWKg
5kLB1RVLH55LelVlkn3ayDXCQvdW9Zl0BiwM3yXI6AjGELijkSon0HgmX+EFhMRLssoBcDwsUplp
tDIrytG7DX8PLC3DDKroF97nF6emXobeBpGxU/10Iq2KG6mn6+MGho+6bX/fU6u/ExYg96XLafHq
2ULyLSJ1lsoSx+gDx2pN2tkTm9p5FrYnwFXZzB86BgT8AqcVmvuNL98EUaYAk0C8p/9OkwTZ/uTg
kdOHj1WX52VHboh9F2lK9ExH6Bcb8KPJKJ1HZsb74jyeqIhdwMk6sFCYZo2k5jWYPYK2quUsUkDw
wtHvDq6pMRLW93jImHJnHO5nM2DP6/gzlFg/yUUm6YfQtVl2csdquc+S8WqKOxPUrc6wYVtsonfn
Vel5elk7CSDhD+sIWu3pEqkWfaol5MroYh3xCSnsHJ8AovFtYw0pLXScbvsLx6oyF7a44FgzPyfe
SKChQAYrv4OLjkqYSgIbdPWJ20f2mlqaPh14iNbnhJRc/J85nejUip1JXU1Sfg6tV4gg2910G82W
fpIrLrtGMebKKhjPuZ43FArKMNvDLQQf13nYZ+3tM/wz7+RJzatAe6BPbCJkwK5nN/5MGSjU7uGY
Cx8RiIHsTg0e89rn8T9WRagqF8fOftjz+sv1bHDpz5MU0362yCZyDTsAABuknKA0ZYkUhymyUQ3e
N9ZafRkhr8lJjGeFjSuD3J9Kd6j0vZq5zZgGOj1cfFseE83wiTrD65ImtVLgCMPrXTyCsvV3b7bX
0RqVkOS0mYzF7Kk6bZRWZtJ1/cj751emMHQ62EAVdWOnnl7VIhEFoP32AmrTSAkVjSVD6i21NpUH
Rw2XZQa5+Gu4PHa1EQL2FCNw8EhwqGOtJProuFUGi/KT9Q9IZRI/plt4omJoBzerJwl6DHppAw2m
tA8Ft8jjl6HSC5i4gNipYX2XTgrXxzaMMaaFeX+h/pAUnjBaVDdXuZ7iZWheu7Ebo3QLO+L14ZpT
AiQhDLFJ8vFwjFlrIVw/TNAhrW3uC/zjoc7Iv24Cr6z3ko5f3TssNWdxn6b2WQKF2mX+CpZl5A8N
j59qGn7TCQm3MhXQIwWfJ20Og4Tz0BR2P/mVF/tULxoAr5RLFX3N79TyWupjSjdTHZWy6M0hB6YR
RJDVK7eAvgTRQvEtXWZMONA2mfnsEunf+9Xv+tnmt0gvzQOVB0C6oOZzYWd5JUW2dTrkjFzg42U6
Zc9BmqKgjvXCZnG8DSAwbwoDXXcH5DE55N8wlT8nHWEx2STdrG81lt+ANDSVqGHzf0HuAFt+3VcG
i3a/67PpaR5Xg9A2V+MJNoeru7ehVDa01yIpThI5YcSAuZ9ONMheWPxfMp/69rYsfrQptbmXWwRb
9OqiEzyGcD5p82YTlyGEip0G5qLZd05oC1w/+lX2/Pz8/GA5BLTpBnIbuVQUhluv2/mTKQY9aqN0
YMbQTh6/NDsc1d+Mj4sa9tkBSZz/9aTv6TBFfJpLXfoqZDOJzJPyQ8tvCajO96K5xWTPRVJtHftf
RgwzjKkieuCMDWuIO3RV6erht7bJIqiWQVmAIj2CCHzdFPNLFdPU3cBD6pcsF1gqYfQ3rfaxxGuP
1F35HCa+JH7dKUop8bccVev0FzM5iJiRQD14viyJOQ8AJt/L3yXWeMOegJKcUK8F3S9VcDmyguyo
XYTu5g+WUED/OJuLlIJfs7tZBsmi0QtN7FUW//98J9doKi4vykVL2t+UtYGybzIzXnC9nqtX1dk2
7fbOS7R1sA952VyJCsJ7HjK/ggQvQypqcQRyFVITZZXgoh0PzvG4cXGJhx/e0Vj3n87tk2oz9hB8
PODn//I55flD+IveECl0LUPWn5qQ5f4y7cgBu5MkdXYJaM+PLOOIf/J3HkHAoJrn+EVN+8hSe82i
fYggbqbaEy3cYH850Z6F6bisOXifg9RohtKCZYrnjZdjKrwSbCL6Bg/glXc+zR9+rDAvXCRlSrHx
6V2flcsEGgV03RWnSjxdhOYbSt4H56dWBzqbx6ycaaoEQfoHCXk62WkMLY7KYS4B4uzpf3fV0RKV
F7AcOCo1F1440MJZZdVFjX4rSnAvWtSBW85Z1Ex+VbjbHpdTuuvKpDJW6YqXgH7DZC3bMMKjZB8f
vpy6PBzMjVrm1r36dICXRDRtwLmz4tssafqcFpNN2U/heDPio47RIkUJi+Kf+PPsfrLBKUpiRLF5
YonyeQFPAZAxys0h83bzy5iGqFth4YS9BY94rfpYSt6LET8WueBVYOEypNa+443tButPYxH1dtCn
8pctZhVu35rmNyBP4bT+oktU7oaq/sQnuhq0MJn+uqPhxduvLi+N6n6I3BxG0X2xvfRgKoy0Y4jO
BtmVbwm05mTb0+Yx0k/8SYu1GNLfPndo+4g7fkkhJopfocTwdmxYoRvz+7stIjEyVq5fGZ89JpKR
hzX6DaEntAboRuvJnUbJkxkoi8EFw4P53m8am6AiqVvDhZmU71Lvu4125tOXaocCECWRFi/+59jO
FiJoOh/Vz24V8rUIefCj9JqZt2cWR9e93zwdQpxNGwDCybbjIYJ1U2gE4StZsE68NxvZYSsrvCtv
gg1/hqbnGfuHJvAocbCMFhXGyWNWyBkP1abpsehSXk1VISvhi8lg0NOBBOygXISa37nNkYoqiO9D
V6M4sMqMA+H/16xGugTzzkVpKo6BBkDeL58keoaSdD4vcdkpEQkRfH2Fo9ccuXevbpQD/xQ83JCV
G/QGkuPloYoTiZ4cbTEGYKoZRy+jIyUKVYLc/nkm5LNDntG9GILOH+xEOzDzaGC6dA5Z849DeZKM
h9GI786dxE6I0nVAytMpX6YEjYNj12/3zY6uTNiGXFEaIW9R9acXeTcbb8iFShFxjin7Cm1tR8H6
TGN1Omo1WBthqhmx1MAoA1W59+tOp9PX6+mIhIZJEyxn/d7Vw2CgqJIqn4AT+eHRTTDXNIaRxMUZ
leMe0oQvcLUZfIAh5zxKZXk5VePgpZMF3Uo99AcldnE9tWLjZHNAU0FPA2pkn2kmI+hMjC3Pcs9m
+hpIh5mWq/DVsXsXtA9mkaDL1qyQu/jUKFwmy5lU89j+ShV5GKhEdwndRVYCefLSIsu9qqGRKvyi
E/pCbcJvr+rCx4K/a/wLQJ8BKzBP2mKFw+PmdGxB7Q3mfRF3Geexb1Nd6cFs6WUketmfwqfAri6n
RQXbgObtB95RXs88ZpfFx5XQvr3CZ3Q2yOOv56GEHXkC+C14qTbhzSkucxMl6xkoGxhsbeBpHf7s
dQMuBwk8khjQQOokbKwml7KXLuvNer2FMTp8TwYwBsSqMjVXiygresrkqqLhE0jwL9wbzz7SkBaz
H1J2cu0DRpGcweqNyk5U0OBlgZey/5RYfvdMYpwZqUYXExmHRTrG4KW1lhATxkYyJIWI4wOW3FDH
+OOAk4RCmbc9TopJ6bDPlrMOLg9RnYzIUwdLIaKkRhdl4qj8JgfRqEtvA2wvc/i4stPcZZtXuE5N
qc0FR1tDq6K/cEYn8KtXEreAZ66FbKa/oHsN1OJ4IWCNbVbU/o7YHPZSPNja0g+i8xv3b3jaxQkL
p/rTliU4TyvKqJvX07/Qg7Zz5sSHdFtzqqrx/44Xq6shKk9mjeiqtTkD9CcyS6E95QR6wVbyCBp+
kB+hcYskl7+cttGD5/iX+fWM5zcuk838EBfFB/Y3grU50TmQwZ2emDaa6neFaU46XnN0Pow1GrKb
ow8+qUKkVJv53zXkUTVsogroAZ9sCRdbcxu0NvIjx/WyPTKH1ReZewkvzw1UXg4YLrzrmHwcof8M
lNJsEtPNBmXgXN6emGYgx6O8h29gGm6pMmswsNJ+Qs7fu9zuL83UtQiINeuYe0f6YJJ/cXnUsXt7
E5Kl3M0nEfpt8o9ZYBdDiws+Z8UdX0Xj0/EGqcfrb0MElNVzLINutm6L+L5dJkE/ghqj0E2aYuzc
N0ffqrixOeP1xn6J2vuektzaIyNolWgLN9JBs45fhHef87GEp+BXFoUYvmBtBAvyttIZx57hSMe3
pV3X2N5yip5w9iIdzr7qr4woNvjnqducZjLp9pKKr/wDaidunsbuDOe9CdmM+FQDzm+4uXfOTf5s
TA113Bjl4ZxibLRc/noBpxkxPNasUwRBJy4BhbjwrcbzuLVvsC0oJjvI2NZwDgKfjaFHHhG4RDqF
nE8aZSrbj4vq9vdW24Pw5roEh9HgsxNya0N0Hzz7/Um7NpSlG6kIq7nnUck6RxMUzIf4hxLMA0vY
NEDbKf+ZPviBySjD0Jex1WRh8A6PZSr7GP7YWNlseqVIqftC5tTdLl6/e7iwOVezNskbpC6R5wYc
addOzm8BY+WUN7wB5uoFLScE39Gb3v1lIvHAeuMSfhLf/R+Sz8OhL/3rcNlpMhqGb+Vfr6dv4vIf
DB3nvIw8JDJ4AV4xsHdVK9LxNa0f+VRkg0L4ZM1e6f/JGz8G5/qfgUfLc/H/NBPP2atFWr+cydrb
ITg9pdhLGySljZosZXyUR7+XdcLNn9AkySKiKYCFh6XS9hnj/Asv8+Dq+Dof2igNQ5WdviPjCHnQ
AW36RZoTyEnPTcSFJ2t0/OGyHfYOEBO8BQv3etmBjsys4LPYJtNKGstk1sfUMc7T/XKPXnj/FyC6
aJQmdIlKmz3hcR65OKE858aPE5Ecyn3y/Iv3QZcnJDBiQkHKtAzdBUtosCveMkntrmpRUNbq8Y1o
E//XfMj5HMBt/qYgRIYC50+E10KFfL2FL4pBxP/zhM3DLiKRa5Xs3cwZ46Gb5RYSjl8xEK4ZED74
7FlKxi7YjEVwJt6itFCPxRmc9nf0psm1+Q8IpzcJHBpYE78+Iyn3WY0lXLqkJl7hBMwMuhy6AXyL
s7z4SJAq7J+faw68+Zcv1ZT5ejhA6kEEfeUeP496j81Cn+Dk6/aqbzqbwffx+sQFWL7kVWdeGm/K
GunfUPi/2eus9AjFn/OjD5IuWjOH3slAGg0eKihMK/nSxqsyHV7fCe6g2OV3ir8vAZB57NbwHCT7
zUe5GD1c0jb58i0B57Ec3ItLEfBH7SGGB+k+Y5vZO19K/DUFn2SbSHoQTkGkOfNlWK6xtek1ezWC
7j6f6fHCeKWu4G5YvUAmhXZ5K4XBYJAoWdBzUYs+tfa4dcXSHm0WNKkQ78Qfo10d6E/1TKgwcqit
7/3l/rrN0IimF5qeCv0hz9zq1a4vIUw+F4nn1iDjeRmGjH0RCGmDJJu/4ZbHi7MsY/atNp10ekOi
VrbQ6LP32ay76RytLBvKd3EkDNQu+AQWJqCV9cyXC6ixhe53owRsvgSJgXDoniCPMKoTZYP6DeX9
YpAteicRS46m5OUEEqj152q1FovShCP5Q+H+C0bhhF9NPzOAa9GGl3gELsC+v3q8KBqsooq0ElEK
UYGUS2U99eW0RwVLlnUv+8cT18S4Zhyq+WiHOWOSrAcvjwsE3RqJ72JFrRym4dlxX18IsufqZhm1
qsvOI7nlR7pKtcT3Ybv01z8gBeU6ZP/D2dTsNualaX5jKvUkY/IyUb53KRE+LtrpkfTP3UaYq3Hu
hbvlghK56DXCQOcYKCJgj+5tMsNgYZbyE2TBP3cDewwaPa22MoVIYJt3caNaFf4aLAG1vekAgGT5
G7SZlJl5cy4HthQQWoA4fJ+lgULf8HRWcUSumsjtkBi2Fdbuer23MANUbkKeZ+oRYijfGFZaGO/1
oI8CoGqK2aNCqSLHGbhif/GIJPc3ok3/gYa3H1RTL/dZnD7/LG5imMj8sv8Q5y7VRzXbDF0UG3Qx
8XaW64525qTGdBiucgr6jJgJuBlAwZRVX7RB2gm+jyV9bPgU53iZYfB3FiftS3lQ1G4KsAqOwDBb
08WtwfR5oJAAw1G54UphimaUsWR9lhRBBfiCGgK2cJ6UWohqJILXe6JeRKGk4pLzGtmK3GM9s8Yw
GSxTs7QjBWP5afzBshpNMr21N3JuwjwR3NItZnZkFvdchbOfCZWDEErz0rnu1T8spkbSSW5s7oog
Fg54YRIJfHSmtEkwztXqfMib70x5s19sm2xBcMTEvEIiM3g4ULWGgLkOIcRSgqx2rGopIvtO8PTK
T0c+NU4XPp2PKivFNocj2wl0voNEz8hLDHvXlHciYvSDoOJ0h0g+TB4MMutcrZ4JUaxATUdMl+8m
3ASQf5XjWrueMi4hPawMcMZGhnVfU3tgTaCKjYHC2WbA2r+2exOZ9SfcSa50DYkFsCJ22ehskcnT
0dYQzmcD5jqjJjKfgnEETcS5oGJsw5sHBHYcMzLWbsk/i7sdsnuUnn/iB7PTqLnRIgV4dFCACLAK
lWbjPAfZjw0Gxm4J9gkca/HSexckfSrWy8eCRbCfIdLvYVyzt+ASjm7U39BcCoTAWR5WuKSN4b0I
k/NT1w4OmHKEnn03o0UCjsss6wNmcxHOJm5GTVaA8BmhSML+LAfB4NmEmSV6KFjoKidib4M9nwiA
1K44hwi3Gr61/PTumJ7xQrQDqFiI1fMROrgxnPlcSfMvwP4kV2E0lTcriuLft15uevy0rvprkeo1
zgbVeQ055+rnqQTPlw80ddiAISgf8rthvF54Y8zjMdgSfCmFAof/c3HVfzkPVa+/DEQvBohDM6hU
h/E56fpoDfvDKYJqHid7SCVhQ0GJ6jPctpIRnFOlPueNBii1gGe94lGMslWurEOjS17LcZr+/fps
NNDKRezpBEcAeh+VqdcgZbXbs+8eNFgaOXEVHrJbiIUJCJH9q3UpDmjTjSK92BUhFaWV7fc/QBPt
cdbvWkuXS79PZn2Vc3XiKeP2HYiy22GId4t2k+Q1R6UY2QoFVRakE0UU5431o+nX6YEfBLgcupTh
VnwApFp/m91CWwaz5JDrs2b5aO/3MydFnRnTwQEXprqfE1VZ4f0yYX4AMcKmOL3hYv+WpCYnclQr
WsT3gEJmmd6nYwAIS9vCDn2dKywK2UnqBi8SKH4u93Mamx7TiHFnLvaJJxa193WsAVlKIJmYD5zi
9K3JdAwUjuVItIwwPDr8K3Q0xCb/0fIx4r1m8A6YO2NqWaiZ55Cw+R9pM/mHGKinybTcspTJ3QlK
IxPKYx7DbIC5lBump/+X1Tr1eA8PSpYR+lXF20gUdqz+cuw7WcH25O08sSHG6HL2m5ah0UuiM+ee
U+TcLmh5v/h0bjH8vQ7IcXE9RZ07pJGYpl3hfSTnAyfuqIoMMs2zIKjhgJgGs6ttJ8EL/G07JbI8
wWWM4rL0oytWdT2d0HBg6+wZ8ebXtHsm0XZz36KOtuKQ7rguYmrsdSBvhNbK34hZ8hw8GClDsKfX
yPUNKwZ18ZkEhRtITBS4iq50jbp9ASU8jI4EM644oGrLKtW8i6ZVxh8a1eGm87BvwwNFTx5vKBhI
74HsETIuafB11GtwfhnutfBJHAG5yKhNG3fYP9knO6WpRr+Brt0J/DB0VAHOFHRV5KJ2Nm22HgUb
YoUstyY5zm1Zn8EfeNujnWNd+0XpQPNk0vv2I/hMKiiuj7pX/OcXrqZegbV3SgIjU3brGPRHWdq2
G7qQoUO0en2xEbgoDsYKDF2bwh48q74jLNkFnNWE04QCo/IlLQgpU0pHyhojLjJMxhxrC78bSqyC
qXsqxXlQmSkuzN+ep/4WVxthM252ej+DObOcKVVz8wq+TO1rphoDxUNTgwC/a5U9dc2AaQ8Eu5hb
fIzF0aWP9LnyKqpx3HUbNjOb5q9snjKSNXYcoBpajq9OH3C+jQaavSK3qigD3URmDWR/rKbwBA31
TMv/p12oC7EmquDL53lmfs1q5ycRVIW+8sNG0jt5uPv7+Dwujdcz5++jpb37pryhAmmnAJ6AqB17
Hr67zUFH3xs6lw5cu/qd1dFJ7jVoDvq9K1pUoCb+8dTtnw4cAAvrn26nAM5SnkLo57vbzcxQZmKW
+A8PEDcghS4CjMapjJMHiQsrymXo/d/EK6dIOZ66PWim8q5j0lgxbSZRDKyTwm1vpzx4RM4+Zs6t
pVqOxOoTvF71rUNpCMYcGyOIpxmzV10XSwi2kzx532HHEIxVM78dEgeCIohKzpR9vS9X6ABzzZg6
Wiik0VExKLKar3BhF316ZsI8q+garWVMNyMpTyOB7nO/x29LeWKV7VOj4NmuKoGFagcdocPsyP92
eWOXcWCxPd3iqkaGhc61C8E0yFMsqTTQv7+BuucevFH5Kf9ywrcExYBs0BSgeuhHLcHrBkFx4tbl
fDTPiNEtgoHGtmuXoMD/FSWUXb3UW+LtZ36iQokGsJPWo9w0SS4OxGJy03+icki2QZmvWxwUDMUL
G2Z/ZtBsYR7Uf/wB2ERN+9YQg93mDwaYLMOGYWvCALnLmcthk6ryqvB7jHmLfau161WcEM86RZvU
Ov9zF7K2SFb+WUlKCn5xnaXbXro3evQRLvXttegOaJAWf3d0l4SO+CE9Y7XI1rxNdlXaD1nvS/PZ
8ozoZTxPEB5pugK8T7WChyYuU2XouG0kSNaLcLBinQfvOgl8y/YCecLEnpJ/5nqsmq6JvpGY9T/4
RXqwpzHJPZyGD4oWLWAB58rAnVjP0XnHFZFY6iAX8HR5o/trwCTUdMdtc8z1hrUkTl5I6ZCoigVq
3YFXectmt6CeyCTPZBzwMKgcaCY+zbU4dxTUxA5kgYaPgF9cTbKvSsRqhWRKoUcaZEuqy4zf4S6i
gvVxi5b80ZxQIGUewBq0qeJGR+iD+JczMvCooaWMm9/LerIIyzGrnM4H0qRAtJphTgXoeWOroZMM
aRuLj0sBcjCJnu9w627n6JXt6vWsFvjQJQzhAgZmGvsh7Q9be8demh5HI+S/HOyTRsc2rZaxycFj
HXtLAKe/WKFze5Tm/A7pGy9k3v/tS7e5OHpUWoa0pSeuNs1jFkXv2J+LTa7FcjsVdRcZR+yUZamu
k//cM6yqUsjXnqJ/c4ga5qMAb+4VASZvN305dgS/sDXsS6ye8CWOTPh/uiupCRvpGZdUJV9ypYCh
Twq/7xlIa6Swz0Q0HrkDoocHwv8Ynud4AImGU6kHYg/nY8QOTZozKlq8Fi3Wv1dSZCwYGGqne4v2
bKeTZeBJteu9M0uoNj/Gr+y9LrcLzgMzvXOJ0VzwX3nqo60CEbXzc9DH3WFhaoCkVXC3MQMHZN3S
ZGSpJM/xM8iyLjcsLcPklphBPIsvU5se7ik2f3lSdRXgBUGQOd4SEXaamIklL/oR7naiowU3ZcTY
OXzjdRJR49DZkOStnrviDf8fXUfUC4No7YkIg9JnOTR1rhgK9m+f/HzKwQhacFpWUyDUzVMFcduI
029S306eleFRurNjSm83nf4tO/ykj2hGcfJyWZ2aCYZzHFV9LPFm0OxYeY1DDYHkWr09XfVTfD/2
lsN6mzjvXg4gK1UuTK1Oq9kAl9KE8RWL6FlU4vGMHpxxmFP5b/+li4svHRz+u1MUvWyCmPlGmPvR
7qYnNvQxz63c4/sO+NJGRpFI1TuOGS3KS0hXc7qXhERioBU6wjOBoVEzgpHcKxaTZd4cqUNoSzV4
a5YjfmrIXc4guPnXFK7dFtnUPNHoJjilomgY9IMvxbWfv0j8UAld37zEqOaIG48rdFpGhpVc6s/1
4CKkqmn0lUcDlEjHdWixyP+RQ7cSzkfjkfID56k+hj5PowVWntpDsvoVlqAHxIhtpitY+kZeiSYr
5Owd5CkQOyfLVnrnDjX8VoZEbJipVaEwIogCoUaolyVLPP9b2CfXfL3DK2NKI0Ig9pY5MI0HDLEI
52oIvpvvV3ddQN6lDrPXGogfPAjFuVFEy42qAulWBurP7aKgeLbsp8yug/gs3U2BCCYJtZdGfsbb
c2xYjgSt5X71Bxfnx4WxguV1038R1S9JoGzAlEd0ZZDrYY37e3/8Ri4MtobbWcERjfnFrOWd0s6F
7brDLnawo/u9QOsESiA3x2GZtsA8OmPTgvpTmZrNYlEQSkwoTgswYjBjiRpJrMcZg9jsU8e1Qq4e
4nzcIiEuvXcjAfmPLbsj/hlzZhADYRB7JrnwIKjVozvLre+x2yzeBUXupJBOHzlOF70R3C6t5+F8
EJWJom+g5t2e+SpEeEGNB986fkU0xOOOUvPDimKesdnJGk2/uoE6n13ZgKtOKUZtncMrX4ONAaiI
Kj6OmUHa6x7rCToaO0F3ablreYheAHrzTzkmABzOm12gSio/5SuvfszlfWJDTq799LKfMP+Izt5N
vsBVFspLDj3lGJgH7mwl8FHYcC3LaV//kAWLxtD8o7dTOqUmEfB1r3UkBEO485hmAXpz8IquojFF
HLT+IIHhBMt2xzieV8dsxzhs6z1Go1VHnUV2kYSnCBebAbp1jm13itJQ7E/blQNV1ledDBsPQssl
G67A1Bossom8RJfdKFEJ3fWOf0RDRqcSU/9cYxyZ4eNmEK3vsnLFvlindF4NSzbCn1oZtob6JOYs
eAQTX4SNL0cASh7QZiwiejNBrA2oH+uoBzg0BvUj59RLUwg3a9lFZ7rdrTnBSVIPPcD4XNx3IuaQ
C49uEuAjtvF5E+4bf0iu7YYhPsktcJaIotTqfbSovNYpgiasguGMbclKcm+01IrS6lyAnSessbWL
4lo3EoZexWyRD0iKwSNphPoR0NKYdosk5U0QRaORx7VzF3LF3/K+6XbJmnidsoVbtOhUTfngpD3z
Ka/BpmQEVOT0Zref0ULX4GsJD8oBviknWJgJ4iD9IV2KZI+DbtGNdOFDhserPcZYabHHrXdzgnnd
JZ31BpJPv2nHhc/agFM295W/Bt+NNXGrSmqV/gekllhE6BKQptCxTOBkq+dgI5laoNCwFhZqOr0S
E3CYP2BSnpWzMr4CM42plGzhpuZ5avuU+VQ3IcYRtoCGhVQOSIpxQK4R8NrWPoWNBWyEM9nw91KM
IU6egJ+hJT3tDWR5n+WOURWvQse/ihe9kUoMDdc6CdlhJS/zctHablZXcyVm16oI/wurI8PuLYY6
HwsoPO9vF1UDZ2+uGc/7S6mKmCZ03MGpMC3Lv81qoDDTzlH/k6acnei47FOPVse1HrFfcLZoyBMX
/0IgMBe12s6BhMpOWMgZRzx/wgUw3QzITlrdvDgmE1H8Qc3JBf4Je+CcJfbTI/+XMTzj3UmCX7kT
YlZxgC2tsqeBV9G14w2Wxrzfddw8QgoWOK+BZPktzBcugXOsr6oDCgmJ/DCFLYhN4sImJA+7W7Y2
2OuYTKSNwOZmcgifyR+He6aCyT7cCz2Ro9rc+Ewu3NMKckeUiQ4QDyknoOGS3mSWkIzIE8FKwohL
WwG/J+43MDkPw0QTvdGLzhNUPv88p2jCaUH4zk6hxmD+qZ8eu/a+Jy5KdzTdoL/PpyfQ5Y4wN1kK
wa5VYQxhmQFgHkUTML9IKC4PMtyY9/Evp/F8psKwfeGibxRj/fJEOCJObkoe9yqy1ONzKtf3ecrO
p2O8RUoiVRELUihZUXDdtPDnyQ5wbOLp1t9TmEZpE95E53MM0g3WGUjeq3XNpgqgijmA8di0fGIP
a92D9DyjsNwRPqoBxi8cgMoPSC+MjkAg06jBAMALio1H5yXM9SWTC+wS453pyqkXXbuBNw1GhxW0
3CqkfDsYXuSFuqWm/OugaYTPQ1gAGgRXtwOHqUOTqbuGWMQRszMxrFxISi+5IelDRdq9gjARYe92
cPoKs+lifGJlD3JiNoQ6cU42hLd1butIEr7MNQ9DdlqTkbes7kS+HP2r6EC+yK7j3v8snHgdJKp9
6Ku0X7MlSIzP8JXiR2HctuOWP0CoYjv52pTy2DLRYyuM1TABitKFOm9a74cJJ965HEDFZbKbRrof
XkzGAhKvLBxNnrM4jdXQAik+mJAvQIQ9x4h5Emr+Eq8GP4uD56SNL4TxXBzk1Zq6Ix2o5nxT0qIj
RrvxPSZZkaNpIeTvFMsevYsxBHh8HGxtvstKHW7KJ7bH7NpqGJMHrlzx+gwfxmVkOyLL5A2uX9rc
MCqY7c9F2eWaGAyQWYOgwIJ0xWdTHE+BTi/p/F9xiKVlmlLzWG6hqNCVuEoFUAVuXZfTruSDdGnx
32GoPoCBpCi5qtfLjlP5ps29XdZAC0+/LG/EtJfKUX25PPBrXoEfMvJrHFjxK9BruvulpbG/CtQU
+IVm6wlMP9LVfpfUG4nkEBQKsxvjr2/G6U+X8OhV8cfg6XT22Yo0QJuCXK2Yyzk3SeUT9ipAX/yH
bIDNvI8y324ov+LFOERMlon+QrluOeCCSP4J5xv/38oO6kIUeLJ07PgkwSoeQYxA0hDbDUj8FOFR
bWXbLPQAe6btB6r0EFDdEH6do4UWjNB3qb2EAMRghIcHWhDdfZEz0pepORsfj2hxzJvELDiokoMz
EtVRZAHuvqsgVr3uJHxevHFM4L07YQnDooMCORluJL39T4JC0X0Uxes7ONqt6asb67Z6xWE3XmR/
zi1gnZ+9JCT7SlxJOx68/GqR67dHm5elzvIh0Raaw6aqSpia6R+FnAkpNnLoHiBDvfp4eIP0f9/E
T1/IubL0/Vn+8hzmOwZiDK93VetIyQPFovlLPaynijqZXKXbVjHijUAMIy2RLB3qsHFkx/wNJepQ
6LBUJkZI+7LsiXyOpfOirkUpYFKemg6xx0J0yPFIDyZhWe4dLSkZwWQYX9I9th4hmkOTafJNy7fX
we0RVZImFPxGWbDCMGKQK4JwYM4ZZ3w5oeTgClFIcuCrUR8mZlyAZgB+yAwqsZczW3sDZ0ipqDfz
xoQ3sgsKKqdRaZXVy8Fa7ZC3iDR7ubxQB10e/OUJ/yaE6NgaaJ3uSBaPFG3NH6vEh7hqnSkUWIFj
HVIiB8I5Njoo5qFT0wL4s0RsvWlFBAFQ/HU/WZTlOasOKGEYK70J+qphQmxycLus+53RDCvxeCIi
ys6K4JKW6Yl+AtIqzG4QRPnwtbs39e1jO95MlhuE6XevCC0FgwDXqRrm9QU6ygHHKSmjFGtUNnnB
xNAEDuwo8QVKuSSwWKwOFfUmo6LH4wRBKGJcbZk0UoDRSD4iu4rRV2XylbLIvkFoRrHkbS0CS6m2
ZJlTuy0IYEeTKpbD+iXTQuCgSzMyid7v22GOWPoZj4zwxNZyzTfBf8LHRIxi2+wKxt152CJK2toP
pRLelzO1o4chkokJ6Y1c+zcwqCgzbIOP1EkB9oT6RtGe7nvRBSTkHbQMqk2Nj0lKEzyK44mhM2G+
xxWgfUJFkTbQR9CocfjMEiypRxsCzwe2D9reYjgdm9oxQ534UHFY/OYa/sIe1nK6RVT9CzPdokGz
72bD9b/Ubtw6d3Q8nb7op8DeH+6EFGQjTKIuQB58dR/0kXRNhPMfBqeyHnyyYJhGsV/OQPMlMd8k
wkwUbNa3o4gvqQUdao1Bf/Y+eManjUOw/FNmlferlgxYayV5tH2u5Ny59dmZ9qmuHS+lUowJjSEB
VEEZItnG1zc7yeKfSnvkuIcwr0DSavfcLxDntppb9D14Qbw73MTqvEoVHHtfquAweFah9ZoUqiI1
94iBS9Q6CyUFUMn6LtfLcAQnkdmJjNL8Aa7wWeR312gHdNE5/xo3CSVehqzqptIAXevHjAgOgBCS
L6VoZWKDBTpjU0PC+ysBnH7FPzXPd7WW5t2rHAIlFyymEorZwE4IZyqQNehdOuhJsXcpenuTYB8X
pMke5oYi5XggVr37Numf926PTLXRteX113DB6qfVFvbybWDHIyT1qviFkj2l00pEw6DadOAP4UUf
m5DuVAfXpj6/rwVuTZWqEtkVqvoiT9a+akMpaudYXGilxz1icUnPJ9m7Z/H1ZISOLCd7dVTMZGsO
pF+qw1diz2QcgBWegtRCCOYkRSDwGqQUNpXd2y5IIUe6LEtme+Fj4FYCrmqBupG7FopQeHdWlZlY
sSmaYgYM85KkgP96zfrhtVKCCGACMvuPJN3G2kwOl2LL7tC+yZ1m8whvHevH4OVNWl1gTrVi2ACw
qtysqu61vHG672n0gIid4yE9zBowB47ynVL5JqHh81h0z/25jiFYAIijUGIuubG0m3XoA8EiHGC7
inXfTyLFCYXLg6ckZfkglj76C9WMVISMy/Sah0kca2VJeU4XlOamBvvL+C+hde6h0Rb9olnYxOE/
yG3vLcX8K5sBPjz88YC18sjbC0taRlNrFk6+oixFJ+3wECHVvlG9sjAoh6tf553BAFMIXnFg4Ndf
lbesbWYV9U9YsZ5lM9HT4ftZrIUjXimXF1L0VXrLCT5fTmIgyqY0FPGYat3Ihua8vb/eJBH1ZzfK
9s3dgAMB8dajCFL0yn31iBma8dp/rXB9q4ZLxGI77QGBOgtI0ymBcRKsNeqU3XNsqzMka2gpQsET
e/DEuqFROJyoMtyA8q+725LY9WqDZLsKkaC1T5DnPyIpiQVhxgwo2PxinBp/VvhxS0wEoCWaruzI
/lXTSiXAx2c3/FrAfDFeZw/WAUB0pZ3dbQ112SNluC30gmwWB6/9z7WCRtDL9/flT3t8uuaH6O0m
oZ457FWsk1A12GMDK8lpgIH/Q9kCoupOAKvyljffa74ng7XdeSKLewYciycZa13+bmoImbzBY6EV
epHhJJa64SPT4JFC/mPTwso4e4wAD3lNsHtM2SJ24Gj3CuH01ADjyVSGfeIF8bO8+KSRZ/rFApV0
lOMN+xoLZ9/DjFGb12ylrEtBwLJPyEkesqh+ZW7Kdvw8/HWIwKP9OqNlkByP2RuPeqwLKetNpc+K
OaVzOVtRhWdZwGqBxabxiO689iUZLKUvOfIfR30ts14ggfvpY7r1BDmZr/yFjYdnZhVSoAd6czF5
rSdUfn1qN70PRCezQmJ6iaFc95jWu17+gLrKHai1SLqV4wr3gZN7QJs46fmMrMzzXGbbXHApFTBX
WDV/VLz7aXPhOuHbQ37Rb1BmEW6kwWQCX9JxHBVGE0b2YpVs6bieqNiUmy+J/pmnz5wwTilPw19t
l9tcIn5PTxXr+QSE3+shjJ+BgQJguOKw26mAWU69/HjpFUzaMkRJmVA76OfOXjyeqy26xVzqI6xa
oejsSct4KjOd2qfVkLrpx6lX+ysysA7BndfgCRexzIC/i8ibOe6UHVyE1Wtxnsi6nRghArOLvIxu
0ERXJHejrHZamPjPHp4EV7vDqA352rO1VLxBYUTYGlNOTVT8w9ZTOOvkYgHN6evMsiWScirupE1e
YQfpt8bZ8v4k6RCB+l+j9t5B8bpEAOhBY21XdtxYeLAfWjzlnpJH7MRQWVB7enVsXqAIw/fZWRGt
8zPavM9jyVDN3fL5FCKfgy0XyFbIfWGFsgDFsFq3+x+Zgbtira9ADNHLBNQXNlr1KVxdvqQO9VqT
lD/qI2OjjSZUTNWcv09+zPWDYMWgtRqAdVm/sinmI3XAHW74JQnZHg/cv3w5TT32I1jwvhuK6YGE
AXcwBrWDvn/mQTAb42K+BWBoaIGz7hqi7/FNj7jHUk1zwsnfB/2yV9w74Qy1j1zwBkPaSrJ7z5EF
q7M90DJCW0wLMNQINmX4vZbL21o+BshO6jz1YdVbqms/4k45GCDGG7ZTRntJwvZ5iz1PX2RwJ35+
dSD3zOsabWYEbTO8dx1Q2v9KpU4jhETJyC7BWt3kdIOwj96QhFWikiI6WWdkO7os2EUUx0bZcyVD
WUlcgeEuVHveFmcOVRsfPYWzKU3N02cTnEH4gU4NLu5XGJhaCOknMHUfWl9TVRh8sva3CxukpDHG
foZrnNV87LMTrO6EQ6Ezt3HVyTkcsm8M/mkAz0feAAuXZSK83KRlZu81uMJQ2pRrJOYs9P340qQ/
HDfFgclv2fRxLDEy1t2PyWNG+ZVfb9ix5O3lDBLsuuZD+RSchHwcaiUbLY9S7xljKqIV+yMVS7gn
lOcXhMI8oUNrLnOs/xJjQgAjoiP8wlS+J9dVN26xRypc9ZUgeBzPI5r/GMP366kNgj4sbcLGNVmU
28IeCHIVerp0hF1PuBt00PwLYfLnWjTJb7xznUdl4kZjFBbJcnqf6sNkBTIaVQ9sWxWsz/32Dtr+
lGjiTuPNdVfHgMSnhjIDHMuDoki76n3DB7QKiMMyCKjU3L4ZOt8/eAZXtZW/ht7SZLAbdHHhzIZk
x+N3B+w8PzjQOhdwanQy+HoaWuwJV9uHCX6UhGSZJChUGNOSfJubaTSZEWBaGn/M7l4iwF+aCJhO
KvZQe7iJCuUhdun2gV24KMtT4Ln09YyStmWSFRWw/cCSthbc7u+xKt4YCtenGLU09MGMMpez2WYD
0bqJMlyhou8a4MEYHhgYg3Ij55cFJMtNZKgEcIrBZH2TxeW7euweG8sI7VvfjwFCPJj/s4z8WJFw
p0q4K0UHDueR0FdGPbsARUQvLoTVvelb7m4DeIYbkl7vUX44kKxn5OZbm/mf+sEQpL7X8VIiKsRQ
pbtVHkiPucWv69lhpYMRgKLVbttCz88sA2FJU4nZE2Wiqa5DvdbhHt2EUTibGYumvhjO3LrnjHiY
Eey8MPjpplpRoAF2XT7qxvDmBaSFY+b6fMxhE3gvYCqxhxTNO1UEMv1g/51orLYxrYWjx6AJl3db
szCZYKeroOW/FRR39wJcaMwLP2kvHxbutFMts2k9a/jhyVr1yrH53z7Z8KANeKJKsMqXDQBU8uyx
y3oCBdeKmy8hYlIwWGuzvfi46qR0sjI1u9jAFTMZBKitEj2mN88RkRib0mRA4HHiF49yys/kYZDk
AYzmOLtZNkRy3wiQlgx0WAIA+zsOW83ln1zy6Nz/j2HxatUkPDZUTG3x6QTtFZ91oIpYp13uPsdf
tecdbLXxsMFGaPNZsOIzVHVFrFuMQly9N81l9nRjX2cl+hRGJ9SWc47EdqYyNHIk+f3dy/+Rh7YT
yjynk00FowGc7iMTlACD1c0hONBtOQguHy0oVrYtBCxbIfHcz48OHcLN7fTF04hAcRLcDnyKWqg5
p81ItFHlnzVRygbaW/3KLoLoHA/RFm28lMopGO/zGyfnjKHFx8+s6xv2sxStqs3eSLd0/OwYNfWo
Eqa+jsRXiIALs5SDVph8P+YgbkZOxqia/S9VjEN7IUn0EwwwhuG1GCFQ3toMjMX9LGTS0QBileAR
/3FOkFl84MST+NsJBGN/9lUI7VYMkhMI9tE7s/ljGxTPyMrLpC2qSOwdbVJeL+oHwOGvQO28iNpb
HTV2Dyh6lZ9uyfbRYxrXcxY7JFtTPKEJFuSyjhtFYLrKfZ5TpocfloX1+rm31znkc5mCOMlgBi9O
sM6JhnYEPdt/rDAmw1VhT37Sr9TpKDcEyLYDyDHN0VASejHf7ik0RJT1eVmXYWhvpnVjjf5Vt1Io
gPO63jsevmGnnmcNxjGESqwDt5jwduLi54aSOkFcfB8VkE7Y7r7FuDbRfAzrq+sl7RtWhnQoPS+l
H4x/MCt2CdG0NYFMtkswJU0Hz9WYG6xdAQK5mpCnj4LcYNlzLPBRIRAjdDwFyU/CAeAx+7RVl+5A
PR5PrHr7KTkwR6l60CWzXl05kW+gCicE3tpMpN+YhgBsL9Rlg5k9PblsMf1W0FIPFk7BsD4xKlab
Y7t/he3UlOfBoDbetM0mkaOkYlu+jtsGkSeDGOs0ssspJKMCbds/JFpVXA+a9EQWdRa5CuUSe3lO
Maak8QfrrmoiPLIZp7/BIIf2tu7bSjyM1mMTRu9rYYnxc3wnUHCFpTeZMG6yonNvwUqhmC1auGps
999R8nUVaVEJNZa0Rq+qvnfgkOuLzsJ1CEXWJDDYXGCaVnvokxpwwZZNNXjTsDwrjSCWb3/QyesW
65qZZaLcXaLZjo6wEQDVvqGsRydC4LZs1WVbjBLg39jMqVutcScBiPFUCDChzNEY5QTW6fYKjJVn
22V7DzkqMhZ6qMyFWv3fcBiEeDPu/hpwCd1t0fON6ruVrCoJDCqXyuQYFEVSKEg2nYFjEmZumCX5
8WksKrUjAEVPn0lRXvW4Tu0KRClKsahMhi7bpk5NFACysR9+La0Smr4v7rYjFtGG6eGwXuXHh+Ia
NrPAvORSIheTBk7eK4LljInYJEyqCGKHn2m+6SnX0eUpVV6g+qU2ic97cWjWthyYo/I8edEURqZE
Tj8pKvKaBI4BM1I4FDiJ6bpo26RDwIPopz3AAtppNsggXnzNjiVfRXb5tLgZigVBNRN+PA4l+dsz
zEFYmo08YYjmlVnZKkbSZjjCF50TI9Uf5Id+nW8HeYAmTMvPnDWgvZ1zpofsN/K/TF1JkH7D0N8Z
vN/HEdGEfGnyG8cKl/C2FjYJbT/hiETspYVY8yjTGjxSgn6AX4zwQqErgf5a19rCyl3QnvTs/IAe
c/uVPTCR9fR7/thiZKQ0AwUJWU5U6zULQvYxAcYM7siXivpM12p8WdStId69DeLxIqEB/6zPVa4d
t+3vNxtl/O9XAJupBlch5ehmY+ZcA4oSo8Onei7qgcrh5SmP/gCyCsQq1/Rf87w95ATu+b/fwQN3
rO7M0YAR5nCDB184JPvmkjxHWDmNRcfOT/DQnkm9L9vnbC/ZpcIQVgmexhGEQRWSadEqJhhw3aOg
zQ1ehszieagxi+Q3dK5l5Kg/XNmGSx24Gnr5ScuiYR2c3bs73uS9wqdp9THIrlDs8D5RyT0qVFY7
6n4C5+UhlBqaizvTKOJ4NvDVyUjbTtEg/mtvsflBHrguYHOdLxvkgg7vrkWgHFQrVbk+74eqErMr
+Z/zt/6S3S8OsM59zwHmJK8wjrI0JYfkWMDDEaihBBDaWg6wenm3AV4UQ9LoOp3A5mHWpmSEUOgv
nZiDs1SJSTfgt3wnCfKvwCZAX+ZCXSpmrv65yPqu4hUq8tXYdmAE1cV8IECaauDVqLgiyO36m03f
HJi7R9nY0SrIFNAyoH3EcXqcXj6BZslfpseHGAitO3/bXEj6p8iqvekQi4n+uyM/OZFJ7YxF3ijC
e6njVb079M6wqMtJpPE+wRu9ua0fHU5FopcK+scWyZCzJA9YUjboCgmwIzbpifwFve0/jYVo9GJi
MqIflEriW7Y0u0+CZf0G3Uudasq+eH3YhAQdc8DWq+yCls64wVvy6YFWLKGpNMsWCS4i4CPJTuao
lbX3Vz/4dpdfRf89nKniZ1eI1RBN0haNqJU7adrBJ84+xOcXhO0D/c6za0WUnY3l5aJSStCEFMWj
yUx3AXNv1c0UkceJ1867wjc/lAcqTygzXMjK634ioVbi9OkgKDKpz3rQflG8nrEj2LWBLHr3V3Ky
LiTKLbDk1lGv7qWaJlQN2NcloEKA/RK1F2fZfZeVdfSUc+6nD5qKhwMrr1fuhecwJK/WEY1aHImO
VSq+vDDnylcaJ41rpLk1qREWKsJL4LaAgDUW8n1N1UOlsaftWwQTD7Hz7qXM0QbMpA47wel0Etau
cCI6XUjSauGrPNHiUqUKbQeoIeOWf0Ckk+XmS3+vIoFREWpUf2p4X8xsmEyymEyt/IRdlXmoKHNW
8HA8jGYGfMn+PUc5iKH2xt5hX65bXJtnLAyKFZW+6d1/9owwaDyA+RMPBe1x+GBuyst5yRe9JEuQ
mB3Skyri0PRXi3D5CeoLpSSg9+B9dIo9t4WChhTbkAodWOmoByHyTb6pmd/PeUfVrnySAWNgUQMs
YzGUTZD6fjNWreN7VcRSnexgYrxxaS7ajS4OddkVTqaCHU+R8TLXOBEV8Qbhu34mw/YZRBaRzuf5
OcVYkWDsYNkVDDtMki6ztKmfONbbXZ9JpKhpc+fcFGf2E+m/pv8Uh5QGLacOp6MS6wkvIjXgMuLH
0jaSFyGBoJTpZzMlSldB2t0cQEelpWSCfmzsEkz5YTG63LsJikB5o0oSEISXpsDE11vGhSs46cEA
chA/FabeFwA7y5dgpF35pKMOwhUyp/Lb5stYb8/ANsZgdjYonMhU9vRXqGOG1K2gi54TFAHkBEoK
p9M02RO+kHp6Jw9DLKl9lJWqVxJct5Pda5ikNJ/12tJe+7UeHKCXKQO42yi8oMyBlIRm5f2MaXXw
7Y7veZ/MeR3ooPbzEkeGYJW0obYBiVDHzRC6wPmZN0O1bq8yCbvWbqh+Fu6reRwHTTp2m/lv8BmI
0Fj2s7/xujiYH7NtSioFaMSh5OW4xH7J51cFt3q/YxrWLFkigwpQswQntrhUXLRRdT2wFTR2cdtZ
Kx+SORNrRvrd3OjC030l1CUQ71ITdbfhXo31bMMbNRejioU0To2Un0QR6rKR4biRTLF+D+ZVwkAe
knpAoNiPPD4hLxgK6YRGT9jW67XlBQvZ1Sp+GhozmUhKK1rQ9csZ7+odImwLDXHjTjILmqN8grEP
d0dj3+DNG1hPVp1Cez8Z4anuvI+ktdSqXcTjUZ3hCX73OJtJmc9WFc+mMsaV7oWwKO64B6QovYp9
3n8DZIps0pGd8UqOD9Ioc4SLd4TJTxUb/L/usuJc2YSu3q459XBGRPiDO3MPpkILUHVQT6ZWO/kJ
scsmR9sxb4D5+2rdRmIz0bw0pWa4RndCRV1PI/C7NFcbg19NriOnGkCIRh7nY6TBYU4DSsuEodHV
iww31toKCYwNc7XQsBcAZCvTf/pvprzSc3yoX35UhimbZO8I/crlEdEnV61Kp0d23zcMAl8+KdvE
d8Vvl2glevcKai+jgsBXNEWOyP4XHFfLVxO4Kr9cgP6pCtfJzq2RzcpcW2YsYABFpMpiDNVHiUhM
0bi6kdS03IMTIGRFHNFaf6aFTmeGA8LCpRecXUUL8nYYCWNWA/p1pr1GY6msyXNDtJa3ibw6uRE6
N4nMNGlZSFHLq0qt3zw/LeSg7LVJmFuRx3YqHCU6rYopPkyBks/AJ+RZEVY9OIOlwqyL2hQwN3xd
zaUd2fN1u/M2u1qMP1ZUE3LtV/nIpAv/upAbzDN68wYcGzyaKNNCIXIBJq3S08AIhzmxKuY70pxJ
Z3Q+dqb6RcEwA5BP2riVqMTq5s0Gn7PGXxlecQXL83IhFFtW/2dCT8tTIJPA5LSs5NY+HLQ3GcKA
WHiuisa3SMYfsoqMLTMnfkpzRaUvZyf95EqsH7GA3L+looTcMyvkk4JHwbR9ODrw3sZ9BrbB4Ico
7OMwKaVjG/1WfEeVyAUbgTwPVjLJGnY9Z5z1b3rDSTojG7ZrdQOxheca2MU2n3PhinQVD3YCWMF3
RMK9sQobGaUUNcQhkKPsPM2TjjsNEy6NbYarUjx1gApbMtbmCL4bO3KYbc9AHYg2D9+FuHaxLIfF
oy25+I5dxHTHZlBrhdnv9nDWQ+jUEm8IZw7A/W86ZVp+wq3wIBTWTXqGzNA25UjxHu0ZZy0WRl6D
rV+rDUUwZALDKrvvI9CFZ8kuWL0pCaLT7nJTpe8XpXDkhEG7G6EgY6ab/nxSXGk96KGLa6aHXpJM
8zufNzz9FLS6G4WWH77J4MUHi26DxVU8hzMzXk0J0+CasEwWW2jRiGFPkeFe5WwYcDrzk0bfnCOv
5tdeEYMolXbAUikLLkE5SD7QvZdupZI3iLMpPBv4w/P4MUiwRLMqhy+pq20bcbSdM/xqSPSt38FA
RU1tUqIgvVNPCSiunzPRLbKoYRxUpI+Or9nwg5btWnPBpVjaXG8TuIz0oC/zgcYnt17DUZQfJ4fl
LZvCe5rkYPPzkmOzKhV1OSnGLrdAnFzZkA1XwLjIY7UC4LcAviQFJQ5DQZKr5SEQP6qriaRufJKx
SZlvWS5MJiXqeGnwAHbr9e/76qT1z9hiH9GI1ttp0EoWbGZpmw8bCayCsgSMLAWDad7cT8k55NO5
B6RIuvcxn8Sk+8Enkk3tmJy+KOfnXzHso5x3Hxm+e9B8YqUP/05z8kUH9ChUXU++Lxwetj1kqX3B
Va9pN+QW70QBbYgtYWD2pyV/V7mPEhjZlEtr/xrzDjeHWbjldH4nldRNHF8YTxhTjwhqtjyHyxFu
xMOQ/9cRijrPM5OZJpUXVQvXPvG6KUc8Di7KI0nweKV0nG7xvZbPJWLBbWp4GdNSVHE+Lbwq2jzq
icjVOuirviUmENUhtdCLCOnLimha5x+i/nZgsyqcR0svuJvCP41h2DoaZwdivHCdjfmVCCUgDeGI
NTJ5PpC6JBXgvv7jDQkNDvsUHpzodFJKzo/HL0xQ+kURLdTnQueVivrNZT67gJC4rlU6ppyE+T14
idM6oC0kyMCX2+3NDVrSy3v/Wjfxbec9MdOuKd+nlo+3mR3dPS3lPhrPTOxy8VPewmO2xB7JiVwJ
3c4JhUkwz/t9mhCltUQ+MLMpkOR3F7mpdUM/Zc47NOV30dVy9CH7T/TENUsIUaEcOnivf1GZZZZ9
lHvOM/bglDHvnDhqmca8SWwjIKUbtjgRBr8lDg8wGxz+kQa4cGZeh5ed/6VSSCoIy46+fNgPkk9X
0vMZ3HPDITkoEMLDXHEVnoo62/RLMFgPqet11B5f+rBj5AnLDaf2Hkxn3qVKrdeHo314Oc/m25nN
Vrtqy0TCahJTBhW5qaFN7P7M8JiDHIzEHCRCzQo7S34YroRk0yfvAUqpeZNmg4eYlYfNz7DJX+Bj
aL+c7oxeQPl6XNiQiRymmU3ClHIEdF5oHtH62wjrApyaq28Vql9ReFnyCete/1EU2qgoUjvqpoNy
dN0CJDNnaSDJJ2ztwtNwY1rgJdyiNOcZor2bgtE1Qp9jS4tT095jjcP6kZqrlNBnTYI28f8sNfsB
DN/z6RnmGHWEFQmOuU0kZ9g9rfrqSnAIv21Ze+2TtuU/ZMGUxBHakMR4Zu0Wde2nNjXbORtlNabh
x8mG4nP4zEDpETl1OsZRJPKhh8T6v+nBOco0uXNeceX47r1DIaf6PHWb0qPpwV6x4T4mJgd/cg01
NehRnq4QlJkHSKD4Bf5hvbzWjqbsOUhiRZ3zD/oS4xB8MP29YijpdUB88pQJRbj+WFgVj+YrOgAh
ZVnP520zo92TdVi0c4HktVPyTh4IJ64WLy45/w0CSJpxVHhOynGsxM2U3E0vB1FW9W+W+fDH3B+j
NKeCBbdH69wzN5mErQGtlk1wc/x7kr674jafnU/LnhBAzt5NIEtjQCdXudymlMC6OyBysYRk7+ds
wGiYflEEt+R+ikGWr7xSGGnhXmR3lsPyGdiOu6NQh8LFHWli061dzNv4LhvATLllopnLJaxo3pAF
buy8d/jOuzXWAmxqNse4IxH419JFEKNqN1yG6Tly62PQo+1axge4L05+eZTj9LYqCEkbci+KK5Gy
8K68LAAHqpyVImKvLMV1td8R0n0PHzCbIS8Kp3NVQUd5SzkF05vkHNgx+Nnw+DVDvgx9NSuMR2h3
SZ0UMt/e6M461x11akqeEl8HfExt285qgaIBUWWMy1MooZjcnQKXTS1YJBYWF2hdsuEe1KOJGQd+
suXt1dvb9e8gF2Ro18OuZlnNK/l8/ZQ7g2CEOtUNoVChbAKK3uDWJSTMOjCILfluP0zrHqwWeQoK
rLDLjrUEpbAYlmG4MTF2zyS0Xa8eS+hY/AkVEPFZEF2W9F6pjgbEmzQGFXW3k+ZB7GgLs/zZtOTW
fw5vowCGy5tIFC6K1HW/E73ALgUlk9n/8S+efP9FIpGp6+JQRwnt3YuXwWLYa592n0pzPKppwNiq
eFwin7guOibLGSs6bNQjD4q8V65+FTIooQo1aXc4A9EVo8RjJFrPxDZfQro0ka2+VaJQU78WZXgi
ZGiGlVzs2zv+Dm2ya/LNTaN5U1Y9bmLooExXvDa7eNJLxC7zpTiVf2C6DqBD6kO7dyvnMblxC29z
1bShj8ihhsIliUsx8kQzbdYkWA2eUlMcqdaAeaUWOx4ygnEVU+zWgQjz69G4Gr4bi5o2O2hPuDQO
ebaRGpPi8Ebglt10qfLRLzSnfPZvGIbZNcWN4JrWSOj1K01A9/RxEpDGlQhyL4JuvOSzbha5PIbe
upyTbktxZpwkQfoqq6BqzcMFjCxsnbp/2gMUpnMcUNay3YNV+Hh22oGolXu7dNrNFFF+7aK7ADUO
7QCydSC2GO/Jpw5jV4BsagAJWxGjsociBGNNAFAvaNdEor0Yq3OQ4amrsre/md1NXg1mp8cHCzzt
wUKzZEUMkXTx8hKULUGgqpCGXF5lwiW9kP8cy8jeZ8vVuPnoSFD6Fw5lXteCL7dAsZa65vKgVpSg
xAchTOo7GdXjfgla3BDTmRG7ogBJ36WHbGe3eWIBzcyzKFSAw6rDJaMkdBXTBbVXIkJ/eh14mdEO
VHg/ncVDPyWn4qRHs5sucd+y7vMq4dZpdNvYqavSoQiwtK9ooyDZRyJNTKFm94eEKAktZ//Unfno
kCvHJtXy/TldVwgW3sC3p9CYKjfe6jg4rTYEgvokt0muXbOkCOSLMyAf0r+qoOKmBQ4nYvVhODC5
cQAI5Agnahn34202kONbwNhH/mfbsHuQHs20uNvJndRi9Lq/OtVaeU9Z/HXAl/owq/TNEPAksA9c
SniU36ovQcM/JEoCrHIxoByNKd5Mb6O092pU6gX2Ie9RJSCDD044U/TjYs7PndA6oyK1uv8cs4+c
ZSDaeO2n8q6SAvHlg/wCdoFo2Kc6Us359kqC3Eap+5F9eUTS+/Wd27D7NY1+2Doye8GEL6qHcvO7
YRqtso5Yc8htOSgifSHf5PEuwbgC41QY58yJNDDmAhPufJP+9JTwC34kowZexr8V5Xd/PO6q4dAE
poC0aPjB3E9ByrrTcXBGz2rQELyKioFHsxKEEdX4mdfwKDxPiZDKilG/zcyowO7InJKDnLkPznhp
Bpcmqn17Etemp0A9WvDOB4zNjGWiADphC5/kwcvDYzZtmMDnFkpB1AN5On9WIuaouFyqiFUycSii
6hUwiJJ0J0AtTdd98i86rV/8veJkAEdCPP3DDahDyVffdUYtshzcLnE0WgduCp2L0DACRsscKX9f
b8n0XEF3mNGJE94+0lq0P5oshrXDvUfWnx8WNcgt+hsJjhtRUVX3eD4Kgts6aptMYG6TbjtXbM5Z
ZPiM3NVqMLSPVOSru1hO7+zQbYtU19LEpRGds9F8ibuIZ6G09rHMqf/+h++VgtHbZvCCgciug26z
+CM9ppmfhpEWirY3MxAhQfouQD3+fkV/bKsMASodfAE+FgsleB1EkTYplY+2DHRy4543grPoAiAV
5TxnF+riFWo7leMyRTL8j6ZaFkalGRTf407NVbth9x71cQbnf/PSlWma3gPG8iOcjuXyemstq42o
zAZcHT67gmvGbxWW4zUGJAjbKIRtfAvr6oSv6vdQewvtIzMjgsITJoqBdqt7zQGnnnuJc07hemx3
yq2mD+YMWqoJR37qsYsHUZVYeGK3KlXvQpTmJ2KA54Uit/0v4BXWT0EZXR4pZdS2Di3zl3VwAgVc
z/s9gGFm3LUMkSfgcvTDUkRCG9tyk6Aanstxw1wE6BEkDftUh7+pHR2OWyrGi2BICsBxGEssHZ2v
VKHFReJ6fYcJaSJvZnQBxNoh/SsR5hFgs4Dnri1id1bz2MOdzdvCx9QS3WKfZZMJfEVF3/CiXB0x
oxsst6riF3DSE8PB8fpt7/FzuIY7SwHvJQPPQ88XoAlLghjyaxMbKYgl0E7aAqrd7Oj99UoFSodM
JS7BLZCYEZmnKQ2l1peu7WWErcneutj53NZ+klY+qzXXOmwXEGDoHdeajOoKgQHqpE+Yau2+mw21
oT3ghx84NCRJVLEgxvZ6wej64hUj54R8C+MXAPbQkMEj47m3oo8syzkdgth+ScuPLnMv6ah0Z5wR
ta0fWYTjP5992j3JGlz9Oeu8UleNvxJkK9Vk8enWNhRAvc0Tk9Jx+G1ARMifRbxzyhMf/vFMz/FG
H1l3Skac+pbSYRaI4eFErHtH41M6fScg9rkfGLNZQtJKgocCgg7rx5wglA7rDUh4nHGuX2CWDOTZ
utwVKpQqOxx04QM8RDcZZ62lXAFhoOa/ZSMB221yGJdPrruemzBzfwVeKWBIuBNzb3uOzwfUQqRk
SuQFDvIs6HF1r46b29fwwWLeoi8bh/5MPKx/GUWwAwGdUGbgNnMpgKQcPS0A6rhegbtMGg6TpctH
yoAu22vk2SP6JIjhcrws2ot/W1J6FSUwzTOdYr3A6ykJFyFeLu89zJQiEsR1gdqg7N/II5utJNzt
7ckjeiSUmtjTwgQOKU9NuZLWuD4H1OR+46ckirF5J81Rg6Taqj9CqlEmkrZ3ITI75dnOjJs3r+oA
cTRnTjKdBQI7olPZxuAGv2IdljbFZznW5hMLEZ+eIs5agfHQtc2mGct86w7ck8+GRHfrOH34fk9L
hn+/AFMHW9k+tmcYTo7PqOG6a4iaLTBStYfFeUbDr+Iihyxtwx5jUdMad93CjMiB1hYz/JgX3tkv
tNOoTYof7WHkEZHYqztnfjw6UMzaCanjURN7iBjESTjDa0Yaxcic8kUHP/7/3DMybhAtDZPFAOqU
baLetrRuUcGJbLg5nab1DwHN1Flv6tYbBtWTEuHCPd1ZhfobNzeHTTgJMbVHQqhS94o185usCnrC
xuVda3ce5MqIMNjtnTDFYjJWjscYr39wR9qNBhWOA9pkJjjuLpGzNM8P4Ygs8/yPKVUTXkUsja65
Wp4bntthX5DcGfpsBRHXy3//El701HCihK9lZzACzpMQrg6GRZZ7SP2pcSbEScaT9gtwoqGhv333
mF2bxwicvnGpmuUWppIUfK6FrGh3TDB5Az6kw5ZeJI5EODMixXQea8N1yAlX/sCcW57yYjbSrj2S
hJQ0oAEPNQ9gv1Y9WFypK5jSR97/PzoACOf7eta0oaQbzmJOP1Bi+QpLDsaSsZsBoEw+GSR3A6os
KmYBuyT1YTh/XT9iovuLU0MZdmABH+1TUOccZC2AmNz7zt4xvKnbgC2qZk20mV0gBhIc2BRokmk/
Ucx0sShP1+hUMBJ09uQiyXG6d27lvcG3RhQ5lgjK1ynZnOo9xm0cuiw/nmOPPFlCVisy2hVtSTlJ
CrO1OoF/CEMyLGoueWh315EZAu3AANzQNvhDAQrng08117SZ6Fvy8Z+iYNu6bPxlXYCrakzA3Ojb
0XuAQGt0urkMnnjh5tnDhqV9bq9rpWCrBwSwdlvwSCNPewSgqE3PUAML2WFlx+jFIT82U/PB5bEZ
fhYLhLIfQvgwMSe/gQyqI9kB1MYkLL/3BKb7oitAsJ5JZL61pHmxeN7iwitPLOi+2R/ARHwtLR2L
muG4nDiXElkCii7v9s4p9dMN4VWmJXYcCvdWJ08VhptQ8VXgOwPZ96Y6xyxYqfZNtzod3VC2oegF
YDb2eyoiJi4hcTdQPi+wk4UI+LlAc40dLlIUrygt9MXMoCa5G5POvkkVuj9NRLBHXgpyqkYWspUb
zblQaa5gPFWG32KX0lCForhCab7JO8isBB2dYOby0ol0tD8g0rBhtdgiQrnF8vWhNTHGgy61bCA6
g1iWJLpKaGw97jNKo6ygRwvnuN9nedcvnsCgS41ZBQGumxuXa2ybuNAx6Me8GI7x+7H1H61w8Vo4
5aDFj0KxpDtkHi9LVuJTk/7r2MdVllY/RxIRImT4Bd5sZGN1MHqwtPDFAGhh2qNqJXZFV47MlHcG
sx30MhwBSg7Fj0Y79klCxu+LhELTtdc4CHoJfi+x1AaA39815lXciC4kD/U07EU+buVg9n39oD/k
KtOsmHZ8BubweGMtCcW1mZ7BdIKaUamhn1OkdrLGb8GU5AR/0zPeHVES0SLPpiCpnjBmbg2DNx5e
mi1sMUOextHj2QI2dkJFHSDAygY9ANeWChrk1tdJbG+le54sVzxVvSPWDma1yjgPaBaEHxKn9Y7v
q3K6FDWx6Ek6VOtfDWoqOfX/Vmq05dr3oI7t+iBVhuw7lcsblYA4Qwozhz7Jo4tiV4SIqoo/wkUC
0fUFvMnGUHXeVQHiKnG+ryqaO2LdbF8DsbkzimSi4hKhJu0up27nubkfyffq2zCB5qK0XTW/0jXP
SZj+bcQzHU/7HHMIjqdWqXBQMVFNmykMAjEDXs3c8IHZf3aBRpqpBQoo1WdMtOelYaKvLBrPReby
EaoMYdG9RlO/dDdLwAhARQv7M8vJlWYFQ3rc2ZTA3kPX6svpcyB+LI9SEuNlqZU0mPUfr3lPj5Gj
BsjRtGdKrITViQYpFGhT/PyJo6GEZY1tqC6T0CupsKa0w6zM9Ym7ZCi9SlYkqOkHQS0XNxdEpGIY
MB8CM+t6CeNdn5Xq5YQvZS448UL9aL3y0ArCl/nENCptJwjxstRphdhkjgEVz9fol25M7u8ZprJH
oX/0DRT0zxfr0XtMIJHAB8Z6a7/fqCaYyFFR284n4pT/JiTITLpwUC0p32Qc40xOBWNrOQfDVmkC
k1qS2Sm3ukZi5JZ+q3WC5YN7yhC1BvjTcA8b3YKN20rT37uSsUmqSwnD2/IwK+bFu8YE7Bcnb4X5
pbIEP0NNUIPhHr/gGIFphD57903l9M24wdmK9/reUzNgQyCYxYLD2+EJPZrC3Gz4CWlKCK8MLN94
0NfLKkfkHYddyAuIsV4ILkwgdzSG335VrBH6aMNG79BNDTpUA0rTFRAp7MRqaBj0QpNKYnS83cdQ
etfQR4E57BuE3SX3r339PwujVNE38Fv2dX0wC8TY2TskLFVDFssox8qy26/HSSEwZ+NzCR/lwWTS
bIFfSMWdj54sO6Iw05Bv4QJE7Vk7S/ctAXOJclK9W++1bVTtGOlIbrIB0yP5DxFcIH4o7nWgrSxM
zyCwL58NtJco9EYm1rg/0/vNKe87RlYRpgzVwU8Y7sHLLcKljpdtgo35zZFUUGeJFEdsjHmCLyqC
Q0Ld1wSBRy48Orw4Wfpwpr5wJgaq0uwbfBk/uxjQYHkCcyOGCkZzDBXqF/NbSMk869SgL+L6RhbC
cDi3art9Y4BuC85OZ3AfrSlLAinJhS9i4S3y1RiJLzFcGAsHMk/TSfRht+Mck1PsA1mhX4T/a5pE
4rr8jo8AVKmeG5CLsouMFmUc4f1WMWndst24yRxtTh6gWaul52FTXZVKoscrTENCTuWd7VleZiXH
es3FLFa5Uo/ntA3gFoah5G+YXAkwbg8iGYkUt0JMFIQXesy4eslQ8IYz9L4ycn/ifgNsizNFk9yA
NpRzLgHFn7BdrgCfdzzJqyGctJDrF/lc5Fm2pKMKHiT9YnddTpH5yfAscrTUkRaQpL4218WiQ92s
SEL6j1rw1omy8xfiWXqfEDuCcJZeQSRi5EWXGReNB7jecusNwV2yZylKbV2H9PtmyRvGK0vLTuyd
RsgljX/zESzDq6j92WafxQQWMSZX5Vtp4vVCuuWvfdexwf/68vX1BheNfAO0/ctx1Ilroy1HiC9f
P6WakixsAowNukAcOPrWOQKLLRW4A2bnCf95jWiS3RGkWnORfBA/OQL+K2dtztWsB73CLTlkiYzo
evep2fRLhoN23eQfacgRKPgErfw7fFiHTwloBYJ3c5u3rSth5TncrvfqhgUjyQV2LcmIFO1LPqam
Nva3LQnwdC78fyt3shDjbV4KGfRUFEBuH/+UGl2ikrj07krPqdygUeQzywih1xxMmo1psxF0l4cg
w8dHeDdFPJFb+qmnXi5aq42EeYLa3xHMxxOrfiTX+xf/GrcKMc2k7JdAX5Scfls2rfiSkA7Zh04O
LvceeISSS0hcf6mSXasY3OqfgIaAF9KVq70N2VKgs+CQNAvMs6ahNzD23UzCjdeBjerhvD0QsAZR
dKskhPeKT5fVW8qd3KTUj3V8uAKwvwj9vTHEcata25wMzEvIKT09Ebw7JLmXW+DBDPs5j1LMSvdC
ajeKaxvB6STuAt1GcHB1t++QNkCBaXjfg2a00CASuRWNvjdCMwe26oIJR6ltTGyJfB3cKGqfDH9C
4ZH5cD9HCQGpuo35YPFzDaXWTtuQfVqTz27PwWTCVpTrtcydafBVCOaIXLVa7qkH22VtSrxGG5iL
PFfI3hp4M+7rwkD7hdX9c8ieGP1B9Gha9aO9flg3+r5+LwMeNBuVRBfxf/vL/FvNL2Y6tp2h022N
vJj+4J35WW54rhXd48p91V50z6/ASiZPcA87DPTVYpRK7nfVidvoKbYhP2g/DmcKEdabHPlDGh+h
/ZrTsGez4INZ0UzteHJ9SwfUPSXCZ1GtN7eMkOtxrGYCkwRtXjGMXM9r92BvoAI5fR68DkXVkrFK
lhdnQOqMAhOaXYWcfvxjDWl8Nl37Gpjsh+Nbg81HJJg5blAaLo+Oy8M1Z2GRxuuRKRFJf53EqYA0
NvL/KKwNwJLswddT20miC54wAOqA82qDQtwod74kABbo+Lb0q/IbTm2Zuot1Q2Q/WKKuVUhs4o7c
ihzHwHqmsQS9KNLORcHv75xFVKpKriwhftBPiSr8ZxVOeISmfaNJBwliO3AphDdso4QXeyftIjOQ
+6WtfosGghhq6/tYkq86F5n8qtDCdNrKZjQaNC+GmXVNBDd3kKn0q6uw+0cQUXommudzydDBCLGu
bFfFdZwqojjhxEbpgKSLqE6TWfOYCkWP8QCdfrSiShPezW2F6iye0um1oSCgbfQKq7S9rMdzFHHR
cMGolP22hS8/Ty6Lm+K5wsd7VckCuSc415td7HNirAtOEyCBIcy5fSGyO8BEndxj+HdLL4NaMp8D
QAupECW30WSxdDeZIcDS/yXlM/zzITJAG0V+bXCKroggeQftChnloDpoPVYYnapFPjNIgyRdEdmb
GYKE+UzvMbwe4qShTNaYEtrYEJeML0x21NebeNSKS3x8BWilb3Of8n9l4YcU34WFN/Qt4/C9HLJP
T6Ql8qFHMDTSe0AM/bYt6WGOUhf0wHelkwFaCvF5aDhCwIP9ugpcB36GWIZm7JD9t7skxIaNxPCF
Jmzut7QEuLVAL9A5qgucX5nlTNOUoGF/IWHNRdKJubR2sDM7/lVQb0RXd4PD04bXFnBDatqNoi+D
zFnqtGvdUuoKhlHPQhalNwfBkPbz+/tYiSbDZOXCFIsXZMRWDhdyBmD03iIfBIgwtXzAGpShwVgz
4LTRlNcCegUY0O0Ic5axAY1wH+dY+lv3MEc0Wy45WoWjkigG5XBCtq63RxSy1P1Nz5CE907lu7w9
VrYb5dqCXLZjbnPrTjuLoU4v6Bk3DKXnNAzYjz989azoqP9VXoNQhVwEv3n+cg64vWSBdSZWZgI8
U1dUuC5VowHbSwB4L3oGReY16ISg+in2oJm5ip5g3InT1XQKfqf75gm45qiHFTwNIUv4/4PntZ9J
bOiiQgkURPjJezYVo6NdeaXR196j5iPBu0FHjSuQmWS3J07qydtPhn4H+H/UghmxvBaHh+8myKup
3kxTeg3q4gHPyrPNXZT18lDTRnPe+doslfFYl8AH9L/EgtPSMNO+bz/k6h7AzmpInBSsASIldo8V
Q1Ycl168sqytNzJNCB67sEuMnU7j5SA8Kv3yk+NlWsSn1YMxVCL7Irt4xDvzQXQ3tkXfwEzm0o/u
2r4fnhsgDmSOTPtjtBjWIoLE01LVXE2WxqYwiY7ZaG5uX4pskrQVIg5gLBSMPGp84qQKU04VKTwa
IudkYWjkGR7BTe8NJ4KJuwIkJist/E3osRmnVqgO4rsFJhBczlDyQE/ZTCh1Inh5/3xK3qlCxvZT
g7bqMzXdb9nfvWJltJl7H799QtBIAGYPps7vEM4lAlAgMd7UOZpBmB74y6JKEM/JzUkdGSEVqQvU
Ven/5joO1GNXdBIz+V1eebKnB6XpVRbhqDS/ykuNnox9ojfFvoJWK/27mcGKKnVn5zNHaXzcANV3
qKgsjOM0xcpxEoc8fdHcvn1T3bJbuMjWTIOgNzW0WKggupoHycgi95ZVy7CY6jodfBA+llX/G5yX
MIJH3ybFhBsbEiM8bD0Fo0MikO+Gvatxrjj3awpCeVUKyrOYHrjPfpCxc7CzbCrHI3MD+Fc65/UV
qjTpRJcdXnUW4T558XIFW5RiWKZBAzQYx0xegbGeTfFh2FKyQUX6bYZknRWDarwjk5lsRBK3KPHj
YZr2t6HE+0KhrmoSW2I2AEqlLagC+kV8DZLSZd6K7B2MV8XsCS4On4ANAsRQRZ3i/R0JGJouVZyf
nD/dT4iV0XU4Ns8T6RkNmadkBKT24Jqr3Gdv0aqwp9zHnnrcADtP+eAx2p1EUp5aYYXw/rVsEVT4
8z5+/3MF1yIsx9IXjG4+6yOcLct429wVcKKxTpvNnd8JMylK/brSqJB+bwqKkBMtWu9sf24CKvL8
T5qOpbj3ZYmnwm3EOtlLQg3NB1us2Smvi9D2KXgkPh1ILaqTgsTOJbgpv4Rqxbd7uoW7gcUhnO6Y
xevT/FXiSGF94Q/rRcuVvej9pBTsTjsk3wLXRPzz3pLO0KPqjhjDoVWCsITXdUzQ/4OEmgihQ56/
Bcl0ACxxDr35UuENL5MNwZPy5DwDChm+5fc9pxCAhBQqQYbxsmDlp77xkhTgTVRoVhPMq8v7Vl2E
nhHs85gpqlbiI3xG2fT9IXV4MwJ9BX7TdL4OxymslzmNEO2oDudtsA6yKtlziDRdcg4zMp2tqPaG
P3nvOUk6kh96yXkZzdD8oV2HyVB3/3cSchpMWPHi+/uy5XwvN5gu76uWrLISjVluEr+0X9Wne/ps
yYT7+/tYq66gdmqKlg+/WVQSr0hAY3auZduw07kBifPUA6LLeQuRzyPa2L6yP2bhfPs42tMOesK0
dcn/Vi2CbvmcrJChE4ugAssh58z6Qu9PLWAGOXtbQM1n7gUJpGNuFSgWquxeu8hdveTLzM/cLrUD
BAWz4EGHULSBueYJZoxrDQf/jv1RTpoTtruwvGw3wk3N4mxXdrtHDbq+dX7ja+1jmkt1xqr/BdvB
U47vO/G4ZcbJh0Oxq//vicp7xwM1H8ajhMjnB8xKeyJx20j0mcmX4lzFhuotiLfehBUqw/uCGIji
ElwRtqV2Yb4+MNk5nqrO6sguY8GO92NaTKl36N4h0IA5uG5AW0hpQkDxM6EgJtywxqe6UsgEWOyr
n1tl1BovmhB+35NPimicnYcBrJXdpKsExvOuEKBN94Q+XuUDDWhqi2SK8HGsV5NlcxCUQ55hOeyO
n7izWLKF2IHQIrCCCRjjSHSD6zr6xKmrzvDDLcZ7hOz86vwRXDlGLwesh7Du5cr5gJ7TSafWuVjo
2qdj9PKlTnUAe3JQTALhjKScy/sMvHDIOaQLOUqPeb4rX5E+eQrgk/nV2E9obUMaDBxCCPwZzIK+
JioA5XlhYREhuLmXfrOhYjo6OqBffArjU2DCfJaPKAG+DwmUunFzRYBg1UoA5yOMqQG6ThvEk0tb
Q6qD2iEMY7En5gUmzLTKBjYBsXyHjLdMKHWa5o5bFqwyQu+s0kd8Lxt50LqMp9CvLuG5oiIfMogq
037iE4aDT+hX5zgdwyceKalPxEyJugC4+e843fYxm0geCeoG5U7QZfSOWHQYTbVbJz8j81JdZG4S
FUHnWNRuvU4KWly0URaw+h1VfXHLuGDnribAufNqcM/nNk8tIvTievBAYI3lq7b3afTvdiyXocgr
VFTBF/2MzvRUhbgUSmE7taHIOI23CnrjrXvanLxfVOywmxq30xWbPXB66Mz019ryVl5yIDndLu3R
1RxuNJLoSsDN8+gtpbZrOuSLZPc+MuIydu4CLTtKCZC6lTC2yIqziGfijmtjkUK4HGwTENE4+zX5
fhZofDCMqW4sCrO6uAdtrQlvUopEOR6lZGfqehI4/3seyf/5nAEQ+dEJZR/VS6609tdVTpQajtTT
/0rRu3II2px//oEmNLYafOo4epQusTgi06EY7DhPgzyThuYcI6FH1IZ5sWEkwUrV1HwxCo9cOG0h
rXHxJTUYdG9cH7bLUE2ZGJHHmMc8Ps25scKta7JMBfHCuRc3lW4Meo8IVs3mCBL8ZwYlvM7eVpkB
oCYtlqlQGVtfgq4tSvReoqHHEBYC+l9P3zJWSL/ldSwvKErcfy6f8E1rEIgRhAXdhPck2GzPxly/
3034kq3mHiuEMVcq7f50sGy79olEggwo2/M5YuXDDhcHgBGqZRAFNawY7ZJ+vcPnqFVeD6QrXd7E
Dh1rTX+Ihf5opQEUWjRBG1g5XEv2f/jEGACPTotTKL+HUFbn4PhTtqH4rPEPWU8PyKLGjrTQRtFl
PBlZoSfie0PPXAANZNrjZAWH1AHbxJgN9V5nPJ1iEmLajTbb5C3vu3TVLXTqLvVL38mil5lkZjvS
aqW+b+VTxcAhWSYJ+I3egiHxYwNtPHuPPmzoGthhZ8IgQ/eDXhIkaQii2UY4RdvlVbjA+11epgkp
8C3eqfwrfutHyBUV0aap7rOsji0pqlPPOeakDRfriIagFHu9Z4A7WY+fRUxCgjbGDf/+qhGxSW8e
yxpaEuy9jp0RL7m5nimy8pkCTE0yoP+KKhcwjL0gjEPf80tcuFztrD7Rf7jx8z37oRzlXMNAWPp3
Kx69rXVYyFDoW9m/xbFpZAT2V+sFiUqdlgO0VlEUV/uFZpm9Ki+sCdA4bP6+bveO5dQZ5S1bCq4/
Jtz3+E+ArqleU0WmvD1rJHxgY7mBI96Fo0Zd/5gGaxvr9VKl3rCUtdRun5Npjv9STcNgi1jRrv+B
nKTq94Z8daq+uZIZ4JWw8G08lfwnF5rxowSgKXyEUovRkV41AU7qDuBL0M/bV2qGAmrOVhLGuihT
Xuse8N7ASVAjy/NrPa6G3PSAGGaDaPGBsW/+bnpufA5La5epvkeuQfu6hGFFo36hMRlP3JiaYHTm
2yspCBxBWcFaOGCbkpwa2473fGBcjNGtw+zcL1rVGgNhAyatq7TO7R5yIdd6h/b5gLILqpQDPKIY
57GJfLqFa0VvC0YDMel5BVGkcqjsGvPX+HiPCC4ORaIl+My4iG0UZZGZntZv3+xQaagvL9OJd9pk
Itp/CaT41F5yNulXJJ9aRievFQZc3+TgH3GS95DtASZPkSdmsCADQUiy30s2lTt/QLlNi0rcAQQL
Y+Hq0b4bKhx61zwGU2QSL4miF7VwBhyNK9AD7qv/jjvJXSMWF3pgVxz2VM07MBySp9Kn9mbauH/c
Mkl+XOUsmDx1ZpXG9yPiEcIIrGYWU5FZX15h0zUkLuS7pyvD/EUPAiAt9leyx5M0KUtssA84GYdG
04y+0gl0nsjbvM9FoppZVKQwbEZXOb3FI6kgPFmWrymFrECkv3hwV9q5C1JQD5dzbKCYGz0lBwD+
gTVEia9hjyrOARTrzPyKKjPzZzCvWsvsMaHSukW2tA+PSKmSbJyxaRVeDbVBLsZMlF1ZmGlI+jrU
3V9Ks1GCICGfX1vtbppAOEKFzQwlUnsVIgnU9+RfKFUg47zh082VpOdP1McBB2LqHnGMaVaK9oZ7
bFng/xJhOhsPlHWPWncUafNAqpKdmvNHy3kjOhVAMPaARxG7wnFd7mK5xPMnAQpxBDV2e5zWuW9N
KgMHNNC3dEvOB2tSh7oM9fzhDo/aWc1UJ/bnmv11tC+Iwsf6OJ1lf+ruRuJI3Y1EZRTkIPgOn3b9
e2frHiZzKE4KHr8suA9Y1UrKfy1JGG9QqLFElvXaOmrp5FBvTCHzMJ/68STMELiCrMwWb8qpgj29
Jep7drspVkmXhdPZ2kHfFrpigFGsfXhHv/za5lmzNJeAS3emtcz/YJIJpaI12kY7NMH9KaQpyel/
2nqoEfJ9LJzZ4fUnp14Wp8x11XEzd/aE/k63V0GODcaLuzMp2Je/BssJeWW47k/G/HCyxZ0PvHYV
45x8ErGcjjel9Q9yoagHqYqDiSNkvNNOyEebUL0iGsUSnr6KECkEERJi643XyVvvG9DPh3gpPrR5
Kq4rD12r/h69NuG1OE5SldtIu6WAYPIBVwlSg023Ktv/ms9fpWuQaSyftPRzJvN+PdQZXg6p7sWe
u+K+BXjRY4UAV7S4TTNI4RTK0Vh6b9+6SIkN45O3HjbyibbZpHUPu/kbhb9opE3k6/6UvB3jNGTB
uUQhVIOlbtHiJZeEvsMke9cjdy4st/iyP2/H5joD4R9u8FR69mj0Fv7abS75+ibpoYqiVZSkYueT
Q8FIlW0YOHPgmfd6NQy01TpW6nimqybxq3e+apExEFJWJWdV8l8FYsPIEWuXuCNCtV3rcy89Z3lc
FYGwVYeQYyKUVzhRnq9C5Ni1PPdZClwuvR83v00+rPtNW+J+Dk12TqoCGKfwLMrLI2sJloPh7xsu
wX8Qx+Lf2s4MkQNyIYUh1dEnf1JeDR2lP8/J+ozcC8dEaA6zfrUPw4b38+raxzFiHKes2PxkFIwE
wNGx7eSND9xl2Pt1eX+ftHy8gSQMUJ4eh53MfIy4/dHpGKZByvANwrMLEdrdUUxEqMoQE2oAKp/y
YX8TVrpvrvvgQB+71jOegI7HND4EU4vPces9XdcTpqwbfl/uXlIg7qEUCPnL3qbtV4BIzw23h0g2
Tn7cC1G0hHTWK8TLaCpcVvUNLYXL5m8XalYgLTHNVbg0mKQ0aFUy8YQAfB0KuAeLRmbeBHcCvAKj
KZCxGDuMNxLtiiw9BuVqPLkLapSQffJZv0v3rcsGzr6zOd1qsidtZiSpdcC6DoKcVO6cdgP+ierZ
qyYi5tAcJUVL7K80EjwcCeR0llNAG+slw7VTMWDMavSEnMo4ZI5mu5ea0XwTvuAgnOd8qNriozv0
aJWGryb4OPlCryjWCaN1t7QDVU5Jogw8ISlwyIMPhzHN36gdgATNe/k1H7u3EHorC4bXApCMKpRJ
eVyRGGuWC1VgMYdTR2lLgErW0n6l5VOCNZdpt5ZO++sAqxNIrHfP/drbZXf2hX53ewZdGFZ8RV74
l1c3hpwEH8zfss5aGUqRCuk0F1ECUtNycmEkz/UzJ664pRWgh1AF1Czux8t9uEULz3CFS/YHHnuD
nHAzHMHR2ofUBFfdKQcp8fewUqSZGfte1nqM7IIVs8MzL1RFZAtxNIISbnGxNgK4veocdP9Q6fTI
5rdE9jv/9fIYoVZKRpdmBfz6O/DtI/hyiaXKpmkb11eYI7pzBYdq3mOmXSp8EkGVdQ/R64ZtViKf
L0kPhVKimCzc2G6OQJd09NROwHcvNUP2SYY8m0CIOKwzbCUejOxq0xL+LbOPSDcWDmYr8WGgnadd
nJJwozZhSXtoVYazRfebSYql/+6hCuc462kIXNo6GExIEHpfoQbWDNmPLEBeuH8efun9/sRwNXno
25xcvHVoDEFx2DRAwyS8/LbK/sSgcK2attFU1NOlLPtL2ZwG9go83aDqnEm0SJmwWz4sE0s7FhqM
AEK22/MgLqwymdNIbm/g/i/rCKnN6AmqfCiZfy1xQNpAYi5UPHEZucwpAPX04vesvdyTgVo3hTrx
Wy1fyOK+GvGgRZTgcFK2oaYDMDFSm/fuUOH5MseOLFULLgdWpu0H/JCZcM2+F8evWgYjEmctIoY/
qJbn+xwJqlV4ZHPQQarPVk+ZTDqiTsjvvvxNfFfIYrofED3xKqlpM5ECy7107pYxoSFzKeX1RBNH
TV7W0TohL98vH7uIuZ+udln/Zvozgej11Ju6DAggoqudRvm0F5COEXOrAzMU//RfIoSTnx9DEbe1
pgd823tIqnYeGrau1Ag3XbJz456q1TFTVEE2GwDmaHo2bj4WsQHgiIcwYN9Qs2vZo7RoIkPKFcrG
FO12slU5XrCqBx9qXRlZff7/ATf9tFvAeyxFoRit4D+S8ceyUDF+/l1dPSZbS1GyPeBXHUDlNbg8
3NPXDXAZabvQ6jaUj5YWoLP4uicpCSJNYWMefvFICbKxaHFcQ5XjYN2asFdinxewHC0AZE9QysZG
li6i1e8FkADxilcAP77haqQykJFV8a34/Qo1dOF3pDwhK2U57n7W4yxXX3+2rYwn6UvoLRpqzUFs
6xAAP7o45P2c4QcZ3Sg5nOxKDB8d/oLUn2AImlVvtiX6XkT3GExgBtZbkGwEqCGB9qNMyywvKVRG
OdDzLx1bL4+raTpVc+AGelXAen0ffQYh6xQidvUvpEhcXOnlPbLSGsuMrCidMj/LBPAW5je4RNDw
aV7EK0/BtzyLwYB9zeFNuG1ZsF/lUNVRlf+LGQIJDedSFpwY4QRXlHuBQS1kl5kNXc/bK40wk3dl
dDEKTAhklzav1ERYv7OSlIDcQ3xbPjYNdtFT6LvlL/K0TwTX7VtHLpZuTTIvTo4PYRB2M5HWjKE7
YOyUcLTTtG+qZVV5T3U+NtwZYrtM09Efa+o5enJAYyo8W7nYI5YtccuuGqJ839/UsO1gYkt7t9Fa
iHvd9LPi2VKhLv9pP+caF9oTjAl1cw+2SQdVuQKUXa0y3k9RNOyohICnFiBdJhMiUwD1+WIFRr/w
KMNtoJWdq2UHG5Cckmhouc48KI+rTqF/s8LVzZ6YWtiVPSg7wWc5fS2mdtVOksrcA29BQcLcHRjF
HgGxkEu6cJK01Qsvz1R/QQMwRN4esspK8J+giGBMbPUco/EueMo+/s6jMQQbJh8IQwhhWTf/k0x7
tgQEj3YdKAjkVptywmi9biFzTjEYyFO5FvV5RV+LjhbB5TWcsG6NdaKpuIdwhQ0ijU0YyjAAK9Su
7JXYw/XsIYZzHuYlCOnijzGuAzb7X48VNZg/OZzfmgKkhiYitOCTNpPoOoDGfaCmjj0gvSHAfN10
R8dOOzNGt68MMyhWqSqVyB6Crf4DuPdD5CEAI9Guokt5WMjflcZ9ieYpEH6AoaR+vcHkUlsrFTtt
Z/5GF4ih44xnKoDVNf1wx+3Dokr8GGWo0h1aprbxK+XT7d10uhNeD01PV4xET46cRzS5Or8TclHL
m8o5chEzQvxl5ZlsrMFINC5HGar/zc+th+NkHQCD6aemw4BBO50yQDr2HMkmDLZyICSr+nukGgVU
OqqC4khrRJ6lX3wwzjR4apmW2KD9qeJhNaQMcx6N79dRCHex/nAQQ1LJ4nEp1ALM4sbQAamkR3iY
5T+sGPBj3G87CXv4+NNDerGxoSO5xO4ZAmCgGDBE4zQOrNRbU30e3Qi2ASeYGNwV61RD4AZjxvzh
sBXt05vVUr+YJhJuWhsEIKsKF099cw9iyQt9EVBeZ5/pJprAY11IDoAVdClCnlYfc3YM1j//FbHa
Nd0iWUxYhyLituKwD2GUxct0GCEhKr21Q1/eJQkhjssvNx3q7rp/KtLWCJGf+dSelWz5t4nxKPof
SR7iWlU/7mfgUy21uCgaa/U/utSP/FKoBUwcudDxTe2LDKOf+ffu22FC9tJCDSLkDVtBFWTu7wYY
gG8p7c+IG3rqFsrGiURz4ksCr89XmGBj+K4/wtPoSrr/fY9ddQy+Pj+0pJxlYP6QNIlQs8GpYpZE
6fSJiYAWiUCEtLyb/18KDX9ZvAs7p3lfLhaY6b6g0y4qGXm0mOshV/EXkFbbaKJWX2V6D/X2j1vd
c+FD/kRJxCRvxwcQcaE9Bhrvq+rmVr5T36Fh1jZUNtWSZjDaCii91ddTvJCYZTL7o07IaXIOJ2R/
7xgub+ee9H7QRCd7DBg9DoDVToyICa3t1+bhiCxukMRBL3sFnV1MLJw8Fwky/Ofkg9puWbOX1pDs
RRHs70wwwpUjCX/UCPRDotdI8cFWHHilwTaDyGE/pX4xVwOga5qqjzE+3uftzJI24ih/aXsNejo0
x3uI/fZbvmYQutkurBrWgqeh5X7iABV5JbTj7f/jjWJvWkuvSMAR1Lg8pS0phWmJ0KJTE/7HGgGL
EyIutbUwrvAZF5y6y7NttI+ECg/NqJhQ0syK7PRtBWt2uvuLbVdK6itMd8YNtB4ZHvd6yKaoXkvx
0euI2mssalEYNHvKbJcxyk+c19hgpvp3ghRvkDwWcDzatAWfRJYm3Ze8iPfpftW/e6mm8zkx36nK
1yRZKOV8apxoFY/vNJxkwWbavf3DvQ1qIKsxlSCZZc8sxL6X59Q1uwpm6Gom1PmseFgfS+kcUOC5
o4YrSvYAsz4SpnLDuuhWUREC520EIa5nRE9vRwnKlUMEUZfP2Ne3gk9tKAkMl2whmy/NisB1tYjU
7R9c6UNGZDrerKvZtvIWQeUfSnLtTTJZykMb4lRYTP5VUNel4wmLatQd5JouWrwnaOf/rilclpPo
mMXaQkcAquNdj8TQROsy4WBdVQYy32nITelsOWp9vAlzx26M+xDQcMz9B9LbwzLdnJsyzNQRk/HY
+lVPjmfrWsoiqB3ElDy9hy9VMarqMNRtTXhVDHxyYrK8pBTcBEI2ncI0Ljk46fwKsuS753lXG6I0
Ao3qRcRif206EoPjpa9gz5JUJuQZFl+B9D9W1B0UZsoiZGZntKjtC6rtNr41ieneOA3NAiQLTjWk
kqWtrG9HTLwYmPLC01DcBiSWd93/luyuliwqQoVo8X1+tlA/6tyhYwbcWJa2hNSx3WHWZtFYzY2L
JfJ4FbZE5t3Eba7wOmOiXq37uNxnNFxrRaR3+NBPUiczILSHKiC+6Wsj3b5ONdMCXIO6Kq8WzkeA
6UVBFGXR5PtI2/rIGpcVZAlxLBDDzXwTNFYW64vl8K0kyL9gbTzjxfEF6SbSt3MW3dRcOPLgm2tf
0nqjU9Hi1iZHFame4RD1zQI4wSuO6joAEnZW/d0Di+wdF4hpatMUFQkzqMMsCn3XaCh+GQDdIyDo
paOTL8Vw8Nm0gJurbspXcFx8NdrXINlDOp5ZwLmdpvYYz21WacvbpSbajqJaUTu2Csu8Pe3Xeilg
hehYpuO7JWbwcm1igX067hZnC84dJNDAUVhePQZbq31TDi7ice1uAajpD50C1S0kiuR9Hw12wiPM
jwBprc+iNARIDZNErHCXCz/pql5qc6ut/a/2texv1iGBdt5ijUbsCiwr3OE6A9nN6e33UoUKGPtj
TjAph5C+tPUa0cGlAXyj5RYJVU3/d7PWS6QtrJHSfzPpON3F51bSV+nELDOLcS8UYaw0np0O9iZm
X2W35azXpDujpZUnn/sXlOItmEPqfAyy7pg7y6Oof8uSi5lukmxnqSWiOemLSsGkJosmdO+amzzn
9b4SYWVnaU2+XhbvNfHYur3kCpQHwWIBwGcR2V89awM8Ni+QDn21N0zbL8GtfNq+LhUEOIABpu/N
UgVB52y9Yq3XhQm/FDsDlBzX7IAFrdtaiBl2T2hJeWaG5ThVQSrWp5tqIjmcNgRK3u69NdJ9P5Tg
ggqeUtMJj1joIzHojr8MzPXJchdkAIwcuR1Doz0DaL3C67OlXifI9x0H022E+KCpXce3ct9fXNGW
R6c0EJaBC1pZxG99wlGrdDc1oM8WrRzyv2BgNbhVq7ydCM3jiBrywqhM3HXukaKBY9SZm0GlpSaE
8HIttCPop+3svySb+Rw5cGHvWId4eSw1rx197JVYyihb7OS9/nXl7p5yRgsRDJOTWp1c0DS1qD18
NEVrPk5tHgjL0lDwg0ycm9aU1w2C6G5Etxv/UlUJQJMbQ0OeQz74qcTh0TnY5JOGJ3qz0m/J1SDs
mE197eFj6adsM0I1YyD5cV+PcQLNMgUKp2tYyAY4/z35nVAy+SQ2AAcH/DNqNOY6yCfv3Jo7J4rX
h4I13g7ui86+1mVcfXum8nLIo765rHYssGBJRsXtlEH1si4dcwKHN9fUfeT0jyaizfJt/sS60chs
+nqzVimOvwqriuRfOthZ1sfLsUr0h1m5jCUUM0jjXpfdI9ErbRnHiQ+Ef+MHaJ9ZBLN2KNqfnjpa
tiM72ZwRmxJipkM9FH9JFT7CRqM4B0SJPsugEfwfjMNEF5mCVhwTzW5jBBXJnrZQ3biAYjUKf0NS
NuVAYamSCeFfbTZm6gvK8q9YBFFSU6h8NbrWi9X29cCXop0YFv5wW9SLnuiyz4OihFfPlvc8vloJ
lF2JaFtO+yBhKrUYlW/9P3a8zNj+nUgrbOKb7SOfps2j2rj9IaqnwJ2gQuy2USBYFJ+RumZcMt8N
QJswa3Na41akrGzDLS57kZcqSXRl9nPtUsu/0hyTU9hdRNkQ88BS6cTrw7GnXjzhHJTQdBM1uiK3
/yz+sESq0eLKQrcklO1t8RNgwWD8e1c/WF+AjCAZ+vKhWtij3bEGvDf5/B11Jfx84DsbDP9i1X8C
CHqUAwO/EshLztGV/xTHla1GYUuaELqTBM3wx6b/p415qcy4US+wmPrrgv5GmssP6W84GdZtJk1M
+LoqUayBqvlkIxSlL+1EJtpfbluZIdOoUVkuJK5RkDMKNuX/MYIti2U+dwTNn3cy5KIZvlX+Up9c
91SRnNRHi5o9poOIcP6tGNF95bfiOV6i7Xyx82ffL2lBiYGM+BXChjSee8acC9O2H53SwO4mq68e
TPRZHldJtaNFe9EJ3DO73OERHOXUEjsJixJ9f8jrmTCdAS1P39Xlcp8y2hPNstnpFRF2RHbu0MBw
8mFttMB4xHc9+eiy/uwMZ5HTnp2hjRxRSnXH0LKplaeTeYtgPoQYnGvUcnXOW56XKA28jpSKztyG
xMRwfGpkNDhvRw03bqUJqRGQf7Bo/vCVGYD1vJ1DJggKhEMBxjndgbmzSNf1Cxm1bgjkPuZCR/0l
4diDWp2KoDUGB5VkVt2mY45i4DEAnm/St1AvOGEbqS+WWeH2P2Sc/Z5dVmWsyDlWqrYF5DX1wO5t
q/iYDMuU9nCddKKlyehtnoCh2w+cHvExyOVAoz/BXwZolQftFFz2e2irQWjo00ZitO2fyvH+GIDM
gxNmioEoEKGSRk7aOAwJXUkGk4UL6mP4vMZaDxEDkk9X8bi3Jebqxotx31dzGjBRgd7mdebIQVOt
rfk1E3D3h2GCrMAdTApf3CrnE6yg1hjk3AIOGZ9aVKP/x0WPrqIR5sAdkLfkemIrVQrZuQKCrsnO
AJoFzG5uwSIIHFCu4BdlDkGdM9Xzi6VGdaRmD0vBSb7GjYQHl3qO/VkyfiHkX2zRH4KrcGcX0uhK
ZxnMKQHrMEM9ICKkIbAhLPJ3jcolXaQYWK9ddW5oIp9zg/8xMPLFLshjBfG25uxVPrJqApkA9hO3
/yHtQBkW0/ca3KiKG5EMaHV4tuOqGDfu0vGbSNo/LIcKCcF5LnnJ2yrb7j1ArrxQWSlGgQX95Um9
KMFTtM1LO8INZ0ZmAzcwyB8n0jS/22XDIyuqSaNa2lOjsg/Fi6cEufX6h+QKp18xtd1AFq3z/Bss
JudsJI8tfCdkwtx/lXVemFEexBOp4e0U0M1laYWqwzr0Jinc5G8fY+k3I6sXYNHOiT8vs1c7cWBU
f1EaLc8Sz2gjpWC7W8Mmu5UkYhIwbmfw9ShJI7nCRUg8ZVv2zi23U7J1bTm6dmRxxivghc91YT+H
Xl2Dx9c43NFDBlVj+R/SVIeY5pFVgvGMjrQ4TIFKDT8KMwu0d8DMAiof7nmHasV6gtn4e5jkl2IE
htwksqjPA9YMA512u+QtmsObOcyRa2A99d0NyRPc5QqfBaQ8LR4eAgBUskzY+18isQugmIF0hkzm
m/zk2CbOkHvSqJ3WaBwHe5ZGBOoeEAAkqnxsxbicGu/v3JYXIMl9OsxAoaHkah9rEKAapcieFmlu
7yJsinsdoMEyrQkSXln6FhtLDTxjBcWHCdN4FesLR+kkv08aRpwv/9/hEoglTzkvKTsTHrCGDJei
ujMbqOcmG7+xhUhLjxtIR3R65fREg+FPALAaomwS345JT1Zb3HW81+mwUiFqzkK20oW5s7dNQ6KH
6AQBsxurGaNW+ewj4RoluPxhz1nUnySU1PFyMd9o4mY2tOIJZ8cpUH4c7IWnJ+rPt8NkRS4fVKLm
XzMxAxJlyBJQox8fQTewAMnWZ4rztGVFB4F7irvsiMZ7uXxCjjmO8Nv0kBSfqFX/f1c6Lw/tLp8M
M9Mj5Gj4kunYMyIsqxWzHGm5I87rAwtw+zOQS+cY42YcXXJBtFahdeGgGzgF2pdr9nH6A9nu+4+J
9wu3nCAGwFZOyB82l/PtuykpBDO3uaKYHW4o+gh9SSahAbMCQHgK8002CE0Q3LT7EQg+4kbi98em
Eq/nla2vArkrKdAKFekIsbRF3LmQfdnCAIpoU0LlfX52KFTb4frpaD7QDWIrOn0RIxooCOeRRFxx
Nrl3o0TeCYWMbnc4ydOkn71d6ZnCssVjFhNZVNQy9uJ55bym6GwnlL7LbcFDmTUtu5CLlGG7I0hX
HymTEg7S/omQtyk3Yhbd3QWT3L9hEXBXIYeoiA+tKLNJKl9Nm5i003pJpRIZapAkFwbNSqNCnt2l
DJJjBsuV2LjmiqH58tzHCx5LRJsgej6zwod1NneYAuKZQB2x/WLD8S1opm0bVfOBCV5n20t4opFe
4USyVASKhgZwms0Wm4Yffd7o8kI47cnJqR/FlWp5eVW2fmqTts0N2OM1J3pUjo6n1SS/sX6hPL3J
HOlA+vS8CMSv9YNKUzWQ09f9OSw5VdTXTu5MO21AIdhHiIxXD9uL8dnE1iipCZvJbljm1KEbLViZ
7+0fOfMHzOzw78lan9775Tiewgz5M18zqxbxH9xD8Nhu6MtUPmGyfSLewQzRlVHGklR1OEpotZVq
LjXNJmJbMqRWi+fS4RPKJx7xu1EXJhdBcAjbyZdF3f18PcJK7UsNDKyWHzFwAwlddperN9aStpgY
Tmnmk1AmSEFP/RKZx9O5V01pef2nA13IjfJVjEcmJ/42/hJ4eObEEsvSC41eHOjEpoPElmiKHOvE
MW/JKwYTDC9k0pM4IrwGRUoTjI2GsONiPJzRV/+k7z4EQItkbGnnBC0hQLM+wySVsXS1x4sIK2ht
mqNRfvgw7h849gXgo3fJgI4AephM2goP/3mu8jhPBu5nBmmLPYqCgqVHYqGxOEEPPSjua5suQc1S
UvuA3CD3eqr4xn7Bgw27zwxJQLO06T9mBPNKDtF87Knm4bMPew1+2IJ/CmGiDSLmcyc8WBS+fPlF
/niJmb7NHc74sCu+yXnGHTC8DRMbh5Vj+hlFNlO32vFMblYSlaubpYa7Cl/AErPyAbbJIeTJctKN
0F4hJTbBPXNMMJpX6hQGej5vm0xhxq/c9yp1xhwuXBwjotKk9l3OOQhovaJ9suhWY3IK0LdOGmwR
2dZUfcYitNdrSeUrfoqABE7/aadlbEM05b3ZZyMpmnGI1v9/JSqLbt0Qlpu4lnXkpEo9Xc/sou63
Tb9GJkUTCJ02Ei4gi3ESiCayG56NM7fBwzHog3C2P5dRwfdGeuxYKAUIkxxf1URjoQSJxkNkQdPj
5SclaB1wAyROIr8FOTh+zl/zrHp94r1270oovdCtqVLPU57Qf5FO7C/i2mg3dduYOOvno8Swm3yo
v/x1zgc7AgXyda03Dlj9qPOlaIN3E7dMGimEH+ujoYTLvKKSus+4Tt0FZMoBzSOifTjG/GQf2+OZ
X0UjF2Qge1NtzdRldQNNiQqPJBXoj1KniieIK0o7Yx4RxYAJhoyJ8Bx0NFVzrXXtMgms7hpZD0Zx
PQpFaoOSg7wI9RRHE7tJhOI79Lk2NNe05Lx9jhWFaqC9uZDolkKxLX48zC5UcsNEikABTOL4Lkzr
RD3ijgnNkIZUSGcQTRezP5bFgZp/WUq+mFNZuTebEl7uVSZFp8GeiXGZ78IMx+Y1UQaE1G1kk7IK
uTF++7jJGIG57UfSCPNinWCEM4FjdORqDH+n/HdUwXL+JWL9eqwNz6sjDJ96znvIVBR+gsZ0DTw4
2lCEdsTtCHH8Xol4z/k2r/j3MeyWfQ/8lrUVPfBqSHemOv1MMoeIKLnifgVW785lLkbkM+FYmKmG
lUjrHRuzDJaPU46aYKQ2fJ5zPSN9hIhPS8UON0M+3g9xNmRTDpaNgI3UHm1cR2tNylTQRKJho9OT
jleuGOxYCP05R915+7bjrHC3t3fkcevWOq7guaF9pN/Q1hEOP3NdcgQX+hRbSMst0THma12+xCwA
Ojz/tYBTA/teVJaiRg4u/EHJ5JFaUNg6NNZ19PfIYHnMwTCWFqFOyY33qzuBSTwbHDh6CBduEOUO
s1ljVePLnGmIkU8gemaIyikcyxiaydd8SNJArhPKyeKsyVAHy5+Yh6C1dF3jfvSPREEgLSoczPE0
mMaeD7Ydol9L4E9tbTMaRwi8vt4mscc/cuwqjq4mvuFXtGewmgWCVedF0rrMz37Jy77JU1O0csCf
XSryGL6Kmrl22scaeUM7zBKjhZp0bLCt1Gl724Jc/9mfTQ/wBbIBU9IkWUFjGQdO0X47EqoOLxOx
YFGRiiShelUGH4V0iHvrefu5AfzYhJWfP4lsUXbk8cdGXIWEaYkcGTg9CwTg5uax4Jlhy8ajA+z2
zjRdTZZqqO4Sc5gq3pd48OLH7XOsN9yN6VmVGUWcS+afVvpUe4eYxx/KjTTnTJVhcqkbG3ME6Q/s
BYkJOpa8gEknzPrqNe65XsSxaTgPykIsj1cnUUzhbxMhiImhNj5jlZZpSo5H6hzg6l6/kwTw3N1+
YsY/J+0shZm1Ztb3oCPp8frEMCokfdGb9k3Cu3A/jve64nRTwX410bNspkTG4GVzNOrp+3yUE1Oy
FmT1qRqa2JXP8Uo1dzl/S5d3PhDpHqN1HFdLiw3VOGuy5Fk16RBocm1AgcCAlHEgJ/4lF/vgb+7s
P8wd6OaOb1QRWDhIPMvk1AUPoV9F7y2ztacbeYr8xmEUAvn4/JstGuBm3B5FQ+Pwzuf1oHvxEyMp
neKg64sSwNrwms3CdZ1jZ15d+Tc3/5Ww9emQ85P/ixk0dyjqLnii6rPBDFmMKCdai1RLBB9Jd9Xt
OmAn1pDVaDCWqrBCGkLaOw9pfXcRG8jzqHEO6keWCih5WulHCtO/5tgAsrXPwejSt7iZp9A6VLVv
fx/jQ4rTKRejgJHA+TWf5BvU6md26X4xAlfLQ3m5LQSw8HFXQ+uEn2fZ+BSWLezcDWW3SMHV3dFd
W3tQDWSIaGaqVw2ZIiu8uL1wLrQb/a4nZnLuE6EFS+4od5z9Y85FJgUWR/EnVrC65WWdvykKRjPX
84L9LY62Zd+BXiE4BlF0X1it09M8r6HwTNlXyQY79Woj22xVM2P5aiV3AiBaqEhQmUgZUh2v5JPe
fA/byojTS8ottLNUfPWwsbZeQRchroZ3GQCESxfEL+DTrNO4lIRkPj/BjU/7QGo9cEGMWigq+onh
4l4JlKLu/llErIAGzRJQJTjgXz4v5s0vZ/TYnu6qGbu8vMofGbkFrjz1xJuGpZj6GoMko8Xdb4h+
5QDaG5E+RMWG4cUiQbjP3Qnvw4xn2q8LUgzZYNdisNp+QDXwOrF8CY0v98eFDLDWbnBdR/lKQoQ6
NVnowhMSSYcX/KjlT2C99uniH1x5/Mf18n9fSh2s5EQgg9GFQNaV8w72UCSbV5cWHUzIRAfx5B9j
U5rlZ+3GUaLzqLM6hbwYYNrVckIwAFdOxUbPLRBHo1nVg7EeUd6rRe7zL9uJhCsfAvVPPS5fNGbD
HHUTy2yVcxq9Z8xr7zHayP98+gz5B58o57lYrTWpYGf6IcKCucsfvLd0IZeYDOxNi70hKAlBWJmy
UAyyohutF5Re+GqUSr7Rsx9SAIwTo26iL3lgoubGB6yoA+ANghDcG2/EEg4UM7/paoRNzm9y0pDj
tNGVD0aLoR7MoJjLD6LUyfxCavCJ1t6FwiYvCdRXgzso/rLGbZDpaTUPvfS9lAdCjSLXhwFOvWnK
TuRMHlVJ3taugG6J4ZCgbmnJTHphUSqsYLQ70uyEQXFVXEGSiCOG4SsxdDYHgMKMVi1slufv/2T5
nxrEAR6IBlpVpwN/wcBfRDuib3SLMNPVkFmywefm6yfdWuOio9yIhAK2sMr52LunaofN76x4eFVH
JROkC1zQ6u72pSqMh5ejFvOsjrrq/Vg4BCPkt5Y7OKdIiG+5QRc3mhZB24sXdyZxz2DlWMizC6BX
X3TKjKCiZDnqaXNS7T+mBY1hrDTOzaCAJRTGkvUV/TxHbHQHcAfYXpM5yBt/OBfbV6cLklItFoN+
LTdE2e8ntMOivCtky/4kyITJpwz/ua1vnhaxyY0Re5/FdvOEUq2FHh6NmQXQbH8blaGE4sp13h1I
uSea8t55PqBEyfifmHjpN3p3N8whAhTbF3hZtkDD4RtkDautcnXGahJuEntYLXIdfZw+tVbvAVQq
6Tflh29P4ZrzZLs7wTXzBRUcqz1DYOBQHWfH7wHcvbk0NUd6h6aoXSZ+LaMcybzdS/9xto66545X
galXap32SoWl75uVWElwWDe/M/OIca/RvOa5rAZ7vVnRP3g+Q/wgYpvAXnINiBQZFsfdTxRK2FBW
YqXstMNArkrUMU/IrOcy7tl7zz2iF+S00R9nyf6eAKQKbNiuaoE81NKK7AXO1i7t2Zc2MeMm5K5I
4LB4/tfTCqPzKX4SuGZK9JD6YDeXNLi72gaZv5i/ONdvhpsGOVxPGfI/t84CFx2AXi45fIQV2hsC
u9KKxMwvdjnfMzlXyE6dhLZYotOnJD22k02eIHCOMkWrt8t2UorulUkdN8gfQaqpstnAVp/1jKet
/ge/t5o+f8LGTMhXdTlCCH9GPKbL54zlVInUmJscsvJuRMSp6n74bxJ8BjzU3zsUdoz0ekXkidN9
gH7ogOp4DYWf+uJyyTm+NUtFbb2hgcCRUv3xNYbE1fBGl0l6AIpYkH1ZyAJuf+WRzkr00Xvq0Yrs
ObRCF+a9DAh052Ma34a7dezaIkQF9+Tj9ytbiMk2Z5wqy1RxqsFLZ5KiDM4KCVEv3GEAfGN/Aq9R
TBO4SszXNvmDbimByPS6T1aij51pANU0tZtKHZOifG7sMBocD1Lp4Z1MZskvqNXjuSDwET/4pfy3
IzrkaJa2DG0QqNKTOfAbeoBVSPhQPAlYRFx1imqTl9IYsSbq+0jQgrCFhirStrztRY3K+Py6xhBG
GCifW8sIX0XN5cIWPB0y9bT6w2j5LzT0qPg1hm0NhyLBCxScy91idni/S01BUy0uOcXjy+8h0XUJ
SEliUZhQRJRuOvYCpkvUBpPIajUioYwsHKzdY4yPhrOkqzSEI0tYqc8HNXpUWHor8b6f/W77GIsR
bPbOqK7U1cMMABOD9KWpE4BWEGv8ZbwtmL2p/4SyvpipMMm6vZBefQG8B7g7tAQQrwSguH4eClbb
0pEb0097T0elCpPsarJvHDCPu3z5gi+eFqwzCeA7Rk+N7tvJVzyRsi0aSxycunWuhBi4yWjqBOLl
wRCpyMjTOso4tRaqjGytU2RYXCV3RPkZs3mpvBGc8crKvJj+5X76/NnVBuxOCOMu/C4LKkIaGl/B
Ln8hSh73ML8wp5WtrnHYA7s3Y9dwS4rykpWCEVghG5tpsY5uOLEPnxfUCJHJa9+aoNnUXbldD+VD
yap9O3y4igYYk1RTNSbydccQ/J4lOhX9oDaa5BXTKWekvAPwtdVfBs4oegFqyOzItNpnFymbRuw/
N54jufp43vqHyjjCQudSaY7a2f/J+3uwSBIou2RWHmPH9/RnsJwBY01zv4T0T8EyCJuru7tNgktD
/uRrk/Q8D9ywvl+A4Q4jaDpOmRmmW2o+gDP1D89C/q9GkvcJkfDm38jvviTXDrniG26X3jw01LoM
HMZrvOh4NCfe1DjR9GfdbBEV2Ucaffq17rWiioK5DGVkcmNuWtb3/xz0Bul1yGZZ/gejDqYBxfNU
tyXOjWtBHD6bJ8eAkbsZJ/A1k9KTSbioI6bgL4Hc+CiuMQ3fy7tuRaBEIOvTd5ilpZDDG9yNYPjI
sKFw8CunYVjU1BtteteE2XObSy7jCoIrTedypzqLLmqLQk9gYVQ+Mv0uveAbgSyZ6DENzJMlcRva
avjYdoEWwDzC2XVd1ZQFY7NwoqR9fXtvcC8HXQEku9iE3ofjBqZcEAMCwHFqjmO3CFIy91ZE4N+b
95UQxvYG7jyyvR/+HRV4QeT2Tjb7M5/Rzgy3Dy1RaiUiaWBV8Yk0Z/TeNY+uVvSQNVvvSpHYZqpF
92338wjxDha34Rss/5u4W7/3EorXgu55O4CqFeZa5cp51/1iSAl6WNJq4MOogRQepJensI20FcA7
bTWYuz5BgeqOAZBzDY0WKlnJp4ZQppHoC7S2FpCDdze6+ZPj43C9RcY8SabN1MBlAT+pKE4zKuh1
4Nanmk/rXAHMGktnBJk5LKzscHzglfIXIglkx3P+47UsZnjYjV+1fpgFL9fMaXUHIzn+xy96/q3l
8pYBMAQRN7uCLo2vJJ4GiwHDaJ9YI4qG1XSR2ogLdzbWWy49IzBvUoYNXfL8sE/RUDkuaU1gjGet
u88nslfUWbGVCEJowhNz737eAKM/fhvnH6iEkGBfyQ/3OzMkM2PYzaKDniK7EgoTUQU2gowsA+vs
DJ7CciNr9y8Ibt/rzqUnr0fZpDh43iqqFpFspoKEm1gnjYt3ds6SlnaikDZUkg6MxhvWqzaB8ov9
r2dBeiXVDisIo0Dv4kidTEfu2aen++L9BXzNFHpzlLNp2h7bExGxUSQmHUQ9QXU5QmcVd/L1bZfD
2qcpcF/zPJQqrOTLXOiX2zGsMzNNZtuR4kZt0rgCJ0VSuSyWBvfSE49WnM4uKywqx7+UWzpDypXf
872jf9KvX6zmux9oMP8jUh+4hjAu6bnPFjd6zbsyjn6HLlQ5ZZmR/B6qCCibyd1+UiPLtuI6h/uD
+Wlh/ca92yCwSrxxW7Ac0BUOOv3ztro1k05yCPL4pwHgiElQaa60PbeDZPwto9a3L8dgHBPunWeu
0fbyiaYh7ewtEwduZhltpIzjuC/m82nAPpb3fhyLdndquD0MqaWTOQNgg/4NmhfOBPRyykbxRPO1
FnDtNHBggDxjmQM6+haG+BW1r6No7iH9yJSCBXbV8z+AldZF7VoXOId/YOFBXtHYS6dDOCFsVyQE
I6bC4smKfDUz88tHR4VNKU3uMWm/txLPzdTM4tUk1P1hF+7mAAifMn3qOfC6ucL6Xt+xZtb3tEe4
otxwdtV++IScGL7UKoUBMgzNIrr5rNJGoR3fl+fBvctGl8rVHoxyiflIALoljI4YMcn/+mYqN8hH
fSjoY5xOAn71eRXSEtPJEHFMKHl1k202mHs/C6+2960cw3/bmX+EZWN5fi6HuwbNrWQCtVrKiRvi
g4VcWQPmzVQPItV3e5O/C3cbyUFYf34ZpMY/FxmiJXwGvdYbXSJ3pAUWxsB27KV5qbXhccnFhEBZ
DOCjuMI1dLeRdGguvSgbbZhNhZhZlqWFQq2m7CPgHSz6e9bpaamh+LWETzhPrBWrH9w0P3C+dgOk
VJD1gQTsBLynXOUNH8PCC01zpAlgUQy1f6dEovT01bCgKKd3vl1vG4fQFcQd8hO3bAX6byKNOKA8
8mmPFo+aLFLOoG51gvtWLPQzZ0PhSEfOewVCBee45fDu2j62ThFoPrS/3G/hW/IOJ8JwymDE1ejA
IctDPAk4LpbybYjHhqKFw0CSJpeRKK96RBlroI4NFNf91Zft5uD7ovexsS/OcEQGeJwG5zySmI6p
2DJvDTcY3rn+Nm6Uqo9jOAbgq/tvfd99MCdKFqeZXrNpU5J1c0rU1xioVe/A3+qZBA6t/aF5e2La
nWE/SYqk8KpDReiVPy6aGR7+G/lMtKBsMKItDzFjh5GI8SvvNk51r6bHp3hxQJm7ZTMLjCp4AzwR
atxQtXmcCbwwHJHpu5RyJ/arTaA6ka0TozWb03ZrjZTGwPmqzoDwd9nuz9rlr6Fb23G/X7Rhn2YI
n57vlZEyAZCfv/5hwGmXyNd6ReFVJQQCDZ6SDfe5hg2fYGZ8gNumNzh1W0eSfmKWf1CAji3o+Iyr
/w+wiFkdkVJgojjYy/DFPN8EK21DCU8cuuU/WQsbgfZTuguNwtG8xMOqjSqrsaGRkJY4i8XzVINg
GwfUrEFngDrKPMdmWFrSellf0uifqZ+z3wGRceeUIa+j+KiP41iVzyqPxDcI9FiuRQ9s9RDYcysC
Qf9MI5j0P90pz3+KoBNJNfUdGjgrBWdGiVBHFMGArwU94tERE2/cTmqp/muuqscNJpsF0eqHCj9d
/WKTtmpg+aqcbL2xb6wjTmVfeVgk+OQhqh92G/grBs2h6hfmebINTxXk/0bnmRR7RBwDlQU816Un
XLgi7GQM6O0gYtEfoAswj8h2jnAumOzLUjR1iq03JeEEALXuQ4wKsIvWqcbPj5Dow9t9q+XOjppn
M13dj+8RQRqKG9o12C7hbv9g0K/FxYdl33XcTykBxrFTcNcALdSavJBgar6t/Wo0zMaDRTdG6y90
Dy+zBKT/0JFDQ+jEkkWokoTzRqkmr1k2tqmEuCTl9sBal6cxYUu3QuVytBAaoelkemUxBVRdKO5V
FDtUMPYRY/58MtghrWcUcg95+IYO9hMQjYBWtFuxVj0A9rRwYi4OyzqK5ojGrKi4CXlpSr8jAn9l
S7kl52SCEVA7ra28gMNUdUyMVK/DFIk2MQit3St3eeN5ng6mryUI6yX9ie+qb7ZIOul+/PA7Non2
Vk/Gn7nwUN5Hl/ItzoQ8nP8+spZhYLcM5aX/dRcyJzwdJvMqhih9Jurv6F6JDvNu9N+iD5gjYjhC
avbH64B99Kn+E/CuJA3tLwn7tk059q31l9CWaKznM1O9vB7T8JoyyYYqPfl8BW0BoYUuc0Zti8Sh
gnxZpz5CVTO/bPEKDir3ugTWUx4K2UHhRZ5dMpl4MfALHTgiihLwO02F/weUucdTTPsfVu1ij7a8
MPgrOHPMasKKZ7UJ3UTj+nsxP6APj0XbzQc8aBTicUqkwmICmJqbrmVbGdF0TY0Sx6dcQ9Huw7TH
zN+9/kV9Sh7LtUwsI/JeaAB/7/4MvgTmWFTAYle1sCX6n3SCiguNzyi0R9fXEjCRAz4dePB2devv
jC878D0hmuYs0PYPAme3ZbMJm0ymG9Hd0NpIFivk8//z/yK+I1xzZ9gwS5uTtSG9jE5rqOBeAe/l
ye7Ejl/dBSn160MQayUN3TmbmytRFcxfAkeUzJhzYiStOAPq5NSHvYf6+EAWCFyJO1BCHx4PfkFD
MyApC3/1w+rj2jha826bkRBnUUh/EgARqWOranStV1DvXELs8X3TmPJPGaqx1qc9Xy5uy/vLrGcx
bQFttqUTHXisx8RrRQba+aA2Eu9ahWBA7Q7HOTaR4gvQwYWMFbNZdTdd0F4ASfrQLZMK//RxLNUh
cjefuRqIJ26RZsRtEmPWvY2F13z81KNXq1lS6DAsGJVvrvbq4/ttjGBx+MZOVJ+TTV/SRj+3HjUk
KzQuTuJFWjjgf02aBfw7cAIp48CCDZZf8o53S2AHHb0Z0IPgqFeBlIQwfn0MJm9WCnLV2lwzObVh
IeI4rXaGk4b0poZ42eDxbhh65Ub3Y6F6P3sRndR5lNfa8ldy6ZQP5mh19oeWSB9Z6Qjje+LRdhib
Evb5syIDVoUXqaD9zRL6B+4+/kNSJRLI4ImGz1rLtigsFe2KdQkF7xgE4E2YuQnFrUhDc1xjG0pb
ZVFYS81X6wm3d5HZkLsbVXCQoTI7TcxK00tdJVjklqc8ETeKK/EK4fynmDwWi67gtohrCrdrMbl/
fxjW4Ayni6LKgHnPv92KbdbaWsfCs4IoVVkr8YA/9CL1r8RXC77Qu1Y69F3rFQ0A4gf6SHLQflJR
+A079XwdW+0irM00GxcqdNCBbZ42JJT6Zi4l5L7ZleLtGWU3xrkcplqFJ7MXirJH8COzujJKPN4y
QG48SwQlEAezaAyygMNCTgbA5RKe1+l5S9z2MYuBdt0IE9tVSoYnpPDzIxj+g4j4+8jp/4GB/vA6
7j4fvxc/G41zgHcdaKYa7W78pYM03juPyyaxHBReXQt2/Rx58aOLGTQmed7PU9i+MUKWt3PUFMgY
yMSyMHfZzchSTXwICZccacGitJOQaFKgaSXvmYy6K+Jd1NmKfFJR0FAMtZ8QQiaX5L4DdCLBNpz1
YKDgRKNe05tYFU4v0+N226bTWub1aiIf2jZXUpQGExj6gtKkFI5BJmwENeg35XecY3c6kdFvjc9l
LYx3okCMm9C5Se0smvYyumy9ouCioFKjVJK+SsiBShKFTgeXB5r9XfXDKHiCAWxucJ5+Q+u1CzMK
1cymJRLK91uv2W4eYXMC9GcgfdnSuR5xDRueot0R1xpgtsyHIqDAWXz3JRXgHQsL5gKeJASmBok+
CaYp5vRZKcbDqbJY/r5QjFI741kXesKx0EiQekslfvEnb48va3yV+9o2rH603KrKqgKaQFgTCBN+
XzkmpfDxYjehIHgyZOG2Kvm3wNSFjMUnBv/cmM6E93b/ZNNf0JbUCCuyZQCUyBxi/Z95yofYI+65
sIDtuPnlUuf/ohgcR6QJHtsEpkPF0HUU6YTTxbH9q3FtXyg4AE0haE4vEXW2LeFxTxZGu0ymTDa6
1o/VHoVnT/OoLwGPAP8f5uZGCAwMugheTi33ZoH0bRcTdgwACi3QaGhV7inaIqij1vARx25fcmF7
TKB+cpxt8dI2HRvgxcjfonqnlzjhUVtLDUhDMLHZ6n6VrhCJSHkaFtlzTBKOD0sBrvmFRXFPJ7+b
WI7eF574dQBVFNw7ItmmtjzZgN92beX9FYV20uIRyXFJFu25CsV/pF/5ksS6gh8acWYgGNP/G7sf
FAhCabDVo8wlu3eMH7iGMEM3h0BRX0yXAKCn7HgEukdmSUp+Zmtrtzpnva6QLQ54ktF77u1pVTKe
6RkYuL7l6s0fxvwnQeerWsdlk0cwprhXpODAyyKa3zKzzu71GbcwmmSmdt/FhFkAkaNpH452818R
eiEmhJAT/sXVUBF7sd4LVL772QeLqbvQtqwUPka7Q5P52qD5Rd4qqlHS3sFq0M+Rriv5DGViykgO
RykODd6uugVImqjPQqNlAtv6t2Y6a+wmbAnpN8k7fTCugPXx5+zxqEv8WC1DKGxY160Hk217d/pV
eb2F3DVznJgFi0McN9CZFnk2gS9vRT/tfd150Q4ljpGhx/bahFgqz1kJEOBzW0Y+NRbQMp78rLPx
MG4/NGbowNLzh6AfokweWPptQPRmoGSGjZq8k5J8O+amzRoKyEPotlAIVXRuNhcEgRCiPCIbyQMu
YUQYp0rYj1Cd6mgu2bSYmpjJWwkbWZ05rpG2kRDpl3HpgbBdmgia350rpWu7hZcvROg5xzhsCI/4
pKmoXfuRyZUklV/89GoaN+S5e51Mp0XSNO3bXdBa7g2e1Wjg9MAmDJa/BqM6pa9fSJXErWjwOjiA
1qfmZyYFfSvsTcOhIjqVy3ZbY9oCkfxO0m06iRa93+lnjN23LGhlPtTTi/lMzk6GQkujTpZt+9z1
FhsFTjNbJYq/F+6SGi3CY00prCi5rCZQs4mAahPAyj3FHHp9lbRtJKACrcxbCxWAgYydlrUDNVQC
1EAHyullIcuCk+kF7klGRsycbSU4PbV1Jiib8kyQnfODZDHNBN9uibkOVrtV0OcNl8jLdX8+Oga6
6MISJoWHGhqLVMQnmSGw8K5rvSIzrVtluINrKocKjIIxJlulB+i9P1wyFdalfcArGx60TInCcpKx
YjXv2fTjvNq2Jnl4wNb7OmpIMqjhw6KnHBwptyvtu8QErksVfz5VSx/FUURAz2uk6RFKgmsM+CFq
OhyXwtEf6rDEg7ZjWgdumcCcShNuk16fnSrJ5ONvr2tp9cSDgl5c7jhcXhM35iNtwvMHQjpJuhyT
Egl0J9l/eip6liCUndTPUNfHuOnxRQSzx2ScIrJ/4kxZBMElM1ai4pAzgpP/eK3PQvUARmk6eLD2
3EYHUdFXQku76RqUTOq3UlleDnt3NXJkodSP6UKoCHojrXuLvicvnd3Pzs25zJ5Oq091X0vtdIay
ynAKob0mIHPJqfLL+UXtmChAxmj+Q4lTpHlUyebngbYAWvhCn/KEipFurajy7E+aPKZZ4laBvKKu
rIu37svTbEAlZnlt/zk1b1gtOz17rXg+JB2GoIs3mWDPmued2HSneXpbZSBYei/c5eQsGLmkrWGb
si0h5qeVKhxqQRUafNsUlgPjCVv7f4H81zafqql81zV4lQLE8+GUm9pzpit4ERHLFSB17GYA7h5h
4W5kf8Sc4Y9y+fKCo7mG7Q35W0bdgJDiuxf33wndjDVZuNv42RGvjjmORKT9RmfHPWgWGt8ppSuG
9cQCNbE+pJxXfHRr89g5Avkg61OSYF90Seri2DRg2uEL82PMSmhYFG5d/mP4+cfayVQXuBNmG3FX
FboLt6gCJmro2AyppF3eUwitJrAipNYjx1pQ38m3pn57NMoc4WYnrf07HEQKGQlGug9oI7JPpHng
0koBS13m6OR2zpHN6fC4kN2rLPERdFECoYkbfFf7haFnoafaJVSNUiGNJxGKKq55+iggbjHeH5Ur
8ofkM95eHPoBPU8oqhyiCV5eGxqFhD1pkADw2hfkwCr1By8HPGi6Q32egYWl1+1U86Eqs8ccfCmG
peF6H7GCMTEdNY5qXrhnFUAfywOB1bHI0G+9AqreGvoswx9CpIksolwZk3m7HP0ZOEOQS+6mjH0K
6ED97OYvMuzE2udwY81Kgg062OtDU4YFyHTyTU/om5tuXbNJWIvpSmS7UeSpIvxp0ZKlU+pI6j/y
cRqo8Wpm6kutjuCdq8B5OSZ1SDDDDzAinu7YgRWL64Ps1ggW6LdZ1MrcX5qw6uH8Gw9/eZ/iQVnD
oqI7SaX7+3v8w3r+RkiCG2qbXChCvBZ2unGXw6b/qpbJxdBkLk+1A5LY16GOQgpBAi48klp35LjT
XLvc26McouICSRZZqkZMVJqTG0zCLoJvcieJgzt48C+Lmi/ZBhIyHFz4cem3OTFdi8cMIZBKKnbc
6gZeAy7U9/mRX5x2p3Nz1+69wFBm6xw7fzydFqfeaEpi3CY0dG8xLkmyo0xS+TEgpwmZTTxLA8gF
XnnoKu9T9yAifJh5sF8JPBs3RMJAZj/TP/t+u9Xmog+5l0tv0YUiziFNH42s6Ua6WZlwfFohqkYC
lca0pmk3x253hngyHMDH9/3t0aSWKX+Pa+rG9j9QDQlRYNi3qkeIW9gmgn5bNhui5CovSwBhIkkE
/z3ZvvDwlnPoIgigjpvLmKKZHNHI0ztpC34kd0gGMih1y/psImdmVddtxV4NyFxqb1V1nd7LOpDm
duGxjIIEWBiZq8ZHaDfiz8Q4n72eumjmX9sAp9RB2KpiumgYfEAi1fRx6KqAgOmogJIkcImateB3
FbWGeqZ05qYLaUO04giNpyjfxTzLNNL5qutDWuCulYWVxhHtC4NqKwmbfx/hkAoPtPnxj9KCBqpt
GFNdIFs6djP83QLz9XqPjfO+Dv8ZRtlxds3qhc+L+BggrM/BSOrmLsm8v/CtzDgZFdNgtxHEahH8
5SaplEU/CK9xdaDtlwVi+RbE5l8Fp9F2xnJJFKamJQKgqBqEdr3aHqwY5vVC39zwyuGCUEoyNBuT
ZVHVvGPLBigv4cy6ZI6J8npaoQUTjG4W4mqYCp8b5OVErS9Fg9cDkKFcfsQKUcmTxgH+eaGrXpU3
SbPg51Hu3chaCvwDw8wT3Y+tsIlUOVfT1BuNzm2lBNAgO2QPTIPPOjYJIz3PE/iEcYjBqNFgVQvC
yFa0rbNEPFXw9CTax4qkzWCDZpPPpst7W/BtQVpvTUnV77Zx0LyxgEPEqDqIsszUmOhyx6vrsGmC
waJ/RjrvbHk6SLYDKEdR0WEyGHjJnCqNXAjNt93nFcZ7CbnEd4gRUD8HQ8TA5aIHdzh4yRTQJcQa
XzpFHLEz2PXtyGY340fhsh1OaIs4oR349a9KOkAlSnFq9xYaQBD7Xja7JSMRPcF70A7L9qg8ideB
XFzNsaUldyJit1LFnwEDEY12riPdIoo4Fw6u0++g6SBGUqp6LBgEBFHck2sNMRDmdJ48KrjX9UAj
i5Z8Jnli0SEnQ70YQfVKBKcNCkV+lbshB8wOHbKLWAC/mNlMscZMDsEzAPPMWjQVdR2soMUJ93TJ
pRCHvPyxDssKfMTR/O1lp8isJpIYmD3WBKcivARYKiDASq2znIKlwrtcru5S+WJM5LvW+zSDpWux
qs7qiWg5lb0thQNEM8xIIIbdMIzDSO9+wlKvzfARiZKIDbNRrvKPimBMIJz2vohKbiCgPeLwJw1H
1ZY2ISf4iMffKYEGgvCMrSmFgyPGBQkt7mtNKQ/apZFZJ4qyhmU0hDHzYbOV6DhM4K3eKo1s0B7d
RSrGeUk1eaulhyudtq5v+9S+mMKJH/yjTOmxIgrrinjw953h/aEZtX7CXE5Uvf0woVn4H1L3Vc81
XkaOZZB+vqGU4axWrqcT9yJpHlexlJMqVTvvOJt32Nyy5uJZnbWNVcfByZM3QPxBaYh3yD+y0KP8
xe4Zm3jPt1RpdClXE6G2zlo1WWCTTHVsEnuEWPRIZ6f3/EmUi/+ZqOSbZHZLbHqC9vMNPEQ40Kmw
jrsddXSNlcwQtASISJ5OmqsWhUZjxy14YUgmHVqdxF6ZSIu+l5pJURpcmq/5sEU0Xhsz+7uEetTt
XMTaU89e2EJf9kDwqLzXQ0s7LO8p3Qlt2fW3etl8F+YLy/D+FFppZfnCtN4L5JEddv/3PsMV+Hxv
fJ7ZAnmoIOJel3JOKUOzFGrNRmPz3F7Pw5p439KpuBg2g/HCbDgCuoLV3rcT7IxfSITtVfV76luz
tAElxGJ7RTmg+j/+6vMRBUZpmkEJqkNxAguGjf6jyhEjzDjTAWWkY9rW6IiVj71C87njYqTzkdfW
6RrnfQS7tGYga5FYSdfhSuajdwyLq0M0N2VlGePRaoF6oDck7IZY+D3au+B65eTA/M4r8g6nKuVe
z5XKW3GCu0SsHt0JwWmJrfTdnrHtCFNtGySBTw1ZudKLzqSIFHBTCRWf58i8JSZYfWWP39+i0pjJ
WM08rCUnOSzKLEPRj2kP2QbgQWof+rYO+tHJdMIuLcva8u65MWwnDIVBEVk5s5eK6iyvpL42bx26
YuL7C+v8CqnDkPD9jbmC9v6KfAa61akjfp+anIKDIeE7DJ2IVQEVdWj1bZQwVRHgB+WA4mXx00Gb
lh/lqvnxw0dYx79XQeQSk1z0h3lxkDnkcHcrfyT8uRNh6MtF0xHY2fkF4Fo8jY7pNfazajlHfcBU
Nu77lo7CJpPHVF1DifGEDKQcKmMa7agPmlaLYkgCGNZePFLXJ0tCyTM8ze1Uniigf7tY+cwQoJaa
40MH4QDPMU3yaIh6WqQGMbkUX8UtxLrmxN97slF6EWynFXqQqhINwTwofBn/JKmPcsCn0iyuFZHv
NQ18YFwgjh2oMaV+VDFmZBbZ+tZm5gT81/XeUwFme2I4ztPC94ivz2h3npwpKtZ62h9ZfMioTLLN
dfNpgSsT0IYhGqU4FiJZZQFXOOU1fZbbJqq4yaFKR8m9OavX/XT3xLCJsiTFVCHDfGtWlYCIVc8q
muiO6WbhUWbWO+yOaF43tBAUTxAyGd/azA2Ky5PzBsATe8A6EuBLRKy979kW0VE0BaziN523mIa7
E2re0BJbx0/lDVwnUPXcLGL1zz5ZlAXaQZDYhzdtMsyAdSMgytPFC1zlpURwKf6OVAdWr7WGmGIK
XkNkQk+h0qq+IGT0fFT3pJP2MicdkIECFmba0KsdwytuCjUwStfDdeer7lzYqCS2PonlyOnpx42e
SmM6EMFrcZUOB9QLCg4gsa/QQaBVvMgx73zzvwedTmR/PnvCEveOghJ1CrilGZW/kQmvNOf24bjE
5Uh9/A4Am2T6nBvLEL4kdlo1wX2R6gVPrG4e/cat6G56AEWoK/LjYuZdYwGywfUJ0GB/lZWbjsBF
/L8Z2SK9wvfKMprvWPuHRoTSlvxg83KbNZp1q/ybJH/UP4tUDEJPtSxatXXtskVe/SXhOXd9JRHW
Ea7dCd/1UiwiPNJZRHVi0NnhMgo82ubcQAwqIEM1iJuylxuXsrGV8EUtggDxNjbyKWB5CZFSSkSy
AL8gW9pRJ4FmtH1saEvDEgSiDvJAEihKHVcRtgWqGtFvogAf+ePYsWMicmirfN6fmgu9VY9WR4Mv
UVVgI2ZDOxt8uGfrzanBZRtQorq7nQjt3Y7LQi3zTWHKgxU14ac53nQxk+1SMWcRbCvmLldm3Ang
OL5ScCoxhAiPHw3erNHOvazpmZ7veuaxF4ryCCSmygOs6sNfpSg+F2mugPL4dMlslWnI4D5mrEwC
fJv/7gPlJeW3rOV/TtVjuF4nCkbps7lAfg5juAgoIkY4DwHR+BgtKySDhUyQuvK65WXHFVofdyeb
y/h9N9cLpAHzddXHJXGuRquQBAj7iOh8APExQ94AgEmbsvBDvSEb1/Klz6ZF5gYFjWBv9P/feQZI
CkFUaS8drZZDpOfdvI5+VrXpDq9W6G8xQhixXS3DrQFGYzBLlyZdchHnLZbXSCTIZonIwZfw6m6i
2faIBqAdCZVMN9mlT7hRXmkGBrMTATVWcOPW5V7Ek6u98Hzx8AySdFd3Mhhi0sG3rBWN1HDYd79I
seYzSdgL/6J3XIZtH2l6dWoSH0RAXFnO9lhaqVkg5mqgEFY1Hkik6i/UKORn+EGSOc5N1mvgFRaE
TVYY+uFfk3otQ5SyYO1I5Evyd6f97FlJARG0Ags+eTb11R9tC/ESsn6feP/WibJ+pQc2pvWUt8Fg
rZlCy/WkAF02Gv5Gah23hAwYNsZpHnepYdx6Zm/GO57xEhtNw4t2cRswpMub4dUqaWCN63D4MlfI
LuKczNn8MOkTX+BHja5LbHEktLtwn2+ZhgQXmlFxP7bILJGz0wZgK+cVl/AyLnKPn4t0LsZnPYPv
b4qD4wfeawiYlfoFjjdH8AO2BNwRgTXjzIq5CIh2Xuc+ThA399+JZvv6bDOH+sKeCfQDjewb/FvS
OQ7IptNBd+NfQ8/V3vZOwbGiYtHVyYBaitbF/dTjBjJQ9QomhO6h/Mpp1M8h7pk0MoGLRF368pbx
4x0uaSE/c3jYzG/WU4hJdJ0SWAzn71y+9pZO9ZEnkP1cYV/sr4OMpwwrEtGfs6Raj2D7oxY/FY4x
vtC4eVkeXtlTow1r0kFn9MHlqII1SNaB6mpx6DrvH33npt4ZY/6L8W936VkbLRPi+uOUOh5ecLfj
FOa6Rmwokn6Hq1VaavApOB5bFkg9ebxGWOh68PFfhU6W/NTjtPT75AzDNK5Hqvsg8rySqhPmka9U
tnN35WhNs2xNh4pyaFqFxGVlPkXAaesSHTLmuUJUVbx+Z1feQ2A35IgpXLZ7dJN3yDaD70BqLw5J
wIzjg1w+YZ7fwrEa/T2DsGERPQZGbdcU6w5r7cjrIFYAaKsCFN/xLdBs1V8SFZ9ASSei5AXn7XYG
qaH1BCGHi0rWjjB2cEjblzndFgUGhyu6gNPEnPiCdShWPPNl0a1oz6tfcR9rlhWjFpzI+Qw+DZru
mEhvdnJb9E2J5nPPipM8+YK5uRSOiLHWdEEiOEPPh2OvRp8/NvTGJB5FDB/26FeMYh6jf2GPrOxg
vDtXSbMJGZk/uIWwnyZ5RDauJiRJHrykeGpPF7rnKDIdG4Azu80S4x5AEP1x+9D0gajJEfeN65nA
2KaRi2/obBCOHvbck7m3xJTW1giqQir7tyQKhKdVrgoJRc0rGXZIrEo5VwZM9u3nd6FS0/59cmXg
7SnVMyd/Ki+73z6XhaI0s8A9FGPymb7pgFUt6D4h4XkpfhcYc9vEG22lFfoqq5AVqcme1WQ9NpG0
BzcNw01enfWGYM7RIg0fmoQwq3dRQZNiHdj844rfKqPVp/xfEw2oqY2LcX1SMY8OPh8DwUQejqYH
yJhRqpdddy8tYn0R0QcGsqd7x+nXJPlupBgsunnbeMjhjibGe68H3uMdOzPLXsTQZ0o/73BHoGcq
8LKvLLOWR4OtBVBd3D0LFeJYG9y9xYR85ero2wuaQcIma0kJgY+9wOg/3v2UQnfHEytj9rFvwdIV
vYJSjl0bz66gAqbQXbaldUJ0fcFL1dslr+lwK1pxuZQCivBmFNj+PyPLTXKVrBmawthcbStHBbEm
cf2vtfyLPadMWdguSe/cPBjCc/KlMG6IublkT1kln4rxDVOtRm6G+hDLvYJd1Ztnu06tRdPQWbFT
ZtdakXX5N0plozQu34xK1Gj9bB0OpKY9Dhwq2hSmL8m2FjbsLz9X9D4kZvL30hNWlOkLE7umwlux
BPpmSomov5K0MAhU9HpMutdyI9o9XEFxHFAzSmr2+VavggsokxwUxyCMMafL2Uk55QGtImHcljKy
czAGmoio1F6O+YIpdjIQbnAijBeefqX07zpqGrdc9Av1WmOThf4nrgz8X1k2oLJyydulW+wcGEKY
tJtaXKWE5gnLlJ4YfAdrmSwKPMlmByMqqH6i1QzaYEWPsuq4XCOnYN3MjEyOjTN7I6iIbJJCiQ2n
W/k86a6eAv9gTbKxKnSUqsVJ4MH3q96VsFpXa96NUYfEQcEcHB1LRuMHXtzcq3DkoQRHoQIiX5sV
7ymIo2ugcdY/muRXBsI1StABOg9vtiv4GdCFTiMXaWSuGsRxnaoIyDeRWwYahV+5Xno7uW7N7Ewf
ngYm/sFwCuj5DaD+b0jNPDenlk0B+IRFpItrXaweyfKNw/9LBzlryFLRGT7lsoHgcnpmir2Jl4JM
dEsUFrS4OCPsR/K0RMuBp82aFHjH44+jgnLb1vRV8rhZw25sthypSnsZnjmX9b1X6yjNSSEBD9UP
RYrREVGW6i64PBggkEtIgkpLxrOYqWZXqG2C1HBQsB2meOYf1fEJeew1DnNYB6BtDE1HgxwKE6ya
UUheHXD2q+X2QX00OeNvJcVM/HRLpKbGbnh+LO/dIFNSle/EZDSVjl2Z+wY+U8L/Ct0N1oY4qDer
70AxnkNmOr7WBTFFgFRa4NDUYDKTY01mxcxRhcTmOtNQaKHKwyAyq9vlmlX62dzt9p5+e2e/TIom
DA+BcOQtD39Njren+d54yAJ4ZCcOzJEdSrkTEt8ecxkzRzjbTvL3pX94Y8VUf6kwH9W5nA7NaSRm
1DYXiGMFgHnoFJdZrZXCT1w1EoA+mGii16Y6PhntRg8k+ieVa8KUpUHTkPQQHKXHZ8pGv11AIzww
bjc0guvxxbdhOTUGF6kw9YChyNMiVI2E4K/ccDEYw1GcWHOjwrEL3PatrAXTn65dKo9htxshjqwI
e2DRiCvQil9iHPZv0Yl4bkKuaL4KitudHnSY6M5DezvM8vA8BvfhSaRe9YIBRNZH0Dg/O+fvIzrr
yDI2PiGieX7+X7l5sQCdEsBROeBrddgS6AWQBKCO+nyMJq6365c3L9moUEsfcMpupa77xPlxL74C
jInGA6Vih0rp+H7YbSymLSCur3Qrb/Fv9sio6iuVreJqMSBxdaev8Afpk1Nwg458ce6+WntsOT9i
k3wZwOcckC9Qi9m9gpPOBMZ2yyaGiRYY5Mt+aNToC2JsgrZ9tQUSkdJ7Nv/yBwfAGhNyJOufNULL
Tgq6zuGL7JQbjZ9vTWYJBw1DjVfheOoxZWk5V5Xp7P0gKsCu5IxyxqAWUhJXP+UnPIo+2qwv+cMT
mPGr6a6Zy2DtFKz7d/RrUEVdWd5FXdf6CTb69ufrQ8hLvyFvbWtlw1YJEd8PLzLfktmogZ44xQDY
MVZolVsyMV3BCK2H7qKcZbvKyZGRG1SSClCBXcdwLvLCgfTHCcic608c0MJNMaqo3kRlfR06Yk6y
W2pOBZPIMknDh/+jtLddb1oRFuIq7+QoHuvdof05Lf7tGotPJ1DC6ZYoef4PEeUrzD6Uy/vooD8E
xNWmezr5wscK3X8MPTHoXTZghRKqTagKCNdL0+B13iLFW7tMWskjGVxilQIzpw/J4JDoEMBE55tj
KD3Wt6kvlLcQGnI7WG4ShmUsxLbg2hdrGTIr0i3GjVaLWhkbeHrL0gqEFxiCxcliUPbV/nh7TfGf
VY6I2tHjO+ZtPFciHdjWkC5nE2hEZS1uTi1NRWqn7ueTJa8OX0/aoLIDLWmU8SU32do64C82j9Ja
2hr0n/Lx0L3584inL/KlksIPosYiIjvm4LeP9OfqmFFXuaD3tVKf6xU4AoofG+xi5N6JM3O85BQo
EqirWj6NsiJYvxTKOe/u2smhCT5YrH/4moX9jjNwAm4NCDmkp2/RA+wv/ljhO+OHLFocVsVINzfA
D2kX1Oc9lT1dJRDN5s2c73kG4FoLO0G5Vug9Y+8V5hQ6VvXBArv9RB+euTrVmiP0Mn+QlLZH4s7I
UKPB6sPE1mG34zkXZA0F8pgMEvOKE16va7hd7Avixdpnsew853vWSeEaXFkyWx2EA7h4ok4OOUC9
14+UvfIp/UG5eeq2Zg5HA+ce4NBjXs9M0c7sQ/MpfFQMpcLSlJOrbEaJjND7l+W9Q10o16u0yOmp
sIjqeR7On8yskgMXFg8AQRoLgSKOr6B21W5t0hCdhemY//0XJAO92ptvbURf7dweKi02pgiTABnj
ylgTeB3gtblUKP5hBclxyfeuyel5SatXoAliT8NVg+xpejuQEGucXC6y4/gLwaPyO8ZgRuZ/G9ZV
RXoXPZKYYeJtwY5WwBXUNbndFfVVk9v4z9rI4H9qo/tYx8PW99hS0gmFr8MQoXAEL/TA8tkpKPMj
2EjhB1ZPZXdyGG2lXM4dJbuWvAha0Z5WQRyjKk1p02IxY0bHzE52mnEPLbWN94VjpnineO9g913M
2hdk80NNLJkDHm+KjrVu5vVbalizbMn2PwJYpKXD9SxB/vNDqyyv729jmV2Joqs/50qBA7ks9856
YcqfMD4DvaYJPL1IGVb2HZ6Saw8mIC90tVu/vf9tiujU16rKpk9hcI84YxoBvjcw8GAzFN5EuOAM
qsfobXvMnQ6FlX7YHozcyd8yV+o6pUmT300Wa3JJx+pXfGlmIQFX7NOlfIqyblEY0nj4YoT7LMJj
icm6I6xaMsqGB8ZMwg/SonYRRvWryDIXo/MsB0tL/jOOmzTE+hyjMv3dmt6kFu6FcTyT2Oh81+pW
/Rak3c/pZf/KOGq8aqqtZMENOKajxjDU1nZ4Y3bvJm4laVGGeRUHJmU8EpeKHdxg1+NoK0QL1c5m
mbxQml2WBmhkKcywyHh7buffqGBLI8yAqDqEkVFOqmypF/57jYliBapdxqTrGOlghpdvuRGQoBKG
IytJrdoNuuH17DVEFOxwN1RqqZ1qsuwsGOc8CIWZUGdIBu3xvydGRhxAieu5AcZVd3l00JjB9bta
E6OL90a2TlvoeSyVpXQv48okfh0CB2nVCy5V5FNcoOCWPL0HDk1TPQsO4BohArlxp+WaCSLnbq/W
IgpuJz9k///Mr/IHnJaBXeSU8BlgqpH2okS1Ptt/cNBYutQhMv6b6wDfjTYWDnFPR5xwGB/+N5Hl
9EVSNIRQeZ10VitgKt1+gBbn7Yst9kGnkBv/HsBOLalAnFs2oeNCXtelTa/1ccKCb5pIpIVw2GiV
FlzSnuhTDELRouSJrxIgHWvp7aumGJIxMPps9lQlnscNBSxXR2Pr0VwcIUU/XzahzvDfRv0RojOg
s1eQ2dztX5ushI/bcE5VBxHzgqA1qbIbrekgSCZ4UumSVurLyFyoIKtO4P5qET3Q4OjycbSDX+Xq
3sprBH7axaqRvkZxxfs6zUXtbHJ4+Bhe/DPRIgq43ctrWdEFqoAOvRZO/Uz3etLsNOU3q8xZNVuh
hKCuJRj35Wprd8TrxOVqO8fYwzGxzAVL5KvE9/LTG7XMWGzD/A+lYd+qO/dCRL3QPze4ae7Jl+Vj
wvpo1VtOC2U/wyAFRBI7bv8OkzEpzdmwdxWoZYhzUMYbAM49y6fzfn15Vux24HfSzrfwFykhZM7a
fuKMHaY/D4rhARmvqvPVTav+HJo2UH0Qt9FT9fKEqwHOA/7ZsgXaEbzlYlWWgJKA/vAN0kyJeEBw
735fk7keeM9bqPN/o/d/+TK7GuVm/IPJMgs+lt9ewwGBCN5mvA/Ds45K8aJLwqKzuGboGRPb7xVL
a3TBLBAzDESIZGgsuiRkS5myWrcwmxWP5Jb9bQfUGHi2bbga8gLkFOc3RqbQcwlR/YqCCUqhWYFy
tOHBEkjHeMLJ7J/dbOLzy2RHLopB5bV8sq0Qhz2FdAwO2x/84CRDQGa3eVI41UJQideSyqqKHWrs
lJgrGKvQkg5akHKbHsUrZdZtTOnd3rVkyrJpSrCse97yc9n8BM0zQuhZnKA6fPB0Srl/nRq1kHYt
P+LaisF5WMeoCZzTsd5vQoJfnqVQ4KAq5f8glUkwfsEGTBhCu171MLbkS0PqHD1XTx5YblEs3pPL
NKw7OBnqcY9TByjUHsQ8lg8TLJQ8LtXp8u6t08CF6wkoFsr0FhtfjTMx/S5uTFMA6a6Gx8ElORZ0
ohPz+ygg0iwWYPd8cjff/9Z5Yys0kLNsjtSGOaHlOEtqYekp7Xt3X1/kBP1BZuA4iwEjios7Jlx0
cnstSfLxLJAROXulzCCtoU0UmLTlN+s2Ac7165vxAFOmnyZ86tuorIRu/SKWOYfFbzSUqIQAw4NX
0GJNMWvKo8WDEBRzGsuiY8DIoARhjeGMRvXiwu+0OsVVSsOAv07dHRfM2i5QXaT0A4MmHMS2qejc
zl+0YkSIX0gFU6Q7XBmwXVAluojHVS8gG8Hn9PveM1DM0caUh5TuSMcp/YwEzJt2u4k+wLny4oo3
fHmVSQjarqc7fa4/3aDBI3KqRWmCaT3NuIREqR8jgagpbeO5teQL0z/FnYv14juAFXsH6GKcZii7
uUmXn+MGABxo/xZwJcTEIv7ZW9I0+iWbPIdta/s/L2Fkd/QCXWr+u//4YepTcXceVKoMg4W7GdnN
tW9ejbipDfOQ6rvQ7N+MSknLXVNgBJxn2vNUXI0XzzpSvyl+AXQrdu61Fo9UnVIP/rXE39Ub/aEe
HpFLjfrq0sHjcatInOeUAcKEAGa3yruGDu3kIBkxigsIR4lmyQqRFZp7WYesCdVBvX8LhtCwSgEN
vkRBF+SJVwSRYwuYlLen2d5vRe+LKdYOWH9V1q868q3OiJKjRwQ8oOETwfDMG+uszG4AnOGqowA9
kxW30M8rl8GSf0XPLSshTb1QCX+mzvYjRgmpT6rEkpxko47UtFBZlvlpizihV0rQE2XVqz0aNAjU
84sVyo6CFaPIpUSXVBYzqdF7ox2B48Xz+n+DbJN4WccrM/bCE1v9MauhUgcdMhW9pyrln3gHKRW1
A0oMVz5uH3TimdK2rJaBfTaiquxJNowzdy5x5+pJBcSM/hZ+yxI3qqgbS3lvTxXjzzkiTk1ul7Ii
ptGtaTmuT9LfeFo/NhqHzGM8iz9+8frwbz4vnBDBFh3gThg4nbkbYrlaug8ww8Wfimv6cdSu4cpj
fXF2Mmp3gBkFsdTU+i71+atPD6mOj1i+7WWXb0fGHopnXjUT5/UfI8Nx6YFfyaEEpsAhTeNeN5od
UlFNNCMFLKbmxbLGL/N5zDg9q2zp96Y4VFN3esITUayATiLymPBx+Zk7nLde087N0HWADAxxu4C6
cLE8wRyD7be4XLOwxK54sLw5yiyh3obpOiNm6WZ+Nn1F6zwvlY6k6YyAk12oxjM6/iI6J1Kf/5i6
AEV5eif+j5lLONM+xmvjAsDNWivZtc4WVQ60zqRb+T6qYIPX1wJaIpKQmSiUV56DhTfKG1rbcjPX
1BZ6L2jTPhiVOLmRc4FGrlVxot1/JVPw/4K1vKxHvzJNxwdPZw6XjAwLL8caU4kaTrS4SYI22Q7u
/HP2JnNsYhX2CWe1KpwIQ86Vb1DTmwzAtC4X8X3kE8vfMCuKHpk315Ov19eIrELsWndn3c/gKYbz
CiPiI+3vrnGeg/tt7V4Lo0VmXhLzhimZ9b98cLnNI78BmJ3gWroKLDlTorM/93x3hN47PmYZ81DN
QbAPjBTaaKT2yF9K9HWcYD8H6SVWfYX7ewfW9iHWPkWB5ETupotoAsrWheF9ILbG86OHWSzkUg96
W+Vh9sUm0AAyChDvQryg5kKnmR6H7wn5LAkLVhKj3XAZEQzsP0S+ZrekPMfdUMaSy5BlulP565Q4
P0ajDzbGXBpEEY7vCiWnVFDT8AhkXQ7/snxOIGbOs+NF7gUOEpzhN064iSwqdTT+n/rp1jYdVbM7
3QcmQ4VkoCkx4S+UPeoGAm6ysVILNuzEEQYrv5B6zPk/wzX58Jv6x3yeNdfbF31jZ61Jej+AKU93
y/YSyZmAg/OsynKdMYpVUox6Tm48A82X6ieMtg/saPAg2ZSIaYxKWF0VnC8grKGi2HFNHrY6CbGV
88AIUbsILyyS7czUH2Vv3wRbUG9GO2kGQ1Yxnnn1ABvnZHB50ApQwDXozLgzD0GzA3NoDmx19eRK
5ZVPsabH1BxRhJsUXmHk+HiTo9e4GhmcmncstObIlzqKgC7UQMmYJjYeoZ/cEr7sTXS4Lj+afDh4
YNeokJRQxhLExgkzXocADn4HWlonZ3t9eknXc/XYA1qIVYCPy962y+fs0z9RDw5MfvkmgByS5j0d
nO5+gF8c0cStwNMARVgnmiBj3J1NxSMrBxMuL8mSgNi1ZEBdbmOiqgzckYjbZN8BPQgNQb/zCMqU
nxs7pipjUvB7kn657DqOGhzotpstvuCNuwEGI9XoqCUe8e6vU0Yffpm4DJArtdogpHA4f7qZrOPY
UYdUEcCLiuL+nZFMmtZ2A4zeMOnQi4UTWLKCFENAmO8g5jxixyND11q7Mesu1cv2LQKcFmOKMyya
zVZ5WTNR0YJ7E6yyKGozUH4iLxcd+OHl4BIOayviZ5xQbaAUy4+zuLHwS3N6DaswPO1SgqV/Owxd
XqdBzVcjdntGGGCX/VKGE+zwJ+d+R3nY1oXGErwnBrJu+rud/RLY4uSrCYxijfp60Ei+xicWB1aq
RPtDOPQXz+RyugrrH+BdfKcwy836Y/Pa68IJtZ+ZrK8EASclTC6+rZ22YwQkhqZo/asK74dq4vfu
+K+qehv7ck+0rjejyqCZm+OTp+O3TTOkuzGpuqqqiVrozjP34jL5JKS/7J8Qxh6p7K5XUoMqUuiO
JBdANalgJDrt+lbCIbeGbpqOfn9QdPohfjgFwAxe8mK3uSsSwj/zk8SR5fsHv+wgjCBLrEl6ltGs
LofNr3haEITca1INKc9Xkvx21W58izJHczaVhfj7QJ0cbEpNZX293lHlHyfv2FAooXEaYM0s/k36
e+q6o+i5pIsDWNMXKjdtWe37490lzk8H8Os7sMuyhzSDOTIT2bUi7WYp5lAhp2Eni7W+lxN2g6Lp
DK0py5nzxgz0zzIvq5IbfoS+ugy1VHsJ50UMetaNnR2pFL2KnHn5SyAsTUdRG4UtqNiHYR0yscDT
vvEP8s74uqETjXTzFrBgfLMw6ez/mmU43JRSJhuLTIaUl94U093RWCMv7tqjpUKBt0xyXI5DJeH3
xbBipgXC9w/5x593FJY/DXlntfu41c9f1zrIeaGT6zAtmbmN7pERvK/FOr95EufxWpk9PZezHDpb
OGvatB9WsIxbQB9IQTKLs5jpYX2otXO8L4Fw6JIEmsAut83TXX03q0+EVLn+YFLdiaKN315D9f6M
8dobE5dbXCMOpqS0J2RnPbxvir8XbSAhypplGL0zhEfsQFmKeW89XypG8sij9zMjco9NBWLO0A/y
Rtf732F8klWe1nJ4bhLPhRFfPymwA26lQKLWoICQ0qrp/KgW4a20qvSdrsweSyZ9t2PgtGogCj/U
7WcrS2Sg52tVmpeRbFYJId/4ZCPVRFa4wb/cOM8YQNH963OFTnx46iz2bMXLhvqaj1mxuxtqrDzv
4bjfsabSCYNfdn4/8UM3hcyyJKh47UTkW2qpgcvQZ1MSgPhOAQWGO74TUJZkb1LNTnuA8kOVICGQ
Re90D+LjCKrxqHmyzdcnsesNhn1Ca7a/RszVhGe3qtT1TxGLfgGTRTSvv8IE+j7SFX6C1T76mpmU
kYQOAMk2J2Bzn3ZjV8LsbvTyu6v7xHSMMfFVOvdEBnHjX1RfXnqo0Q6iD4EEgi6iTPsox/e3+iPO
eCq6TyR8zjyFm+5izKpw5EsQZQWlkY+DGp5g078lJ/zCloAB17xB7kQgbgRVjRxImEQX3WMFuW4I
Kc8r7wChgW7vokQ+hUoBIJMu47McbgGRChn+niFDdWDaXC8Byqwe9QNm8F3nltEI9HTFj3S7m2bf
grBd8fdNJT0BpJV8Fnp+hwp/aVoj0ZiUCbq1ZTodG+TndrdPaAjlyVgyWikmPc0o3rLEflkV2DN9
nn61WEzn7YsRuJjBss5m7yacEDYiR4NAC+T3iXerswlozEjNrowMyRQx38B5/DN3hnoVCtbS7PTZ
N9jaturTZRqvRuBRUg7r4AzxStvroOps4EUD3xtbWoHmFfQ1+IhCrqfsx/asc/4vwaxwYLFj0RTQ
Z7xQilTQUcg24po88rNxVaCAYA2t26xEvuUaDjfAzwBAKoWQVczZCpe29q9VL1rVdzoJhaK8W/P+
75oCK4cV5oUnDs73jFscJ44qwuCyqDFEhHtEnYcHs9M0DZQEryxqauzJDah9E7QLKo4O+k22Oy6M
r9pAmFQEg3rpLqoAbTcuiaT/bYbJKgk0KVubu4acdPsFFqdEZAuS1xN9cBZvmXxwJul21Jo8S2oh
yEv/mGiK61UWS6ARLSLtJXdexfljA4qxCTnhSUNr6NUoYmRipQtQtiSGpnaAiamgPtHUqkppnOAx
0luK7vDlpjldrAAaNd62xCJCeNy+EQ/myEfrdpUmGsMNiUAbQiThOy8Lhw6YrgBVq13Em7Xro3ZL
PpcJueyk+AhN2sCl8f9+kqGqhq226WyS9e3OII5PS4YW36hNHPH9IFUmMb/JBOoplOLWYPkJhNCI
KNgNlSgEhy7+Gdf6HWqNsAHZR2ba2sJ/AKx1dUqrfZy74CqS9AXX+3JDeUFgoIbe5W3EAFK+fZ56
hzlkzCInMqg3QqZ62Fu+E88lzC/Px8gZImt7AsclZT87eDT6Jsmi+KXymd4xU9r/YBCA/bW/JLOZ
K0jH0CtRoIOBHr3QGDycGtYIWCpvj82+PgWAr+t0aNX5OnGa4MVM9HukWlSB/OlJf5FJOPQIALMR
I0+sUYBQjPWbviFVelydppjdUBj3fTpXGIhJzKmHPhXYSVTpqYqTKxsFHdWIZme/cRS+k/HGLSTR
Mc6YdLgxkiFC8H7jjTKbyOTE5l+ZFFHIgVACA1YkC4Ogv8eyCxffZEQo9vcz8/jp1qsTSkpcE0u/
m2+ir3e+4nxd5hwn0LUxHF/ObXdkYFmjOMCfBqGROgTQfAjx9NDxfC1GX6+Wz726+oKqPKE3K08s
IRma4sHcfMPXo4W+049XVO138tD6KkMHmAN+xbVIYxg+YIQTbFAwnzYmOOzt/WW6MpwuLuazle2y
xa/EBgrmF+QZK8ZDT3dEh2txn441BVFgeu5shw3DWqwyxLjkY6oaJKEhJk3Ign4Wm9lWjWmRDrq6
CwGfz9OrCWZFiRHLLSLT4LE6GNhFKgVKpw2NvOuCLk8WMpN1QMiqhrqeK+VSjuci5xnuzcPbnUIx
ChUch7Pp4DM4HBpQ8R6gaj/OwsrxBEy2ryCnvzcD8zm1dSGfE5SF+JC10X4YVOwT+hmeq1RZWTRX
Tx48nP3S5Mcp0rK7WBfK2BtZwCjNrsH59gvr2OPh4AxrpYUhGyiiUS2KhVcVqhx6mAKxIEisacOe
zJxL7EwbP3HqB7T7qKWkdjzVwJgY8TQNn3UpUzlVKT3j1QbYnZrnzPlRbwr2TcESR8KwqH9hle6/
y9enEGRLg+OOm2X9XA6N2I5UvRGHWp5ba7giHo3jMltdSNqSjwTETlkTrDY4DN2qpbMIef8x1rH/
eWtbaMkXzNJ6dFJPMw7Kc+zNl/C6jrdIvpNu5xvylBIpQiO7UKwjfG+pDc3yVISqMCbVaXop8y0l
233pK/aq448ogTbTsoVeBXCk4AYtYv99YUE/jmtotmlm/veZ52Rdf0TMFLOnVBguSCvqfDqMgpW3
Ym5pDQhumGIlLdg4KPPCMIrPr+xGFlI2PmAo2Zf/zJNLRAKtnHAzUGjJi+cWegc3khgd86ps71OT
Tf3sKhfOecePX6fxuSW8AlnpSUSoJERIEgSsZSW7p98MZ/B3pSAvqr4Uf/GUPWoTvsRsABJjDbJh
81DJaWaXELM6Bspr3sCpet5IaT9ZumXyLSWplc0wGw5wAl2CAmLpvWPp5Omuym6IDL61oeulMtlt
8yg2wjy/eyvwo0C6AmBPm1k7djxAZ3ozMs36dytWRESFerWI7zgMpLqSbDWHpZJpd/M88E48RmdX
oYzOqkxlcBd4tcXWVDfleAj6d/qg2Hq8v31lFMyPUQ2anlKvVIybDQdPOG8KEvuYIU89Tl7+4yYi
U2hqdOktrEE04wXaznRb2gv4RwLH1a7quiUeVgu5SeCLbpqp+4nc7u573xxMRywMqZYKoOi2kz8D
pYxJd+R7R+FNBR3kZpIGgRdnqYTUQnpBw/JP5n2JXinf/J/bpmZwhgFJSz9rku4OUEU4osNSbfzh
sCBTMr660hBYxBenyYb5Y2FY33UkY1EzXgrqorY5nonyWRiwYy9A8BMB7O+a/6mBaGV9Kha39QVK
09x5ZIQCoWgLj1jgzfo6FOw7hvxzYPpKuReY10wpbyHwkdxWWDK8Hmcde0OXxx6aScuYqvHa4N/J
+G+z4IddkLVjAGHN2t+cjjEyPQpNpijRVR8Rnk6CbDH5GXuuSGgZXzEmKu/JoxYBxJ+Srqmq1f2D
ZW/VhFULV8zWxtxJM0/QCJUf+LXO4AgdQDD+8IOgPVn4NA17eZHgA9A4o+BmH+6UIahkHelazKth
JJiDv093x9GQzbZ+8zgmT0mb0s0YSE4RRDvCfP9eVSLk459SnEiqG3ZuseUJ/OHOFe2YEs8Y+60q
SgM33s1Q9Kvdr/X+wxU2ZxO06IfTSJImS7R1Yj/dY5YPKiIrZtF6UEgC0WFJ4vXZr0WtISUmh3r3
qdtwIX/k89K5IzWwZMHE7zUcj8/G5vgF+TQMD2DkUR1seUqKM3W5FgU43FUHIEknEXdr0HAmev+1
WMswQzj/c8oU9mlgXJrsi2y1AK5D09zLA5G3C24U4S3MYluDrGp2REonsA/e1F1vDlM6KKlbkL2t
yw/9VpGxyFGV0J81ynyrNMefuTDhDDDBqpcllQWg0H8g1wxeoafsNzqC3qEWUcbpo+X9rUtGCQ8y
SPwKkr/6BvoF4Njru3E/rAjtunAL/z1wrceupYTHnvKP6yKd653ebJfbuaT/cgd92jxpgklVw11x
96nVf12+QF2k8sR2nAmbqf3nuAjIAJ9R305ElGOpgNzZ1tQ8sMQDegopZxJCKil0QeCoFOICVKIY
oGfxH7Yh0LJ0wbzpSTZWxmXzqfNtThzl2Ra0DU6fpNb2aiW0IqCt+IYkyDuF2Sb6wOu5ht1qmZtG
mNhVLA0hD61AdPyMU4UxP1aTHubI5CBzLMyywAJkjD9lsu07Gwa/VPZdUSRrp8HxujOQ2J8qIzUr
GTttzR5qnUy0nNTJxYRoyIyFZfAxPIUtgdVXYwhze7vXH8VLZeQ/Gvvj2t5T85f3crDxzOSbjDuw
jplPQOFu6RcYeyNev7G3j6s2XrXl8GIDhBUSqduWuoowSOz4Ybd0ktMkikIBtpQ6qkdD+KQYU7QJ
VJyuKdtCVDhp4/7L1mpAFP7dZWO4ryuTcuTbXG+7U//pje+JbZYf07kwacLikdwhXIsl2D7O8P3L
fvI9Oqz2VFyzDpmzTwvh7YWWbFy4YsIXWlo9eLnS+Sk6OkOQ8gEfWhvfHaRB5hfItdPZ8zv+w8EL
QCsTasOu07Pytpp7ytDRfem47nWpCGa7bMrrNCC3FDtWydX+wkymmB5rGxuMauiiDdzC2r+ENaJ8
cb+r3NRs4RRaDS6Dj+6rnP8caia2lLKquZ/5uJGeMGLwivcizbiVGmhUIYyTLdeuVxSgbMmByL3X
XIIpFQsm9D7QiYOEAFhpdLOp8bYa3h9s/mx5zrSNvQzExySd6ljlNip4fwWRO1MQ3hjvSIUMY04G
shbDsDF8FmIE+u4H3VKEoVV6ihlCjw8BLW1W8d4W+7DjKWch5fx3+eHKPFP5+q1Wh7nILa/F/ReM
1lUmshqATu0wpX4VbyL75iOSmFN7hFy7M+Q11WFzXtkY/4CCoOAZadglkyA3O+NyQcXDnZKhEUIZ
QhgKTxJYd0n1iAVLCw+AhZ0PGnC5WQwGSjpvZAg/ajfrNWR97n5Taz1KZBPxHCQmVTRb5FuunxW2
F5oUQYzU4t8v3F77BJ0y75ExFFtQ8LsvwF7oaHim5fgv008VHND/Xefju+D6CM2Pjs524lx+9h74
XLCQcLM8+N/iAjRnk4rVInBY5UTYVWsll5ReUXugACU6MbP4QmkLgGB6NoslqNNqNcU6gr0cwtmL
3dhXMA6333EVTZXTdLaor18rSqS0X2vHnjefm+LIXixWRpAdHBxRg+tahIkv+X49NHOnGUM9xQZD
/N9ud6A9vcroi0A9DjRppNWak2eyFPahKWgTCuGCJvHWn4+IXrMPH08T1HAGBcT5HH8M8pdFIe3B
8/IpiSkbrW8rkPBUZpT3NWut3lUUHEdUmn7ADXG6zdNijLBQ2BpGJAyT3VIm+GsvcGseF3kyCP7V
/VzlIQfCVseK7Bp9moCBil+DHVq/St8tmNr/YlHF7zKIWG37fMJU+ZZVsUlYX9bh1VYX6F7FtTCS
jO+kvlyz3g9H9V1LofBAb7Tw7ICiZHaanNpmtoV3TQex1OJdvWDVTMa2ctDJ2wbIcLZG3CvlKteg
hW5x/57DYHGbOcmp5Inf7YrwocBp3zVlUEiAKx/pKo8gCcrow3B9eCG3r/eZBgEI/vnhbBvACGBD
11tHAeD6DKysXvp5rWJ8rncIfh89WwB+r8qqUkInjnF/dWZkByQ89wdOkVNIzMcOr6DcOxK6OXqG
ZvdS0O4O8zq2Q0T8+xYrYV4FtxdMdwMVrmzbuNu+PGND98zWQIfAErf4mjssnIntwEOZVq79hY8V
K8Rf4aXXhMIVIDkbkUhlYHmY1dL6nhfAJm3ZNBL0GGpl9pK4w3I8X589NdVj3AnWqyciCw/8I8f9
svwLVoX1n1RZj8kE+zdl45top0MtBtcoLf6vsiZg2/41OspupDtuxWWHcGljikv5AbirQjkguRE/
Gvw0xmRZ8KsyTFAJx5xN+GAYeoi3soNdK7G0WymcQp+n/pnCXUQGPBxbzSv9kOdXgegkTcBteKQu
zikQk7ujpmgSMbfSH1l9ZJW+hK1p29PuyxFQ978Md2LzU3Wz02MFdGAag0MoisfWiu/TG0aLN5Uk
gQrDptBPFwDBP6YtzmDX4vr/E+KMY/1R3xCtDd61BBhaqKOs4LkNmaEA5AytfGc+D9MuUTt/exOa
Tkiqn2wFLcNY2/t9aYmSbGM0UXwpTpBLCJIGaTY4HFakrnun9yV6Et0271RN0MJ/Nn7nFaWmijnW
B3w6yjP6Y3J1/UQ0+PkuY870xs43jZpQXZGpjji/LVgQgH8yYnek+hko/cQQKzQKmXritF3vu2f4
FIgyn2slpKLn5bDZdhNoLo+0Qfc2XzT/g37nw9tATce50kyuNNxSMiJQA8VvE2zgAimYgwZxmweV
mUx3ouukT0P/DrjA3c9VXfaW2QOqQBv1ptagSUAuXQzLPjniq9637KdTtkHl/jkXRa2kDXHNeF7k
1GZvs8L/TcXIeQvtYgjYThl7+uDzpVP916YmPYtLlwv5w8Tu2rKxzHLkkjF0G52rbJuM4oy0c/JC
Lx8bw6wOdH8IDUOjcxKRHNBB/0CL27vppuF3M8R+o8mdBeuoehhJqymoZy0xGHUQ2K4id0Fx2NHc
jOH6bNEYQo1cVkbLEJ1niNj/IvyO8SHuOOofncqbvsd25cf5fXQDQN+uLVp1tIzcveHfUUWxASM/
Wi5Sg/KCmBLIFsu9W6l1Z9ZzIXcvrSQK8bcG2/RHimmaKHC75y3w3Yh3x6b0Cut61Aa0QzMfx3Ny
Ko4OZkFWbi4Bos+JXrem5uc8uoOJThLnmOeYaytHREvVwFofDDt17Fez/uPXOI26r5CyNfuXbO5I
z8T4QS4sfKmIqBWMDxzJLuIE/BknlfaKZFH/DlW4/BDdwC0UiZxwG/GiTOZD5VCfAx209/K5y+38
g2ma3NeORjaSjOdwivYVndIRBd19xURKGPEOHhoQ2XOTu6poRNB9gDXDYm+z5ZbuOFbe6SkAPPV7
mHYsZ04SI08TfXYiCwzVY64aIurQkFw7qRujF7Ng0p0rOBHGkqLyyZuSkbL1Prgvy+f9xzJ+GV30
Z+RRqU6yZDtls731wupk9aYoCV/sqxjKpEYhMMRwPgJGLYaGvOT+ZCSN3oyADJ4nxPoWJxOaYPPE
BMD4/f1BU8Dfhaep/jcHVKIw3G0/O39Ila1ON/l54PKEUAfZXcOH8+hqq6zcnA1rh2v6t6Jl/d8I
iyxSbndDVEDelueCAMcofk8ltY+jVb+SioL0Y0jHBQFiKgSiJSSWraHLevwUm3cmjahHlsg2W005
d/A3shHMkeSLqgpLcYCPlYjQtlnCRAKukmn4O1BO+ybqmNWowgRVgPOksFISIARJPSxqJPyWOTxe
68VablzNuQ4/4hQZfB8KPIOCHo7FtGdTxbLN/m6PY6PT5N11zwnkoGJGJ+j83xWX9iSEkfxEgujg
D8euU2ClQwnVP7SdY5IXWQSGOQ7NDtkFM5H+6uf0HLaI58orprmiwhKoZTbloC55XWYNMUxpCGxO
5YOYqZUkuOtyeqygdu0o+fl0beqsfmc9AiPy3K3z/c8IXf2drQ7LX+CILnoF1cIqEZsV+w4/ZQ7j
thZuK8DpQQf2ZMDEV67F9Mc3L9hI+kROZxeFFO85l5bkEzuPie4+LZE4Y2Y5T2O3w0nj3LRcVNBm
wN1Gu4VpP2dqPiPJyEJZ8beWzac4kI1BBBFYC+hNq8kaUb5CJ5XMlLPeext6d5WU09lLIth4rwsb
8sIKCGi1/FZ4bzwkiQQiMDSewlxmKIUY0HK+gjADCI/Y8+Vadvpo03RyBXK+4EFbmDvoUkzK0+tX
O+gEi7UrQaYyF2Lr3UdSNHz2t7XJPe0eDkAB1HcfHX880yjL595J+IZHsiZEJLak4icPzz1oa0Ej
s5SCDgfh2MwK/Iohx9NaoMVU1T1E+sjUzsjeQhoHd+UzQ4k6sxb9UqJQKhqlU86ljLTz4MlH+bJa
3TjEjsdWWFMDDOCzReRiia/qdVTuC9WI6OUWpJ0RTrHIJA5YLF3GU5CMWeqZYgMQiDum1n1W4Tq3
sepUJjUrPw7WSA7XbsOj53cLd4YsV6sa/jaRuT0yLfyNSOVjMdV7ARPuxkuyjRQmMgBcaGGAC9KP
1SZ8y6X0qF12qO6bl1QgfxKCsEARbC9T9h2q7MAABqKRIwRd5grPWDVtnBqm9YM9kr/x7ZuSLtXY
AIrIsM/WbnHScUwr2P3Aa1MYxUIN+WPHA1uOyZnxhpyhDf2pMydvaavVdZxdri69yUbnlVh6XCSC
ooktQYqN4f/uyJ0U/uIeTQW1bztaHfsUSw8n4/8bw9rePPlPMRcqHttOguvx5m4djymiZIPLPSkI
/CNnIAbZYb/Ya9si/30A8enHr4EgAxwTmlY1VKMh8OAIJlIFbDupg7pUJa8s4veAubCmj1kvjUn7
bB1I18hWefUTlp5yP2ZAVhgkH1sIc2xNPFde3yKG9rqaxUTOcJOgXKuHimnOtvfnC1FNQUmqBxJI
/BEBadLbpRKIKHeVNKq0MtQK3fnpUF2sAFltOvPGTax6sDOJ4Qsc2GqIjv+XxUQ29N4wX8W//kga
nXjYVE9oOClbE3ew2dUdjL0fUNkVZXm0f9bENKCurF1VFpM6VdhEngUou4PHbmMVw4vy7ylX4Cr/
MGzpmAeqScmwy2qCAHrJRCatL+sPo7HnSzOmGDWLX/03Otj55nn+BgCw51/iV6cVmsqIc1sXQfGA
Kj50koCMohhup3T3ntBvon++moZ1hKCsT41D2D2IyfydBAs0e2B1mBybWZNoW/OoF60pvxaTw1Ti
StSVSLYUtr8vBfxiDl4b3LqbYHoeG+HJeT1fq/9lXKrSIzezE7FaB5rwhv9jpf3aQzCOhyN+fde5
Tee+UbxaAJxcAVAqfiDtcx7XNANu3juSi2QdLIBRTeHHuwT6mOVYVF4laQuJo3jIJF+r/PVag3Xg
XutiFDQ4XIunN5KqJbWQJZwjam0BWeoY7RmJ5BRTgFRCvOm7D1xF4/HnxKL4AzkZ1T0CUaIAXRVF
yeAfXT4QWo17rZpWjwhEwbWk3KrFXrtDZSSyVUfksWYabVkA/4zQWDeJhD2NgM5Wepp7KOF27QrY
LcN+MNyYhtRGZt1vgs7Tzb1QKV0BxFfr842E4BUAoLFH0X9KmYWAAfdvUyZJTwHft+SvFA8ZUKCJ
eL7AuAZz99kdMQmhpnIJVKUp/MHevxYGEM+BEGiy4gFZsMxTMWhaO+KZgCxKg+cn+LAy3h7AdnpI
J3pDyON1lCCXmbRBY0wO8gdc3Kq/uOBR1GDPaECAP+NGduIEygtZNFvx0uePNXjF/0+oBcCTxmmA
zND1VswkynVh79vqClgdi3paWJ9olDDQhfS2DfYZotNLfgxCCcKA2nbRjfvys1G0gzySGbl2QeAI
6mkPZEfmuoiLG+xljdwgE4TdNQSsmiss6KzYH0q1qNn7j/b9fonMHHhlr8WmIhtucVwA/S3Ngj8y
4kmHG4i71Fes+uBUwgIhZ6i5wjRZ/3pbqoW13GV8cT5iwPfR0/3qcj0fbSXetuWre5ijRa2s8VQC
u1h7fB0Ftu8NVU1PnE0pUhCoQ7cGchbExvFSn3yUksYTiQnhVa2/D/gUWLUk4FOu7ZWLZ5KNBr91
tK11wWE2uNjsIDmvKsGMPGG2FRCqKZ2zRbJjdRDHrTN1lsVghAqbYsnvjtxo5KWqbdPbAyWsPTUT
+q7Ep6arJ62fBEU5nA7rk53yWQupiQJATJg0QnzqwJ8O39LlcFQpFmOelZ5ozsuGdwGaaI43zsaQ
fEJl4lhvUYc6/0aXBymqG0PkQJtd4yQ2pBdXvVfvj46mL2TyAHSCI9YslGtNLeenZi78+oukForn
rsLC9nleTCmBq4H13f7zTcjy3jMwRXnQz0HPQy044XtxcyEiLCxbuMsKPUzfjcwmahB+WPSGn6SW
3cYILJDvyfRafTl1NjOJCgslFgUkuBfNHpBMkvOQEiIoLkLXRjETA6fJJ1+alFaTWdWW7WTYtSrE
M43T2p5T4eutT2eEr0T1MwFd3fOrp+V/9U3UWDCt3IlA6kZeUKFnZkV/WmI5RpT6xwzdlkhkKJna
5wdMzSlCPEIiMqEwlfZifh1RSRpNKC1u/APymWNAIhBwOjOVnGjrB6+rcnHEC/p8bxW2uFEFz0+y
4iHSV+0wR64gcHgp+ccEGnLOJwyLcoP+Nanf/gnERHJnK9bBypn1sVN1xTXypX1qH+TLELmfdp3W
5Iile8lXhVfvZc4h7UtBUudByMArzr6/ZpwoWvkgkssAg2mgwiTS4dg4XhDVlVfhBponaxRozjBh
jYWTBzWE9AwdUk5nCqs9LQM21IiQULyaoPJv6agAmI+Nx0SvNsj+S2zMcF/CF/QIHCmwqn7UzzVo
r7sVhMxzoqcZlaXcvMB9TAfj+8cwyJkpkdSVdC7+k04EKzmu/roLLe+10xJZgUQwpaH62cprIDfI
xSuuSyVz+kHPN8Otnol+O4JcXYexHJi2L8EaYoQsaMYXUV7YM2e69iOTc59fhz07onICaJP0OeRD
7uM28ZFPpRkpT6BM1j+FRyDeIEXPYiGkLAogAEQgdL6usw0AOBwZqsIHUNYRsKbinBSNkjhhmRdc
LPQcNLyGincCtSgI1k0bXtdROJps7g6fiPu7lumnHrgrKZBbap7ywyCKkUmftNnDjbCbxiY4jvOW
VjPDqN/nr7nWm04vKByWLVCtmHqa8Xefa9qX5onLtxNu5BBWER27BPK5msDMbxFTyL5K6BmLomPK
eKHmuXagWmd6zZmhIk43YnSR98WFbIGVvvCXfl/Fx5o9RuHTz2AjL/gp9oYVbuhRptMvY6bdgT8q
ndBBNzcN5HMKhLt18vxNPacYbX44jfYAXE3P7x4IYMno/m+zql8XCsTrpxaYVrXxA/ovBnDbPn1E
v+xtIc1wPdk+cRu3ZGmZNxXJnThIQ+TuBrSCHoR6kFgAkyvUQLxxi/WEuQDadfaCASO5RJgEEfnq
WKSNVZcV3iMpxdTditKdNBXlZaI/FtqiSC6gjo4Ms+JXViNpcgIc9JmsDFSIM9zS2wRUcVCol+t4
aUbwM0RG7cfukTSnxfykot1iPgRGywbj+uxGJLrF6JSe8FXqbG4s1WCrvm5Tap5cN3xpaTFQESIP
hAuAhyukwkteVsWbS873AMFI70T+3IqetXTLcMYbO74LRPdtzBeKfwp/M/Iu1jek1yVnVx6wt5ZR
caujjBHrscQYMcd3Riy45XJh5p1H4do+4kNVJj1cyGD6jiCArWIIQpQ3S0KvidAdVjf5+IIY0QLx
aw8fTAr1bby35qU80pzkL9PjlYR2Jr3/pshlD9otXnVLJpUnaNWesSwmmdtS841nyCe7QJccEeKY
QQKvZXMAWEwiooY4ozY+WuoiAqvoAiG2WiHHnDJXvy2nbx1kPMCNO8UCO5ta7+hn8JFE9utJ4+is
jOrRsI4i3D3CipdpuxusrvEhK5TBHaBBGKEkc+28kybaRkwKmZA4HHmZcwROjxWsRnutfbvNwZfn
8n7iAZUTLz7aU9V8bBYkj0xrgoLz0iI8s/VsLnSXHa6LEUBYe0gyyDkYyIIwEH/WAdGjXSHG9qGT
IEd2g1X/Obcyy69afzsVHeyOta0ASWf9eGkTXkJ9Ycbp2MthjyMl5nXHZTy8W1VSjM0cUv97T0fh
DGyAzEgBalyUIEw1gLIpQs1SOfjnjN8YETrK0a2bmpYM+5Qm39N9M7ZsR9yAjtQgtZ9ueDxLTQoH
3eLiHJn07/lZw6qc/Y4fsTUI1GpfdsKARxm0115I4WO7SY8iAmL4zBWsE0KjEXNXZKVGbBl06ar7
e8kKGgQzDpz+3n+uJ9st2CSr5C4rrQ207BqQ4r1Q7MEjojis9sbCr6jvw17GDYYFXzGbzj8/z8SY
F40HimnUc0/nhQbxmOgPs2mlL2QlHskdEASK+5upvglW+dkjVs6YT2kYamCSNIMviG+OY4DDJ1H/
iy+mRX0NZ4VrGWdKzckRhUZ3D0cjX78PBndjhZFY1i2w/W7DTxIN4rnfQg4/bpwfNzMQd0NVm/g2
RBomcGOx0EGfW/di/S6X0tgS5ZjQgoq2nOWsQVPjQznYiWsARCURdgfEdb+EOqFZ+Lg+6mUsfeFc
gtxvjFRIQ2bhbVRs50atwt/ekIE6+n8M6aQXgjA8W00OUfVbyHAf/I8Q7Cn0vcuk9wgZYKYSWZAy
yHQmKxmyQp7lcJ633gjTHEnaFe9MMW2QmlaEyEYdayokVOCeYgsmJT1VGegBaQcLWf3vbWnO7NlF
jh2ejiu2OaDgzcvXGAhOUycpcIZ2EHgl3SNwz+sJrVgb8UGmYeRIbQyMMY4W1GLvwWlzQYXDxtaG
j2Ped5amI7/F8J4WMB2+vdub9usfjsod1hpyr6HFjS8tdHmGRavREGpo+Wcx+Y+kwuBHRDZRifzx
uQjwLuZREU8NfLLQfmHrVgusbxnV7Hh2lYHX1hC0wxMyDCYywqC/HFNGjEx8UhLrlHuwtro1Prp9
70281mZgp/BdF8hmeeWHn7WmQz4CHkA6d9BzAaZze+T7S28uWWyv0tJJQrCfVD97vBbW0B5skQXg
UEOzlCfqSLBbrwKXcwsxOohoToCD0xLokRbkoqHqeKaBSyx2rtkbr6yTKqnh6WPOnbBnetwDD40y
oFPyZFnxZYCq6hKxi9iTtWdL/9ykrAqU18UyhOkgqVKkBo0gfiN6q7APFzyl4Bzm6gwEekdCFnqV
3w3tTWuPlrTWRMuDPMa+z9MJVpknIwxNXF9/j0lModAOoLxqmhBru7n5hIqbcSZfYumzybfK1MhI
H9/J5rPvljMbhpNnu8qxRBmbxbfbHkdeAsU4OgIOuCFaK2k4OtNXJSW1ZEtuSlOD5nKlWFkJtzBm
lbXChCdBHBTO4tgrt7bnJ24KAy+LZ2RNFTpgaNDxU9rhG9ij96hZ8kYX0sKi9KGNDt+Fbc0POaUh
CpRbPPZ9rY/i0QORlW0Bhlvs0LL58EYf1p1YK3sduy6TRzYZJ9EpSBNWCzJ6oFGyJ2D4MH3yRNhI
LWR6m4SVC11PP+MQsxwqaE2oCE2uFThXWSIM9QdmBvtllxFZkEathrS2N4LmNk7VRasgrsFR4d2m
dl8/g3NZkKn3aGFkVzg2PJOCAU+vo3x2o5PgGOI3pC1O5w0JEAz3I+4gSOT1ediasuhrIST4jIWJ
+++5Mc4CgMjJiSEfXFrcuvFIq51P+k3d+Tl67IPcrJU6zs2Ctc1/CXJH0jUmkvq46byamXbozW97
vh+pxCh4BiuWK9xEHaXTSa7JsH9tB+88j9M5h4HThA16zUfHSEnOJR8o9zO2GrXFbi11d9kCI2Yl
Iz9ZAyczy7ZT2g5npItTlhwddheV1XeHz2neaLbrsjE7WjSY7a2ADa9cKwTZr2DsycMO8HET8fUn
/6BqVO27l4sUg89isJt4eqBRebQmhEAslyHcFNQazmT57ocDsNB3myOyw/2bsSiir+euMqdjX32I
DzOaK60v5tPwRnXJsM4+I79t1o0nyVyxxGJddqKWWzEBEqlm5m4R9O1fdpF3c2Go+XXzsAoIxV+H
DtCKBnipNS+ZmGC9EW78GeN7ucKYHyfEbBv4384MyJiaXPaEMSpbGezOFWa1nLLGVMKXxD9Z/1tO
4gem+nEv1dm7JH5WNG8bUgBQVYtI6Q9LNhFcwikx3gE0xla27W12T2yQEScAssHj5dxAZW8CVTvx
DQLJ6GClC06AOo85W2t0GaV4YRgWcab/MPij0QnrIOVfE3m3uitHpVd8AMmLqmn08MnM19QIZ1e7
yqnqW27RYJ/ZNZtLoLLfpMvBTPO/0XQ2tTTrYiwyFNnbxkmKwUKbd86d2DR/fYpXg/sZKrnAZEJH
L5QJndWntfryyYq0m7oV16ySHxXP3Pnalh1SNZy8mDjJOnp3lrdubyIvUgpeNmTJY5gnxsHabyQX
N2OpWhhajFlb9KvGxCHDT6Lptw5vUbkYJ8q16+j+SmjGVJQ5JOaH/hT1j10wcXXO+Bzed/pSWxVs
zkazE7zH/pUNkioSVvfXGIG0W7KLpcE42DzLnYH88nJylj5XcV/hB9rYvX0iaP3szNr80L3aa+8Y
LbIQX3MrNE+U1aZW8Z0bkaZ3XIEZ8MbIDoNcYu0mgVhTYExiPUKuWRz6d1KmZnmny2OjzTfbuS8G
uIdZq9pHr+nyFQnHnqQhcDLogZ4ymyfsBw9vdJL8neD1IeGFPIZL9t+BXxOb0Sx9+BCuEzV+/9Qk
XUX+xX1UVxQiCcAJaBJd8aLB8aHo8lCHlCSaY9mTxaJlc/cupx0hLKiUy4YtUzvwPM9sewCK6iTf
xtJ28v1loD4b9/xHwvJrOd+GSXjnc0n/gAcM9dLEvzPld1SMRvPay0OZXFH8m59yyqHcZfdR95S8
4Dd9q5G/NoIhpdwk2TNLVvt33/NvZAqKNtgB4mVHR2bGGViB5fQKCDbEJ2NsSZhkFTNwXkHe6Oeh
HuxT1kZpEWSFCttdzuHxbqi7PwQ7RNdSBuhLRdfCRd6nwMuAdbRM9H5I3EK6Z/InXYLzifpQ0zV8
EvWtgNAsGM++P03PGMnPvGaJz9lpGua7qzOaOqdzai4rt6Hij+xFW+kIGkVr5O8aCi3Yylc+5ms2
8f1tVu6eSPAYI9wjhdwAOOOQTS+Qh8O+Dx2dM9wxJFF1sGkYi5KXIMOfQxfNQVDcrYHpuViv5xnB
GW5y3f17yfb8mtP9L4hZO+0PkcvlXGygbMGgdKwN47IvnocmdXWJPoXRaNHlhUYFBF3/wu8OOzHz
uH1lDgZgT59XACzXJIM3AVmoXaZ6GSCeZkTXe4NduBqKKuCF2tSQmdi4VR6q+ws7jPy0Rl5lsRUC
azPPd08aRwOt4Gcnxt2pMcDUefV67vkshIM005XhMoeUodxC2t2O1drciANS7SPLASdnS8tiWuPZ
IuNG+sCGHqZQEby35chtN2ZhzhWi57m9593TlGB0d9T3u20niM4ZaCAjsieJsb3QglS0xt/u1dQX
EhJ2tqhFtU+zj1oQ0eCSrpmBBJqlLkaaCYH1BGWX2t+W6rOvl1zvzAbg0QGRRRzp8Iz4kvQhj7DL
x01/0i4zvNWwinoCZ5J31ocaIHoEvhTCXj82pr9rxih/VoDqvUwWNK/C4h4aRAvAp74oUK+xt7nK
uKkndQOExzbo5AMQuq/GEGz5tD5NB3TRc5fnAF6qwoBqbcqqusCE3lBJbKfLwuGJ6NS7grVez04Y
Crs3KBWFpw5c75gqukKRDthqNJp+PMaKC8xe+GCsVhHFD9O9GTZF7Dv5PlnFEOI9/t4UmhG1ie6r
wfTW6gTK8d/Bk5pFbgoJnKQKe4uMdKRtntCrKwCUdetR5UlsSIhsAO602qtFrfOJdnxsjoCl517W
FeynlPC5YEQBLSovgcyWnPga1YYDOFJtutiUMHyzmY1H225blBd/tXgAqkRc7C2S1D8oZyzMc0tc
8/Jl+IfXj2Dd+F03qaIqmvkBq0rpVXBv4w9wcgxCHrrPgo11+BaosnfxsxzcCmuSoBIqb88H+hQn
Pc7Z/Nn1uVQjM5bDpC8Z4kbhgYWPx/QwvFOUWCfXHjmsb+dpvvgHT8UKGDWgj4KbgEXGkvkBreap
kNCy+jMUqh+kUJlHIQMCE+AdzjBLDLJsT0TgoSYUi1GXFy0G5PxRGshPn01ZJ/kp0dWvFULIVgrt
HOOb6rXLn8wpZB2R5r5aY9J5MFzsLS1uJXncfqJ7RyHljtMS9eJk8KgBGIKjS7wIjWz3QBcPkuaw
Z61bKzWnb35M8KLH+D8vE7vAp8a8xVq8REbfpKKcX8FHOOXO3BOctXRKQ22z6p9HfCs2Z3n6Foit
fMh45dPqAb6yrPh3ywbnGuPjtgtpxGRg60XBljmHNR3B2wY7KPiW/l6caI92h0wBf3WlT9XIPSAP
hj5US2wEBa9tPp/HxDJmF3KVXqLKlko6NFZn6MYTikSOOcRcBVvIff07y/xrutlOkzrbcqfndD7B
N8s96HEC3OqF5pTbYEdQ80pdDmbEvN67DL6vxwQQDVislSy6yuA+pgTLctqmkJ0YYiWAHxIijh/k
wEECzlBcUfdj7M0YeVUeqrpAZ7iwt+GeH21pV355LtMNtV9wUoY1uUKdmv90Uw2eB4ooainBTrz4
V29i0F5Lm1upa1+D1mNpr/xGMDTYhK+BlMtNkGi/jx9kdiMWumTZWSywoyVT3w/AeMoghUANgOff
hsqfUEeAMEQrCqMmRHjUI/f+MczVS+QUe5/Y8VVwUaS5ChbKWzWLTYr+8lmXnocoE6RothzPqIk6
JMJuno2crI7/IlinQNeSw1YH/Ucl6Ho7Aud6W5KRNeXBDSKoidlLf5jegmzuL8OI1NWPItlNuQ8H
tq2uE/73TkjiZ+mmzttQ82s+YN1sOdzvE5uDqclOCrXbu5bOZf6IP3Xpx52AXaZqE6uhISrgcsoY
Tkfgo/cZGrbFMV64+svnIDq60xqVXHR43Uo+pBR0Kl7lkP6XlgpYGMNO87TzKFk1NIrDXzEa7NVa
RBaG/zguRx+kBksmMaupIh+FOh0UZ4yIo17o0nkPCzPHHIsInsjHA0JtvTQDMQHiL56ztW/ZmHnj
uvh3YDyTlsead98KfWPrHmoc7NUP1ozB9Xtzxjya/3qLKSmOajBATk729EIaHfChFPXgywi6hbUz
f9i1eKs/ZP/a5ZbePsBHAbYHlgCViNDeRokX8hsKqqMr9VOEkgKCIr+0Vhhtfuwi0as58jrc5Scq
BCJgahCjQ5Jngzghj0d5KwR9EUcJInPo/xzBUzAMga+XATYH6VTW8apwOrZ7VTzNiVIlfdy1HDXw
NeJZjexk+Ylx32Dqeem4rKC5hVvMGNrhBQy+m6oTlp5fKjxXSaBZx0uy7CsWGbQOSg+JQAnI5CVp
LX1kU4M1LWNjY8TUheo6T3k81kRjf2UtQ2aWyF6yYPrHzx1IHF+jjuXaImg/5AUuTKQ/eYSdXcu4
x2P2Jx3dyIdzbXcBk+M00WhF9yiHgn2EWpR0zDFkdhjxf6hiXLY/xtuyTh8QQm/5pFMO4qYoXpM3
LoKjf14bkXLoWSYltcIelzt5Eda52oBke8TSAmnVsMY7SgrxW9mIBKhBVYUauT1lsRSvUCfvDGBQ
OfhbJJEJcdkWBISZHRwEpTIxIV2jbn1HYmDcKqqQ7Pgca1qVPc7pYx6Gt6fRc7seT7xElJvCH99U
PlAT6vyoYPNHVCm9oFZaVuRzeQN1Wd3z43BTWmu/Aj5I5wr5ushb0kP1T34fVwTiQpM4VESNH6Y2
sR8uB5AY2R6vOeN4GC4bZscyjYcmVHD4fVNfj8VnoHINNPRRRyazIwGSr63i3+/66kl7vfY3I0yR
e+nHmZZG1TWtaXKRT0QMyTUBd02DH/uXqcBLgh2Sw/Wh1z0LlzkboqxPKKaYgFL8rXgVVdsDNfQO
GpREr4xjSNJJGVoRCNYuBiMa71pi8U9UGJ6UooGGD9ykiiSiCQzTrwL1GwnudX1LAudNRv9JdxTR
S04S4jphLrDeFFbQhTPn0bTtiJasmMoVIRPkeBCDSJG2L4ivcagY4k6DV/aD64GQ8dg/qnXt0dcT
aL1RSJb/2gRbMuvIsTCZpbnSbd1Km4WoAjsnx8Cd8UN9D+4ZIyhs2iLFzLbof+VqSOjNXOpsMn++
jEz+X9GS4cq8tiYayZhDB7PLXE4J7/Dfv+hdrNYCfsHh6d4GzZ/X6yQiXiIuG+6TV5MhZoQhS/OJ
XaHfRPeY3IVsxzsyi21uNgSQb6YhNE9yRUbS8thrqff6ZuwlT7FRbkoDyCyzrQ/50bsJ7+sOwGnq
Iz+qvN9lr1aprCgvwS7xFq7DjkIXUBLh9vD56SCeJcWCjad6YXTaflXcpfOEFKnWEiOpTfuK3/9p
H1TmAaYogV/0OGZaqUQA/FVXd7VSTwIdD+CJ/0uKKQ2PgkVLnI5i0rKdbsuPAzjsGNs2XPZr0UzY
R78Nwh5JQM9OX8pyjCFVr0pzanB9euY9k1BeBvNE8IBghMVoZQC/nlUO6GBHjEexqmK5qsxk9z0h
lS9jMqNCAehDAXRnC7IWtZguJqtW27XdKxfSxAjm5OP8vvCLCnFo+dYkwP1NaZNvhBd+nc3dJSkV
L/7v51iofzdob9aWCOjPIcQ5c2GPtc6isfQ1P4ajstEdUYiWcB8I37jMsugkfGdk4DCHQg/MWSmN
rtjquvKIOTzuuN7VIfTWxS2m6Ju/aWSx54W1Zhi7V19TF+lTjNBZW0WY5KdvJ5xFC0bfboVAdoVl
Pe+ASK/5IHFMLHoy6tiObnTC4VHqTCuvyCYuwC/bj/fiek8eGJzFrAsE16pgrbb4/krJMIYUFvFg
Tt6gn0a+txAFZ9JQ3GRCy6w7q7naNnTwr2VCm+6B+8HUnDmyof+I+wbJKhNOLjmYrAq3ejBxeWDJ
KeN953ZfSHbvet5AxlirriQNk2IsqhzaP+bGt/35+arTQj4c6Q3lzS5MJM+Ga+LnLeWswmO/se3G
/CxcjfAnPOutGu6jhrJfqe0i0JUI2azUs2usM7xcPVRhI17s2zpDazOulVYACFS/bEt5WwSVI3Qz
VmHxbbF03Myr7pv8g3D+Pm1zEtvhg8RJmt6hgOfcH7xjGmq7LwodBNzV1g5gIoj6jrNATwYZMn6X
3eqPZytnv4pSoECAtM6+84b0vz6nadwDrT0RmwPd4mu3HmHtxaUF3Lsj8rjp7grjAfJuNptCDT1/
5Nz5h2VPYQFcvVrMUES3EoRLNX31E+lD38GLm6WcYAKc5XruD3gSXyp2eXocNaUClo3w5KA624ny
JMRiUi/6Z28uObxp+WyfeQMc0TzgyJNhIpVRVzv5XyHeGbSM6HG68qZqKelgCmmx5z8GjUYYRD26
Ft5avA9A0cIwcXMlPkNUyou+2CCti8rDHyqJIXXS09nSbr/H9IyCQfUCwfm5CW1SXhNKtK/iZhfi
W6m1kWLpxQELItkHoWEOo5DLVN7vEHBtTeMS2oKsdtwmtifHKkDB5gUiOFPgRc3dPpVEBfTsLDYc
1TSvQoZ46gNy7KaxqQpFhwuFwStoH56MZ7wVrLc59aI5dEQ3UEQPCQA2AF/YrdUE158f2Nf47nr5
/YgMh6WunojsEaoeqin6IcUCTNSgSpEKpncgUMOaj2CVvd9p8FmQOlxC6QOFG+Kz1OD1X8QAg033
XpAO4B0aJeHU1U/TbeNIJ98C4Dr1GCg1P9gbFEp0Z8kwph0FrtFKty97K9Igu5ZhSjMQSGGUyTIz
m0HcoMUDcqu6uOJiVhZdejPITMt2sTvrESuEdMitVVbwJlLJn2XP7u9aKaRv+ko6Fj+CWEb8vcse
qMuH5Y3rOBCLujL3muA7lTciOI8eG1hPUG1xj4kbFE/+oxt6gu96wLnlE7pf5/+f0GP1wnMMoUBl
IiTDZX3YJIxyYHg1J3oQ8xOiay1IMjWNl99A78/dyqKuyDZjm793xi5TDtFN1xqWkP7zHG7xhcMn
JJg2AgikwnuP5nVOgMxDimbsoAO+Yk5818ipivg+FdjvzKnKIeE1xEawVUxI9RQngsf4sLrG98Qy
b/q9LlKLKLdEOBhnWNbhkMAJmziDEwqCHK9Eg7neFy8y7lA7cS1GIb/rLgVd8aYKksUm3Z0mlHPf
JA9zfzXmZx3gJqSP4rfH7uBOT1O4Pot6JYPRlALK7cnl0qxg2qhHHk1nPyKOCiQYyHp5Op1l5vuM
VWfhZBSCOx27ro5LmfAXMVdgPueqfDARrD23+IOtxu32RYlYGgAiwvyo81IRgGIzyvcZr2z5C2n0
hYQA88o2LqHx1wUJuPGx/xSKOckVqTzQoga409j0cf5BbQK9v71LauTSZJOWeQNoqAnFfzTQRCnN
BBjhRWcumFOOHXm3lxoUIODrWkWC3bEoi65vcHZnbzR3Qlkjv31HnX/bYzSK/9RycTrdbjCTnxYM
cpvtvPilZBFkQqahuHNv54WJkPO8h9XZhtJsZqz4x0iUMxaeamGhc/ICkTvxwlmDtUwRaZ9LVKQ7
+50JpqFmXWJOvsQSG3WVw+vkPTqrJiXADVKrrtV72cbSWmhDUKShgA2Y9sqLquTyKfxtgB08YNJQ
fz8UmYeHmxS6kcVp3NyUGA0omxTPR5ICs7hGiVk2DoOGy8iRdzA2aoDwAcNIs6f1SDbkPuWDin3S
Hvl3Ow3YvC7Ko9apdeOjKgS9q2VhqWR0bJYBD3jjh46UK9wT2BIo0xTiqIJPJUPPcfM8Qt5WAXf+
8ChejkJozpyvJc8IxtdSk1IV8So8H90LIJ+ckw39zv/m9J+jhCbdd0saPi7aQLDIh9cQTiUHNpHQ
Qk1q3enVYX5aX1CFlh06bWOKsCz9NcMbQNYTCJYQB/aK8o5WAam+ohmPJM3+ktKcp1r//hrx/B0F
V/OzW60q9t1CngT5T0/1qV9yGjEHYEbpx3aqXklsTlv28uF6VN9dT5rAZF1fPfLUhlvxvPyhU6bL
ee4/Mg6vnEqza/XtD1J3u/VY7/1fDSQovo62XNhbBFhsoUTxU5YDRfcFZ8AHG+/l5N4HKbXysrrS
Tnr6/BwNZzd21JSqYxwQ2vnXrOcqzdfPo7jqLe1vgssdHtVwUSLbMdrsnII9Ryu/Q6XIZxUFAHSz
C46tm/2/2prLJDLM6mCDL3z+zsXhceDnURPELEkyzYAPeBA5h/KiN5Bs2AecNmLZJjxlJpMkDN4x
56Ph0oUrV4GEICJ8rIHF8nXGY4TrnOC2yPQPC0UfMqzH7XZiyIZQz3w/iAqWsFXLhIzOHaeDKGlq
drvl4y+9cL5CnlvJMm6ingaGcj0+K7dVVNVwePG/SwE1xUAovFUz/7mIuSbst7zCnlgX/2Xb0aXY
SK4RDdyKkMpRdVfKro08bORsP1x6cN0oKsZsXB19TOIJH09cwdHQy/b+p3Tap2fTMvxT2Km6N2hn
NeFLWyecRes5VXbHr9ywDvfIPys1XV29kh3HxEN3SbJc8eO+Cgvq8ADF2rn+GgNKVdPCziElH+A6
g3UOaej0tfVnsInuPHUVLCKjFSGYb3hIW56nmTzpdjeB75Fr9nf24Vb8SZBdzskxrH+vBhxuc69l
ftIT/l5eTj+WqOWWpOVcRQwiJgXk8rHhP98GP5URLnU5wWGbRGB3JvaYz4jjtE/XU7BuNdMEeEsW
K4SG138XCVyu9cDB2+h+gpEhxFBdotZmrH/QR3XQ9Y6eh2NBms4/VRvCc0t8fYw+0rzAHCFu2nrU
nms+e0NoKu4G+HSZLIOq+drzKmazKph2spApIrBEdYACAlXJhtIYa840W046O0apzY4iwxgzuQqq
CBXS/469/qfTDl38DwowOxFEA6lylAJv6G+jj2pIZ2+olcASu2HFe/3r8qJ9huGHEBDrMSXT/oZ7
IazsVxBD3shpjbvv1FYsuonk3SiNdDyGwt4umZjo7xj9pDU4uBFuiptAtC27HAkBvf/7wG2yoiQ5
iCbguFL7kGow+E8nNi2flbw1SDI1DFvzZx2t2yq4QUTPYD4kgUuKFt+RYvO6cQVjXBSJgS2Q1nbI
9wp6575XPJpdJOYOsVo6CRBsiyIJUk9gQd1ZZzBrJ98wbQ81fZv8Mj8/v0+3cLWUUORJ8Gjuragw
KpnZ9IyqovVKaY8fEvNzSkNBLjIPreXKYDEFrfSuMMRe2Ms1jzYo572FANVPqllbhpU/kN8RqEv1
Nc9Y9Ln289NoUdVefyoSd/nQqaCSFMyESboO7qkJu0OYAcTtjlSi0ccgBcsUbmLwQUX4j/pBHpBI
BGPoDIFywuwgGLfrTN9j9I+8eCjyUxMA5yn5zlxsOpG6eBwz4lAnBuQWc2t9gg+0hxXZ1L4iwpQn
RvkIC513iD/RrhvetetHkOlRAZfsL7+9SNHJSZYNJFN7P/1aX3Yt4d+bupJ9vbH+w9i0oCf8OQCM
qhEdjIqmdmr4YfCDhr19X95h+CcDTe2gedZEEThS9+HAvKprrRIHo8t+DL/B2+6z4x3FAvb4gOGh
0Y3/lSILGgjeBss5v9lVelFufxX2fqxLeHw/uo2D9HOxKrJvF9he2WJ4XxkguD9zMrydnk5WJgxy
1+/4Y4pRE5ZWrwS2KUJY5jR8SKi/6xtXiJXa2Ch6gJ+n+sypqH07wXZPuCmVCRdfx6+KmmuOMQHB
crNTVMJylfBzsOBUWRKkx4e5Ui62EQvjmMTJvswtofsByQeC9DVLlH/JTk4r8hmoxeTH6YAzlEAE
+fNkJEQ7MvvbGlvXIA4ZcHen1qGNPIFhikltRdhjx7F8gNpS1YyyQfyaCJRiFIjkWv7bfZbbLa8o
zs5hOaK2/zbPZRduSiocByMojkDCBXmpPX8Jei0hwhxuB7X99BqCz8QidKiwONIv1HBqSSuqunI1
kZU847PGz95rQ/l6JC8/I21RIgHrhMZcILaQoFCQWeU+RccvlOEtKq6baNF82t80RcYp9/KiSlEl
fqM96cf/u7XjMMR0+pJeOIz55O2ftguSt5RIvKCT/VQ/K00pMNWYeUs9h6v+Dc5Sn6eNuJwsBXuG
DfCwuYENX/2dPivDAnsJP2+l6V8YkBH4Wrt41bd2VtQMfnGMjCRLzbsBjHERiACUWku4CMUTDh7/
wC00yeMdVg9wV9S0ditULQC1WjYxBmzTjqbk+7JJUpT26bKeOXOHVoV4tJGHDo8MPYBxHB4JfO1g
LW2/Kyjw45KCrl0ODCwAg/2vLirXJnGJsPoAGCBHa42PNZZx3jvvY6UmqMy+LMpEMAxV9xDm4Yat
+YLd1C6oNBLPpAyWQSt/rOXmEn0MSRWUlgOVhrOQngmP6spbdvbuzLzSutymHvJWmIaRzgV2h2ia
FdJZ1UgMdf6LOwZ9i7fDK2r1AABF+pc3+ebku8KYX6qHaxvKWF+iPoWvOBIThUgrdyENdLCPJqn4
3SLPgmVecAI910BJ8/APPMnjbtPE2hPDq3pEk/hF/605HcqwsUcyvR/DIv3VbNJmd7NtkVWKP9rc
LnFsZ6qRnQ85YToZY6fdidT8exn9/a4+NOnxQAPJNlAksbq0r+PO6/hLJabOXNnSIhhopQIa3wo2
tyAq22GMAxR/1+OtaPzBb5MjvcrxbN50jkSW2q7RNE58yVJrxmiR2ecnlig2pMUkTMiBSk+gya/R
6fGBiGZWT4JFJaVXc82UX+uU+RLem8pE3lUO4+HCFGaKpqJCcdzBAkhhEQkakgYIhZyF10WuBaQ2
laFvwySLVYZcfE001ikxU0jrbDgyDnoQaFCPTmhsSnB+OCojNWcwrWZJ7b70UeBt9m48j2CHxmP4
7zrND07Ri9tbEX1QQb2iAPGQQABGGxgxsyfiDja5AbbKuiqvywTM6dIk/cW+ZC3xVIvg0b9p6w+S
5w5qzpdCqmBXg0f+xOcPdFoQSzV79H04qB1tU30Km5jr9T+ahn1qrTa3ytXgqbbfWUCTjij5E+Xz
qzs48kfwFFl1zl0Mod7Xiv8DwfwqsHjMYHbd43YAxwGxqx2XgrlKcaxlV6vVUyuLDBAFgD0JhHYH
ioYB3J/MEz8jUGChHf+nq639On0RhJ5Qbvu2F5EZxVuxNnVuhy7P0lwO2iDLfp53P/gx3nSFHFQn
rvsSQN/MC1txDvnh6+qoIuWBlDUwIQTcBsQ1jCQnpNZUOBlVLBUO500fJ+WtGGA9K3TLjJ1NepbF
hpEZySuuKrnE0rH1w8eimmJO1jJtNZ9fr3q1YD4SVNniW6bP6fEjSq5PkIlAR6Qu3io7y9Ri2COk
Q8LGGV3n7evhjLiSO7GxX7q3jydCnUZFtPEyLJIA6TbkSRwQhSRbX1iU+CIksgA30jfBVHuKsIT/
zDVUIFqyRgiQgeEYSGZs7cTUooETWJkhrNJhABUO4eVpUodhmQZFgnZIic3eG7iK1eGJRbI1NI95
zbaJvm/lUQ6f3rsC6/fX6T5pR3zG4JdwGgeWBvexVy6S8r0YsNQjzj2T+ssTN5v+7neaoQPbC62W
9e7i5a5qJA/ulfpAnN+LJ895V2EU4MtHMbS1SIEZk+0j5F9cIlsg2b5aWGtDOBRgM4yIduOa3N4L
IvCyKf4wh9dwMQdlb+HIGFU9GPr4tM4OSjZ9ycR/5SNjjpQJg1G5jKuS8NBwPhY9oWsaXsywYyaQ
vd4wTIDZqS00g+8Wo21tqnocbAFCic69VzuYku8csapf/JrIjgMFGNbyjHBfzDVahqhJoMtkZM+U
lGEvM4/5ZOU2cVZxnzX7cD57ER1caN+NOd5G5UBJKd3zpP5snjdxZG/aHtU3w7DS35iyyPrsTWjk
2w6t9PzYkCrfoMmY7FvOiMJNcIwTIiEUNy671bqLxg4FTGpROOiiOfTm5z/48pcqfEvE18Iti7B4
L0oUcm3qNoZ4baZ+gUYCOLMuVMKrU5YpmotI7VmWI9X8QmDlAlACIz9LNQuhdDftkKJlN/Twg7v/
6w4HdshNiodbUQY9Fi08ZuRiAh4t0pkYP9BgYqwgXxA0MbDFgiIP2EbaKnWdEC7pusY1PwoGdPRB
mv3QM54sX7IB26/nVW31FBc8YRNUrqT8KeqeE4oYDjDrS57wxIRfq9IFSFhT6T7d9vz8660+Hmo0
x+SFy69ez02nLQZGVFg7W7CUsXdlLGFC2jvno4bb81H29/kr1CGdi/m6UO9iDZDKOQi64Ot8RQUU
AbCmqQ29GXtDulRH4LBQR3WXiRZCUt36yOu9Pe2jN7V+KMoFQtYt2nnwkjCitweranWy2czc7mCG
YpQucR+Tt3bpJMi2QOMgAdRRSXPJqooKlIbbg+s2ZAqVtE9pGEaoFNpWU5xRxmyakp2o4vBppSac
d2XZ2YpTr4whAK6PfocIgxuy5/GKQ4JWNsg5P/r1KLlT/dND+NO6diMDt3ST8skprYOohBTNJkTJ
GpCIIkrh4beYhwB1zCZmeXnkQ9mcle7+BV8SlwfxW/QD9QO6q7phVG6Y6VzOSxeWk6dpi4Sz/Uk7
NwArIeZHEnkoHObQPRjX7RdOwR/qJCQRftsgDqbOFR+NwqZPnBEx9BWcdBQMulLKn3S/IW1m0Adn
FnyDB+rOr3kgy/wGRDEFhmXZtPEqEXOIqXjuuLEoEEZnJVPPcIZWrsbQeamYRuK6rIwvLhyv22Fi
JijxZ7hyiP4JSf8UvQiIK57jEWwXuYNKGziMepnMtsKGeA0M+wiOSiFGwzLuQsZEB8vr8/kOQJN4
DOHmP5WatXwoNLaDqSt/gkxkVlvTAyj4CzE52C8EpLpVMTNWxi9eIgw9OWlyPrbH5h2i76c2x3jG
mf17HXTx1cYRUdYHKhHpvWT7JiuWmnQUlrK71+vsq3JD1ektl+sl04ijAr3O1zEhHsSHK/bcJEHj
B7dUvd53WPPeSR2vDWsN8TPSo26lRRN151cOL/f63EzEJEOFwUKc/hLeK5YZNUpZSrOUsNLTPUkY
2Nqz8Q7/tFtulYWgIrgR67jioi7kxdUe+xaqX4nuju87ia78bFdnOB4CTiAq1LfToireY0utb4FV
AROK7ST2Tb2VmwJr/kdH5uUzGPHIm6xJRAW34LjBOuUwFns1APQy1K5M1maL7dtOVSAIM/PfpXdb
35jFs0ZCYuDicIcOfN14OEev07CeqkGguky4y4d9U+T185qW4dE7gwg6tNUUIexWF/hZHbsXwiuA
eRDBy6wA7UldiCZX5684oL7h7GB4pM/7vpMpU30Yv8esbvaYECCZVdCy/mvP13kyft3Q/vxuEDdo
d/AeNsu5PgfHTLIyw47ybNgVexRUIKfKdyziSxJoDMkwoTLYKWDH1dkKwHX5NH8/dK67cR9HHawi
6OT0KrMtC2r8BP2TJgbKHUBakexbzXgIo8IIGC/T4q0mgr1SV6nzaXbbzvWRbc7leUpYuKijgaH5
/ptr17d4hhmO9qQOt1YyC1m5Imsqxngp0QnDyus/JVJOdSuWJ0kC2rAHoamUQwpsX2WK27N7OC2d
gWre185ao5lgmoOQ0NqNUnIfzX1ga+ldV1OtsJDRzwxwPgDHqbmtQgenXTaZGdQpdRz6Rnaarq6P
gAYttfnaFGTXg7o4WI9oFciYNZMU5cK70gpfDh4ZHTe+slPxS1II1kfjwnM9cvhJRHf7kR8e/o5o
3gqTTyT5++1pNx4d/3qy4W/0FgqsNx2x6D8HZ/2TgG8rQQS2X0eNJn+gbhn4f01yz6hZIf5tvrAE
Q+GkHhwK/DQyFdcfInoI9VRVlvWOeOlDP6GWFRGWt9oKzx+zgqnsEPXVZtHRyAKoUVpEgwSX3j++
dF2C7weGHLhX9w5WJBk5IxQ1gOu4ZQeft9WLmdrVqLLuQMPNLVkM6RHdLfi56VDTONxTwAqwSgpE
POnQv09eFS7sFQ46JVz5M/iYKOpowWXRSIoXagM+1prJsZj+IR3KOgr2skqlbG0fgQlZFkcdlnAS
2FM2diKLzOEpseZ5t5PWANoAGpJ/WFFpOjfJ6nr/eA7Ip7K+eeL4/DmZiNgrKj2DmVUyZjBxSKD0
TIw/PY4RkXtXBRNqPNJM6qj5yuKpFP2nM/gbu/Muj4GQB2VVbJV2BH55lNCyn6oz8w12TB7yaa/S
GA3y/2Q9WXwTeOpzFvHiFaejidJgG+acjFZHXSVQqiGz5GjAdV80qss/WpEEPTDOyIzml19ei8ZB
LHSaMolrYyKzbpfSev4sGQuu9XiVFDgovT4sZyTFWlXApYLtC/XY4w8CwNqmfVbP8jQuZbm506od
582YGPy1Rqtb+wedQIu484TUSyjfaztjNiWImHVV8/crt4UcBpSkvDv0ncdtc06HiswAx4tH+MJJ
cSKZre+5SK26/TOkaZMYb+uWxe+PRXxhFMhMJve9G9Z8CbeAoBqERDfdgo0A+YehmLTZQX/+EIlZ
1l0Q8q96VR8JLoApIRxSIw3KfMtK5IuEtIwIJ9Tuxv8xQXz8fQpax+1PLSuG9+hHtynGYfXYSHj1
ZCuOXrg+9YtXoP+Gkh1dZqqHsWKUUz3KXpr9xdgLEUu+e9lcMQJvPYBiBEeA7gRDj2qySon6w8EG
nUMNUteTyXkK6lAIWuvJFxVQaJUV0kGyFH4mgcok++LMSkz4pBsjEkwOtX69DwjPax8THgskFWBD
J553mqVew6BODjo1bBaw39rYcaMkBz6DLR/kaftZSpm/4eT3HYSNp5jdtuxhs3atgaxw+jBL2oyk
hav/8hXeYxBlGAsgWaOQmGdTpqzmxyu0lEOycdnAg4DZwCoLag7NAbR+zOYpbqxwYvwOEBN3xyBl
y1kReWfGSglB6OZGZqwHfaGGi5hSzB/f2RaecpZ56zrlo6I0zPHbEarjBlZofurZpvLXDdo8Y0zz
vVoP8f2fG24z1Dfdc0zADnZWoq08xImhUp/jCdlffhL0YmipMXSIavABNINFDwZc4ix4hG1aA3tH
o1kUEgYgPiXkNXTagYs5M7+uqFQTt4/HOmJyygyBFh3EveZtAryECJNb0viWfJe+um/NXsVFY+sA
ll98qpu41lfuagLXbT559KtCR+BytSd0vfFU5Y76VXM3qM7YtjS+lR11tiTHDZA7L6GH3oOP2l9N
2tG0d9GfISrzj5FsugX4DClAoeYOwYYcTx0cKvvAACFP20xAqb96JsMl2G68P78+mQznbxNp7rk/
Gj0WGprIg2QRTBUTwPQoZg/5sA0prxUO45D/BN0jfvWeQGf9xhvX0sheFgZ6k8fuLVhGm6HA3DaT
cXL+rbP6BglbAJ5bQbq6kSyhL1v6j92Rs11Cb3gVufP9nTalwWfur5Tm4l6UA4xYly56pv3yghML
/xmykRuUpaufWVTF2D2ektmX8yHI5sdFMiZyc/kmJInOI2n2pemWNqBQ4KE/rmTQ9jOXSpchj+Pu
pyczFl57fWOtk6++Pg4STZfZCo9Ba3ivO5VlSGHUCdq4bWOONb+3848E8yn8DWgiDZvVeswHg54z
+nFmXSt76/GN4OR8VwFwqcrBRifGuqT8/+DzL0exASoe7z7vDlUkB16viMjCFEz7Og2g+nPgYIoO
vNVwgpf+WxC5Gm2BpawBOvlcVh434tJAsV3S+WdOMNg0mxMyzjNH6ipoWHJBN234FSospYviYWRD
AvjNdEI2qLbJOQAZXrO3A0UJyE0YgEutg8TzBIB11X/AsnJc6Qczog21bWPwrqRxxIq+HlKlCoVt
mL5x31GTLxDFrbDIR65Q5xLeIfRNlMKvIt535wQHX7/AnxXwnXwuG58DE+ig0VcpuTEwjWx0Gbsd
yqGzfFwwjsFOR2rbpnrWISiAdvw5EFNmcMV4xyo54FBsy8WTk8HvKZFGYORa1+oSKCGP1r4ZmQAV
xeWT0Lfa68mjNNehkSihybUc98xqPv0Tw7shHER2pddxRwbpKAFaA7X9I5Ra1yLlvJJKAg0OyMXX
EdH5CirOZHze7yD8WwPoS3xMhKjxmnNWycfK7jP3BHedh2mWptfBrgEEkaU2+dhIlcE8Hlolu62c
Rh9ad8zwGJJmWeXOt3Qvfsp7pgSw8Frk1LheREyvKWVTPULX1owXspj/EpgIFk5VnIxLlWW5qT4c
zRTL77xCkomF2USU5No1igf7eSrtR9tqs3tbr4KZUFArmpjcEUOS4qlEhlDrdhMqklSEA9l0E6Xp
VBcCILotWc94dYe9f6o0fgt5sni7Msk1wF6ySDjwHRW6FdQoB8+YNcWCDHbtvlAMfSArkRxfl43z
6XaFBtUgByJvv+fZ4u1iErBUKS7tmK1SXGhW1Ml/4To+lSjNvzSyAJAC29Bn7Lq34p07bTWBc531
/4i+xbx74GqxHjIGPcDTBmhD9U8SrYBof1TZ2GBEOir1gtu4mk3gkZoi8l1LNkLpF1oW+Y+NThSz
SiJYJ0nTbTNq/s/aAbHTSsOPF+xSpr/8C07ceU6J+nXMvldL6s9HwFf/A5U6CLBQ+W0UtXJhVA2N
xS91fc2G4V+RjDvSO8nwcdOnUrZIPfrTjOE7yZ3kvjpkIZffOjeZ2cd4SS/TmIHiLdCUa5vQMpe9
QREdLtmQ36Lgz/CTp6cKO6s3FoxmhUfJgykubJrI4lXxuOTeFnwiMcUSEoY6ASgzZekbV0WRFQwC
SLCHkU4S/P0EsCvh7ZEUJMCWcsWWv0WlmRQWsNSbvCZ21yzLygZ4G/oZ64Am/6ubfD/sjfX0+D+0
PJTGqqsLJBF59w+WnEHXUMvmZQjhK4VGfeZWkUu/fyVo23rfJo9XZlCBs4DnbtZsUqjzpvaB94sU
HfUyEvxlIud4H7Qf/YGI5vItuwcxpWDlMipljZawCcl266f3rq9HDmNjzrUxTGovvL9T/c4HPHxu
rlWtg1Gxx2QuBieVce2nltQbfxr1jhZm1ecW1r3k/SbtbD8dK3ffsxgG41Cpey+KwkQO6dKe/xM7
7IpAXDcPFu8chmDa2yfECUhGSSDgarKd5py54rdCo3z/ZPZDagjyDn1JiavDsKPVSh3n9oTBS3U4
40wvWq2u3DyJqB8HmXu07afYUR2VqoZ+mLgtZrAzy1fJk8WyQKqlUpzMrPkROIqFENPQL/EKliRo
i7PUs0CyUMLWKsFaQlJaRMo9sL5KmN7kWAAtBHLEw9RbIj68yUAtxi83npWvwPfI8/+lM1MoTzuq
Tk+mGjTfR4QNWsVOJ5WBUWjwoKmBgePElwqZKcu952fkRUM3b//UYMNcHjmSZ/bUhHZOBgdl8Zmk
SBQ/ahGx4OTVINQmp2tOTwS4W2RFrDKJTzLSIqHzv6V0W7WPS4ko0HJ4fWuLad4Ga7SAi10lmS3B
WuvqNQ3m81ygREMqQvvK1ePRTYyiWEXciEUW1C0JqjdPtCLXwMIdB9HCFfdRY+HLAGmchllYhrZ1
FwnAUuto3HVxvMxCCJeOT8uT6Je9O8OtN2UpgGOmiM9HyfY6SgZI/zGFG2L0O6GI9m7S76MIep4P
e+nPB1uQiIjj5BzpnRdawwkyujcmjZxCZyjwChXdowIF8SmKt+7sCj1+MUT7jxuCy0/e3/lJd2jx
KqRcTHMQ90003ZN+1+5Vxb+Nk3UrGoFQEPjcGLSlApImFoWem0ZX+ZJoBmmsYloP8ekiz0KuirsI
Kma4mSjMJfYNRJNkpks2KhkeSERYJSW502SL8fnVWlc3IbNmoJ/iwgj6xqMn5mylLUOGQTc9IX19
4fw7KmGDr9aD/PE5IWrRUYSPGvpUMCKBhKMbiRKeYAv8VbldMKYAz1sQEH9gcLcnTsEBRgUQDp5O
+WnDNBOXXPvz33dCuLduLKDSdKD9GelU2LV9FF9KSWAfBUf+klo/Hvq9nSroAdDRUlO4gYDqz6Zb
7KPZIujN4ujB3Z8XrpLLQoxe209VaApowgtmfP1Ro7M5GdoQglugsiHxVXA1PMuCQs+xhRa0NA5l
hVl+TY7Le2eJWtYQB0CEY+9BA4H+6qsSmhezA8NqYfLBZTla0jSnP94yHt1tIO8/U8DRtcI0CbJr
wBzgxGPojJHAWSab39dRtzD/x6pYNPktDz56IyiNFW2vqhulNVCoxC5t1vtWdtM0qQ0RokKnHSXY
gIba5Jp889o16IAThbeWXzG3sHyjeGqk0PrCXgcMiqUddN+WtlemUuXLjfsP4uvSh26/57FO9qyf
OY8+ibgHvcYUVnaPtXkh8Hpx5H8nrK6NEcZFAim0vJwT7Y/wNLjj30t4I51J5hWcpz/d+08i3dDs
7TFGJaOCS3DLuGkftrotHTlI2nA4ZX+dE8TvawFaUCqtnykvEMPWzJXBEdw0qPHVdSwXILjjQ7GQ
S9KCNvMUmj+ZiqAvynMtWg8cPVW1M7sn0PDBCz0CvoHuAWaWAAdZUaIvZnYRvK35qoQT8jCOR3SL
BCz9hKMJOZVT68Pq3zrhmwY6Gar7ROwrA2RUL0/imuaPKqSTvoYu50MedCrtY8hqjO29x8YosMlX
IpqMHJfMo6w4QtUW2T20tJVPFNs4l6wSFO4JfY8hOU0sTPNwvvvftwLZZpsP+gRUo/oomQoInm8x
dDjL3Mh4Q7KGqsRN4PhNB1JYXKhzoIt8fhkakNhP7yBkiDlpLag1TbgseosaELAGATyclJ9SlJxz
1dVipEDT0cYgzhlIBwIUYiJFTKZ7Cmhl/AML3FqNx1Fgwv5qYAcy6EmxefXyXzTBH8MehJrS1nmk
QCMvpOQPXXmaZrf2emj8iccbGznhd8GHtuPfbcPaonSlzLDtiMCLbjRUIDPNREr3xegdiwgxX2bR
UJrABAsEhB5psE3w5U1+j56NSWstVA6IzL3KS26UQEyfYCohqJcHTdemwy08BcjOOdZQCh3MKdR9
dyt70XajQYHiR7iMQ5e6hZuWuyzDbgAFHQe/r7iZQPTHUq+up7Y1ROyKjtLdioZK0+hGBzOQc6+o
wUcrhbSSYRX98bKXFLl7BQbewTHSHoJ4AtT9jH4IgJ48dHfUQYX0WbE5YOm8vj7OVQiXeIozHXi4
q3ie8JeAF44EI4nMS8rqw19Gv9q7fq6MDKp87AZV97MsO58hVja6U8VxxUD7hy1X/46VFQ7spq0P
r1MJaPEv5etq/WURtiiCL/j/HmZSX803USuuOnSxla7xNHpLEn+NzE0Lb9w7M1O18lizEuM4QCIZ
UPhV2vjeGKx5aj+p9st0cPjS8DIRLUEwEB5556nqe+LGKLCivg5BDy/O8uVttMS61o/V0vFjnd6H
lSGqXQBC0KRY8j8SwuCD8AbhIFXHFu/7942sXdk+yGKql6l20oLzKM+W7JxQlu/6/8Item2WBoti
p2cFrwHyRiR9JwhEvynaQfxOt24e0kGuljx+4kpJvDKv7lcgrrF6MVN+nwhaUtZETIUyOGFR2zpx
XEkagAFyKbmapjEl3Mvn9XgNMj6M095rXrlyjtslx/oqPhMgEe0gGjU6xwAl5jgQTbn7hyHTTZyu
3NOzeURx/S+UYoamiGHZcTLN5AmMj38kLVR1nT6w6m34rUKXEOCmtOgu2pb/OQXbkhxwS3AWcCl6
mD7oHoi/AbHpjlIn8cQpqoVgZTeWc59YdBRXKjIkKaptlUWRlpLl8LiTR87N5nkwlEa71/g4HJYe
rmlDi6U4FU8HMV9NPMjDu0YSg9Wk6i8pLFpbpa/Iy93zeTFMKz0YvyUWgczCHHdrK7EiPO+09ngg
aony1ij0LYIluERlXTxKn5zF8Zl3u/cz5Sro9+LNlLzrWMhmGua4Bn16v8NLvQcawi+kPbsv7Di4
M/bkoEhj6jLTr/cLy16gKXWoylrxoBuAdWM1xY8vYXGdj+t+KgbdZYK5gDxQt80MtwY/WvoB55+y
QnyzXo60aaunHAaGxihNEAkvHMfn2w+V/sk76tm0jiiodzOoHa8mo8U1IZCDRtXTRwBe5F4BPhz1
GNMG70KrfQPDILHCKsxEqdz4XNAGx6x3/WSX4RLY2erewf5x77/SG6iBU+fB1x3KkaIl1VXt4uJd
sEM8Dnmhvp4yIx4hUi/EcVWzxZ0gESuwaOMtIF1GhQe+WS8J6AdvrJWSN5NSvInckddxL+yvmcM0
VNr9K0YD+9tnHo5tM20g1sxyLyWpfIeK+W8TOxfQX+kz0bJEZiuO+1Na1caARi51Z+563FzRD754
g7xX5dxvYb3cBvVI2ZUa18U9V8sNzLtKeIGQ6ygnqJkWCwykEG22RXAbXQPP48gRg5XYq59flXsC
ZkIiNhR8WU1/ODhRPsIqL9E09fwLhljpRdEZUAg+FcWXUgmXsbK77Q2JL01RZORkdRhvQU5BUjPr
PKNsiKRIhn25SxK0D7KRXwQSTVx9Us0dQYx373wMcZtXsVvGIcIRiCThfZ464F0YSoAVbSFJsear
aepDqD0/0jcGJwc1AoMENsKb/B2/L55c7DDfMqe4ZjXrKfSSrI401PJT5/LsX5j1I1xfLNcK1c2T
is9RJhcEap2hI0LuC94hCIUflAGYz8GtiUPNwfqqLSDJPRHjAeHyq1C6HhyOzOhQdBO3cNA15zk7
yajSZhM+JKse4ob5LfAeSrYhjsyB+BkeBOcW3/unilWH8lFuEMKz2/QVjgsH+DZ+/MfLkutzDR9j
JJBsVYvHrDQJyzRVysxboftp+BjZhNcCWq6AO4TsKOURpy2zcE1gbRPv2gE5zWH3ScR0GYQhbfR4
iuEeSA7L+CUXEn7m6uQjxEi3apNIgLc96ChWH4tJbdJi2zpuYRay92Op8KAB66g9yf7sMGgOHQNy
I4tVbQEy0bOVkOxd1tSYpnjbupBZaMWdXpnq7Sce019Gz/JSYUY9MuaUFnnxFdYWO4JlF830F4vb
lvhesjZ1ACkANxLS7idGhZvV8gthDgGvAtNnza8YeODcrNihNiKkfd3L+SKlJ7tHvt5EuyP931Wc
/3Y8qoo+oNEeNh+zmyNcJWHfyPmXtfuiECXAgrGMHPppOAdCHoLbklq1dZ7j8I3HtBXUGR/HehGW
lSDQzHYpW8Ju0xYnoGDGdnV+WjPUSuDzujot5l6U/CENqET9JorBTWNxfqsiHGVj8giguuosVyv0
H5WZH2CCmEPO8AR8rpLxDrqt6/ktgQ/UO1ryGak5UuOysNZaroPbyC9Kb/D3ysodd5hNEc5TpjmF
Jao/gE0oNNJa3JNSml92/o/jYzXfW3xlNdXU6EmxjJ14R+LuqJ+GoiUP45GzRrU6YlIHY/KQ4XG1
63E2AlauPy1PkWN2v9MhlYZzAuMqxzUVE3mNSO8m1a92VbjKZpDz7teApBrjX0r1Wq8VaV8cMGWb
MhO2ahc+Ug8Ulgunjls10Z68me8/qLm51XI9UnPEMRS8oIGxQoT64LHlqGoX5pw6KTpbaMKHNH6Q
nQqmQoSSoCF/NyaWVQ/t4wpFNa99J5Yj+0a6UGPQjFL2yWQaoMGo/ZXoYXpHKf0d3YDiRAL2pYWe
wy0QfCjegeltVEv2JnIhnhTG1NHqnmwITY0wqzhW3GPyKnSQ27lN+eA94XkHXdss2/gykyMed5i2
6i5NfHQ3iXdlWJIaLTKJxaTO2TYStIzVMQ2tJ76RCQ4BHd5tXtBkwlQgVVvPv73dwYbfuFN86C1m
1Qe3FatLqADziZUNUYN71CjNYvtW7YIfyqTCrpeDyiVuVYrXgTamaCJJNBd5vYsi3E9AZlIvT+5C
VZnz0uhJlfICMklbRLR3y3cMpHAkRgoFo/FvOxGx15A1nhsglqY2lDaGoKIOaEgf+k60GHoP2SoF
cpHRPR5aQItOo3s/Fec0mkmrSFhsqFKkrcp3KAqLaMA2vTy5Ip14cKMQ+FKDGK6Pfy+h/IvAZ8pB
rIw5EmQcgtz7bI04cgaGZsIQJQp3S91sU9It6NJV8gfutJ2ihj7oqdvVDQvDOEBQOiFej15YfBdl
IAo+e1ahpFceMsBo2p2nykZj9GAqrsBC4V+hDODE2o+UNzO3I5laAvzYemjZmr1/oxTl0ovVt/uN
8YUPkfIeI/aki1I2u/DMqpeJgHArWaOlHmdHneWiqYjhAZnYvlcynXKCUYef43VhD31kTpIx05Ot
ftjN0yZzpvIOJ+Mcn9VbayRQSwPhvsqd0amU91MKw7c40axVQo+NRWpirv7TQuafO18ZaqqN70pX
ZWo1CAbW3/GnWwyybeHnOCdIxQ1VjmxgyQmLwfI8T8ElkMvATo54lpLwTOEIdvSwjLQcYwq8oy5z
xl7JqNVDlzaRG9pIP3YZZxlPAYCVy4QmKT+8o1CvK6qktA/NjQMIy3jmjt0L1CIJ6EK6kKyYp+NI
9ROgrSWjq7HdojW98PA+XzODHMDdrE/+uMm1L3FQcJaPBpT3jlJwp21bZ494GlDwTXWm+93bAgpN
MkmT81UZ/3kEG+2NUDLhlpS6wM8ZNlbQASvS2NwQxJPaJGRNdSRCYzBml1NKuVOpc0C8+ctPjOdL
erxwxncNsP5EG2PYNftlLjZ5Fd4P1TY6SvWXq7iqOsx9lFfQ/lEfGChqzGatrAhkebtqKu/qXmjM
4YYkXsSaPKWlMd3uScPCnTofxtRUU3FBkZBGgg+Zd5ZQJ66p/J7qluqCX8wJy8pagX2tumYbxcIE
ybqzm0xB9/UnJ/jHj105E32snM1NAx/RLE7GnNMrP4i4isp4KZFdV5qDhv1dC3EKcdhWTsWmoAZI
OG2FUaREEYYV6h3XneMOSl4lODmu1YzHZ0lhoB+QecioP1ekdrt0qYtEcb6uIbokT5aGu5W1Kb0V
FyXGTJkAcstOGfT7ti8xBgOisB/rlBGNdAv4KBtArqvuAveSgV7ntWb1k5Bn3Y+ZX0N7ajXdPdrm
qMY6l/gW+BYF3Gm4+cvFY+Vprg51rOYA3x2MbkUwz6lCAiX/FVvg+cerMxfjxlLzwOLze9SWienP
Mdx9c3UbROXZwX4dfV32vxRU1hxLAtEbhVrBBsSZUrNzb/e+C9KpjNPLu1b2gTGoyIW9SfD/7Kap
YVLu4N6jl6HYO2H3bmMv7qeTyVZX7FiwL9XBHDE0DDTnBkP0yGeCFb/BVD+NTPr3bpzLc+9w6UBw
9rjQlPz6+2X9EO7k4giGmnsJNa94UXymEb02rU6HkhC19XA1sp3Uo7Pm5U7tIbMq9j800KWhZkBz
k7pZBvnDTmZ907kGzs2q/BdMEMU+dFtYQI/3/jCeJTDoPkExHbnKd3fUIm+BxSWuJcsXJyojj6iu
3uWdPxfKUxMVa+ctIAWzmvUui9ZUD6iDFcrHVWD/VE2wTSAF/Salo648Ul/12XbqVGT5B8iHjzj5
Y/PzkpVjKZGGPwfUF3cU3XWLEMKBMrRrMLK+GaQm/Xcgd22S5BLVI/YIwUQyN6/HcNXA764EpJb4
fGrT4aGVfgqQZRyoYWtzhJuPaRVEGCp/h7HWRv16Z2EPjD5h2vzmFLSHRfAEWP6PfqIAqrDr+lvT
hSC8CKfn4HHFkjwNf8QkQ6j0C2i3Zm3R2cAdxRJNCSc+hynTcepGJRHsqTPQ/rT9zGzNZZB8EuU4
KiihScO2o/NkP7WprOBc0VOr0QMhrEssxU8HgxjvvLgYg2p43mOqxX0zcggkF7gFkAbZL8U77tt3
iYGeG+Pe244p9UABk0H8r8gnWv8mLAxuRrZigEBdDpfKqfrJ6QAZq5lH5j3pe8Js/c+PUTRe4hUy
wWUUFeuvaUAUjMM1g4Ca83/isbodMGd4W1IjacgcP3//sq2or2XaeJEwxpOudAGSwCDqTUWAOQ3x
7v6g5UU33KIMuJP614mBb/1LP4q7QAsoas+JjB9ulKD/gWHv/pYD4MILRM7UQvVRNEHfopIku1b3
zdPM7GdRpz6y/rBtu1PX4P6HxeJWJuiq7xLDzMevRKuztZRM4DhzaSXnpkFwW3IfcG9eUs6u9ku8
HC4AIiUAl1LjWAF97FCxy8p/ft6wzhFbakn7tWFm+sNgGDK8pQK05rmvE9o/JqFWuxUQ+ORiKaSk
+o5f92FcnhM3Bx60tSefjuMH1IK2qjzyhjfsOwp/+CEs6S7qpCAWETqyOKmk6O3Jw3csWGozrrEd
hygnf6kbvmbvzwQX1ZQ3fAbMkoU0duxsek17VGgQzQ4h7le6aV8fX8TpWWz9YZkwbv9VElm2B0n0
LGnS2AKPS6liG9YGn3PoYSN2l0jUG3waUjo2eqRGlSiWLWSJa7qafx2piOxgIfMQg0sm/f8DZXhp
DapiM1NMkRxBNB0OukOORYoIEBlDnZmuapBaJslsDfEXmvRSYim6UqIAyGLs0QITxtUR2+Z99/Yv
NnPFgye+XKhkew9f5PHXCG8gNqKXJmzo4z/aUOwuX+iV3KtXFByZsl7aGaHsdes/4jagnSlxnucI
fTGBzZixnAplhOt5pFWYvQerhaXfqZNrWfiPPmj1aUKgAmz9EiNNJ/53H+UWO71hQlqleRnYoZaO
4QGxKjyo8CrS4ZiObR1LkOAe1ucaNIQXLkWzBHi538pwD1OBIbnyRRGWED8NcP9bYUbbJtGzxpmH
gXLohRrbDI5yXWZ4n3XfoDoP91m6YwCD2a2aFGsVHvd7/s5mbmo2/rFcpgixMjmuoLYam1h5Xhsv
KZVA2v8E5XgyinjzYbgLpLZdY+v0R0WA7Y5QGFYPLmYtdYqDosHEokq/mOKXmWT7kdtgP4mVFdxU
m4uN7+2sci8aqWK1ZeAzMS+QuhbkF6PzQKv+6pnYyNYxnWMQNXOG3Z5mZI9anUvDVqOdqNx55r4W
6Q6KpUC2vQ8D2OogpYnL1V5S3F3jlRq1htvffVpXC8qE1cp0v1C6ZEezJSIBMX1IT3LJ5u4L4OWB
WxjIysRU+rONe79ReoDhGrsbUE+1GqHstufjy3TuifLi8lzG92ZFUFxLv50cj+3VziPt8CSjnXij
JEIUGC9ABfNIS5qXR81nISfc+hGrHU2MgVJd/nytAdkWpZBWahc29f/+lCbfL8uDMpywVaxhsmok
PRlSieVd3R1CdkHXJHumFI94PtG0py8dw+rRHKXx2Y1vuflbd9y1g5APUuD+BWfSkCgp1MbcOHd6
8gPtNsekVh0DDr1pQPHEnqGg4PGjmam/+0p70hruuY3zk3fKLvA4eTflj9EEjbnBAQET+c399jS8
r7a9fYPcE+WzlfrfXyQgs92Amh/yPMn5sKIK0n68n7fNVR6/rpm/RxiiwK5CDAL3EEVydXrNa5Ak
h9URPSBO22mKB1ctMfMkHjScGk77XIzo0CjEbem+uq5R6lMMZhPAAZ42n6ORjmec2GTJvKaBZA6f
B2SkQNWMH8J0EH2+dIBVfoIv+h0aFwg7s489trecNLdZvR3vl2DrDmAPaXXHfJ3sFMeUbeM70QgY
baUQ4vqntHii4UOy6hKxPb+oteapMLjvYOhwlINXrPwF68UYeWXfdxsKK580JsLhFNpvBcaLSgxH
hnkwHHHLQVNFcHrWKdiJzQjNsst95vv+xjwTIT698wKyi1pjr9/iDFDsUrsxZcXTI3KTLYdWFzAF
ySNczUM/28rqSFySvPPaepHY3ifNzc1PLBo7j8PMm2RH/flW7ObD+rfiF1hA4GQWdz9dnimUNnJ9
ASDSJSod/u9htZU60x3R5c0Bzt+DkNO5SvkFzj0lp9D8X8YrL+qAokWZKJkoAreym7susQa3E9ED
bxbLXNxEDZGIfFw7kTAh+7FgzJ+eSiDHDgM1qTo9p5AXyfA+3KErKYegLI+i2W0wxXQ7pmRGnh7g
TgF5UTpOlh64ZENBYvYuL6K7zRCjLCZKYY3P4NmU5RthcU7R2kDzt/BZJVjc4JQM/L+hZO70JDBq
BsuTqniiPBfWrRBX/f6epuOHxTIpLnztFUqiWcRqLtauQEXeHFR3CtU2Ddr3lqBLOLZ0AONdbyYJ
/WP/SI6h1o5ehlbTtZ78XwCXBwN6djoiw9/WxkhagstJ+5VUtI5yufHvoDj7cgfsG9mqy8F/C7eu
cfPmsv7HlxGcSMRSFfpyIdv1oVrJ5niKgGNSnLjrWF7xpafm+c1vcChsKjdAy+S3DaCmvL85c10k
VNkdKHzzoVW3Pdg8eomyYpWc/pC57nLhdiOiNUcHw65niE/XFQkX0cww5A8iRmzLR1FFwwctkkyZ
qXzoey16rT2MtdstG2BHsNEhVK0nmE9iS756SPc/bEp6Mt00OGW22nvsoL1Q6dM+P3QkBIzgFJnI
WINXu+KxwI8ZQvkaz4vE/Yc2/aKVFZXM1It30o+LESRqs5hdirKJAQlXeLFu3mWvq3f/DyIL1o+t
H9NjmApwxp9V4IY0L/Rl8PCb8uMdeb7enpBB2UhjUi+QMmmXnBRpjx9BB6kFXSJlR2D8wZlYjpyU
EWH4FwCPbCqHf3qVOrm9IwAQvpEZ9ujpxOATrOmYuf5v2r4eF1giD6YRy4m+n5WPCJFMYKqMukWO
Enl242qZ8pGwUbPVaUDy6jXrrRA/e8e0AD3jvDGMpaurPNRWrCk9sA0e57Yr69l4pl3bhJY3I7jG
JDg1n/vndkK0h4d/RHWLO78G0/0K+NGpqoESLljZZoBumdw/rUCsJOpZwohcuIaBfdEBO86GT4hj
QF7K22KCKXYIWM0F2pc3XOPioX0GLmTOuwY1rkJ/fXJWIMl85JoFqruaoscriZOwEg9NFfTAPGZ8
sBH2heRdYi6jgxuYwl4Zg0Ao4FrYB5Rth0+MD67eAr/GOnS7U5nBMBL7TCDWLWmnKQQYGOsILZNW
P1nGu7hHN8UogX6PmLHxvNGRcSjKbv1IiOCO5L3R1Mgjq+HxtMAw1uoxZe8Gzz0TiVaaobkINO+m
1gq0R39QUPCzFmIItwwltNmmj9kKN7wm7g3xfaIpF02lf7I9110xSMs/0cMA53lweXhmwad1Jwef
WCzU840SOI0sq+C8signvz5djb1MFGD/d3YJnqFNe+oNqR5fer+GCCyCbWDVUAcADWeoQqsBtDxi
JOHGGuvEijjRg7qPM5BTmxjYdrhFJyjk9NiWh3MQI7EA+1FvGkOp+BZcWWZxi8ybPn5OwcKsTRxA
yqxf1m6aZtDbuYl22ZCZL6nT3PcyYS7PxObkVCcCGXktQ/4qgkYcYdjPY5xk8BY1Z7veZ6ic3TlP
LopF5ilB24j0JFEsrUU8KdfIwiJUr/BZ/k3T2bCTEeZs4D6fJIW18jFsaKaHjKkVdhcbXJOZ/axb
lPgMEyKUH+5gtYf/QF1d9apxR5DtL8jIHtuKCiwu8BhdQNsxRSX2pwugKt8AvvfH37JgfF5rD22V
53UMjhjL6igdabH9K0xp1cBUqX8Ya6AskNiW1Rp+jjmEUJ3MnxVbHDwBnfkuJ0Prh4sdFhDXoBh+
XlUYaq7QZ8gSd92HGKpxOJMHXTsv8c6LVCm0u/mxmIRMRivamiLoOfKT5pB0Ng1kjvmr3yK4NH90
k4zICFHgWNbO3lAMr48WiJGO0umAKyyAg2+IurQywGFSfNmJKqwglPCyoiYRNfzYi/7lZQbfyL9/
fvZboiNzrCYVcAw47Zg+UBbCdB/Vg0ZunVdGQ65t/znMeySGrx6kGrizhZsE/fZlgZYJKO7qDblY
KmBNzgMYE9KTdIl+m8K7jSH+pIuCqN6SaFeLZXtbxjm5noMpXfzcu1eYeTIV+GpuLO0y3Z/51jwn
I1Eypu/b8qKKOEIN+U7wxL0gp4b5OK2D2k/CVydX78TMHQFV6EByNgm+MZzJL8tF6VffO7omcE5t
Gfh0vPDKboF3dpPmE9iLKRD6NFrFCYsvh4z0Fn4A7bgKLBwWYlAbKK68toKp9NpL3CpNFIgIQseh
uxIgyFVTStQstvBGML76laHBj+GeO2M6FurNhAluoV+kJ0LyEoUO3It8Ry1e/3JcTO4mBXANCN/b
X9WdIJHAvwrALzS/7JZVyFMs0xHMSm7eOR4ZKUaEDU0LsIc+wVCQWhfHf1m/6GItSa45ncPV3NoG
Js+1ljAt7m290Txe6Mexp0rsvQ7NEsNlMhHsWkzoX9aZHHO5lp6aCy0J0Q9LlH9ilsblCLyCd70z
SRR+8cuNR1PEM5Kvg8wyZHrsjRSANW1ePx5YJDCa8pBUnxEE56n12wsKEAD2R28iaklIrrlqMNVZ
QyFPsAMz8qqMS0zcrm6YwfZ+slbmDbO07xX+xik38jDEFbIcBT5TV9LVypaVxWad9o5ho4Z9U+bU
Xk0jr48phbhOIsZbDO/vYA2obxnpaUYeubodq/lfSuPOWx9O2zL0cUenPMUyhA1WpgJ8zsYT92lo
V0u3AToINqsgT+nwtYA1QVC76M8XGywmzYCVJahu9OtF3FVP6z7QzeeL3/+hLrhGTjQqR6Fpnlt5
S4L1Jjq0yHOojic607n8tJb/4EDWmdbHGk6ZCis/UwSMaRqamD8c4QsVr298nzQm4xJbqm/aaerB
D+GWExmUFksXFlnTzc0tJJG/hif5x6YI9gsXI9ndA2rl2GwiUbLKrHcsnKT4snwJiUXvDJDLCm0/
4Ggs/mvEfO0HLq4GJ4Zch+w/24topUpkr4B+SQdSDpPnp/VWWk1UWrauoz37m6vsBlux83QIxR4K
XoaCU/AGSq1bC6xVMkkKUf1T0zIRm/K9OfTgWQe2HQajUkQb75B/mME6G+vKfxFOV4s2cyFp0h6X
dhIxHzyJxd+NrsPrXDnLTxj5Pe3jS1t4A8SW3eQpV0Lpe+FoshWBMUPrR2NdhvvudzZsEo8ERpYc
MkSK3agwojgqgu7xMM/drd/Y6COt4JwAccrX/U2y0qADdDIaCCsrhpcYRoF652WM2QjtC0hL0era
tDyvmEpcgW/ESEOJka9a6mujOjFXgfuBfXa2+5fpozlWQE9TDdhMAxfIlvI1MfxR8XH2ZH8MgjNG
k/BwkXncdutVHQ9PEwaVeAwDOIU3edIniuduB8bdQyxs7SMMgl81IFB9NyqR45FZAKY/zbNg49MD
133hOLP37YAlFDW4bdUP4wWz5jM65P+uIL/GF2NYysQvUaU8Q3Zq8dqWLN/0tqYEZJCsqGUn9BeB
0vj6lv4IM8S43p2rxD1YB/YXqVnCYTutuVhHs8nEhiGaSn5kUuOTqw6qkSMCIt4z/FvJA7oyLN+n
oRpbxY8QCkXZ/uVO0NyhaiYS4ukm7DGBC5c1dRrBlj8UWDzsk7o7Q+bjfTAdQl5OG157NEUWE0mF
aGLgDHaB81oDNe6vclpz9qbPzxNXdgA+94hL+YxXnzE1Arelgk82s6gWOduKE28sOH2LhT2NEI//
AMghxXZjgvGr2lAEJ01yskSc4RwYdFIptngN8yypXzq9uQZRJZO78ihB6OTSW2G7B2gUGKJvW038
xOopZXRJOGGRNgYF0d6balqk8ZIrxtY6DKRLzKk5urlSo74fV9IbAMpCgba158UX7h4YyFphbGJl
vQnPwSBaLIWoYgt1rSZChKcV+Z7blTz0+4/+AEvvK1u88TOk4FdVkp2VYJwwmZfkqtaYcYZIx2v3
UNnfHY/MiSyOOGoP/gSpcoGrWIKoKtSmua3CeWnGW2rb+QSOPoBnA60qU/n9iVvSE9Wl8vasCgqt
3teJhXD6kx9qR7d0002OkEkpD3ziptgXyLS/1wc2t8+aUvg9uCIypW972J6kUZ+JSx+KGwIvqywJ
krZIK0WIf+cVI4m5OpCm/6m09oRh2z9NckZDHKoxzm7rnVrh1wU54GFIUwujpN6lz2CD9/aZP24I
0B/tNnVnsTm5HpOVmd+el7VWxBFMfrJ9oCLWrRw1gTS8kGOREuCj/hKIf6YHctk1JaIJS8nGgOxO
MmiKZkvhAjCsnXTeYJjfOMbrAHnguPkotOHlVfhtmSRPbSP/LnzK4E4rlrkoisJaGjRzDAVPN4Xf
GwN9sEnG17m1+Ey1MS1CLnYKjOVBCf5h6Yv4BxWXD83MaFcD4KzhRAwVnAcopfkzNE/+6hwu40M7
do85D2aPXpTGOpXy+xrgQzxLxnZEnYvVBflwTZrB7zM7rMYGk6fAE2AhSeDNTVjhzJpriTAoro03
v+aNa+iTo0mThcLLN+NH+nA58XPYBvbaUlV5MyFOr6YgCSlGes8q3pDa2aW2Wd1a0nQwl6FFAipY
tklW3QrMnJJtwsGqKPV2TnBE//0XrAb2x/D53vzAiGnUCMOpXT11uOLsXmKPT7Z/+TuRfBnpy8Cq
+72bSc4kD1EuNhB2NClIKgOzFICM6fAxr/F6azpQFIL67Vl/9ht5k5jGaeCccN1PYQGWGiE/Pr2W
wzr3o+0ulRkcNr94eqhsMPWJh9oxf+JSiUAQ83P3CSLf845vg8zWsutesUiMttcyQrf2YnYZVTqY
7ATLy9w0e2s+cWXZtNYHM1Hw0JOehD286jUzul1g+XeMAEMHMBa2H8Ty0Whi64Cn1A0WI9gMpEwc
B3deqcv44yRVusS8D0YOcU+Yu4Zj5bypdRH3JBQdkAUeYl8Lxl+Ieuq5XFvH98MMNutlxE4xV8rD
6ep1QwBm4t482YXFjcMvy26ukD+piwiLuGKZ6EgwedGaXrUJAxbRJiDKYWOwSJwm5O7/0LQhFHGb
a1Bsj9uDzz3Mi5np8bMp/8w99oKUO+rhiS0J0vt8kde1yCeGC6VKpzaSJUwO7gF1Xv29yFrB42E3
lA3l6mLnSmVtAbS4l1UbRKQYkdaxTunHtGZoN/NXLETpNlUWFdib0d/bHuBkiOOJxHGZZnqtBw4l
AHwma18rrdIbczMxYb+7M8yxeAc+z2uJbjEOVKpIXL6X77M38RQYtIU3tezwBpo2PQOTDnTFIMUb
0OMlBDbVzGIW4htXAKEZZddxB2M2HXZ/I5VTub9adCHjo3jFs9tdVkV9IvQcHOrmMH1PfRBKErbF
/8MYRk9VCCzSTQEfCaPPQTOgPOEg7ry76F3nvGg9Vzrol8bIONDet+hdejhC+bV0PxwAgwHKc9vD
NZ82117Vt+2WtbEL4nkJLRo9npEoHq0CUQJLdLtvhi0kC8hqJsYYdsq8A9J2X7HfM1ioGziwhFVP
LNhDWegE4+m7LySL2XjVlTMmaN26LOf3c02eU4t0zMxCqAUWiFtAdWaxlj4yugQQ7lGEY3w6lZvC
obosHTnwlTZcVmJ/4wUI8twyqpWs1RKOsfMd9lsxVpo4qyiVA/62EY7mT+jNXuP3TfEXlVulvIyi
fU2J5xTJgzIXGf8YtYUiThIhAJeOn95E1vFVvklyOiU/tP4gdeHvSXXEyMtpIVjAut1bmz4JEUr5
tMCG7o5byq7GeBy6uqX5uAZZPgxzFQY0CqHda4NJiVyM0YDoWm4moH8MZGq1rfNiihd+soTv7CFa
AYyoTH+I5QpBW6wfPwHnNBEA+DmGQheec33thEvIwJg7/T05e9LrJSFZHz/QmS7VBcrGuJCq/CIb
VuEeVn2is1ZPskk2Auv3gnIKW4I0r+PcUYxCU0gyt5IXoHICApgDp2FPyuDyoWItwphTT9HdYZ/y
MZMj/SG91PR3P4iL29AChVtv5P477ucWsGrrwdfIiq2JO66eQT9Kcm6dVujSJODQC9YB8wzrg0bP
34gmG8F5QrFsAF47WfePrQpyNkvATyjgPkLPPRa8FbYIsQavTgBinReeafWLMRjFlHXuADVWicM1
5kqze8E9uCNKN5trlhLbZxehXiitReLctd9hpziP3BYL+OdzJAUqmc19klDCV/kz/DKthQBEFKhs
8Ge+B/GIqZy4fdEAu5FLJ3jAybGGFtwi5cSQsxrxNVYZBcAZYeqviEvOx9UohcGFx4yEIpH2fv/Q
JFXJMp6o4LfQTHo8FQz73byoP5FZX+LQS3zf26zPRugWx1Bhq/wCbims6qmAS4UcPe5tr4cQzfS9
06GCKmhXXuQE8GDkhn1Xkl26bnRiBrRp7TIS6oDcvwekVTxChMyHkUJ6+sKAfKVKTCJtsESOYAac
+UiFtOoA1f3J12k9R3Q88IBu+lbFPpG6Hw5pzS0z/UHNLIZZ/BMMDJXD+7IeQarXBUKCUA9ZhPN5
55y41sHk36oK7KtSIihhmCrP+M47y+UieGOBClVaYLqKM7Sh0NshuFzMwjaAwAc+w/aoBsg47TO5
Ya5ul/IfezNPB1N2hOHlIUcVopwWiJXzN4bz39F2Z2khJoDQHaFUVUUcWiK3noSrrg+HtZP5KKvG
uzsWDA3WRaeGTGJa1q2X9EvaGZ3AIU9E96mTIv9NcMmphJmgYxucvqFT39kGXHhw7R7OQJre6ql+
G2O7AhB5/WGvtJk+/yPQ3QPdYFS+Hc6WiORALj7xECaPk8wwlOfX/UxeWtvfpT5yIa/O/GuKGr3Y
yVcpB9J7b7JhAcZaK9lYTGHVc94ZdfH3zaZCStlM897lq3DJ+eflzo0zmy4lmAt2V95mcaGGYnrt
YIUasFAupD+mkUXmZTigH7+yl+7NVuPrGLHIoG73lJLW0DJ6F3Y8YrDF9gOX0tphr10nhj0LR6ER
aassv3zg/MLU+BRmqGJbvXiuPGG0NSESMbqOtGvSXpFtjXnkf1HhbGmI5yGRIX6J4MxegzP1rAxw
sxa86NuVC8FR6mccsc7hTzdrZqxilvYIEHVwIfcKgs3m9wGE7xZgRHMUyzmyFw7z8NFAy+yez74B
v5iuUdzfRQEoPcOt64NyhdNYAnh6NshCmZn2DNGcAJ62PloqvqlwVJj4gFUqEztTQiWJSWAdmhRI
exeugSzAxBD0/YNKNv23rfDwfoBgOKViep1xBOBmSX/U1U1657/DGpz+X6ClB3BU+2HHFYXJ0LeI
gQT/+cX5vA8eOp4JKtoHypugqG+R0R41FtZkXzKoq+MzpBiQDrhfMLNwy5/Ag9+Lfl5NbFABMRQH
koSS+k9kRfglMt3Kmg+LwN2AxYGKfDhm+zXb6AA9cvhWD5Dg9/lGgQvIBJzSgjk4nRz3Ndcch1Lb
+sU32tDzS1EcAa1UE8uf/e0DKLaNopqxAdhCPCCLndoJV0ALNMfwgKaYmWBWfeBqONVAS3y/GpNd
5FyGnIyv8Fp7u2sX2w2r4sucdXKmn9F9b4/7QNSKjkq5qB9DziqWtP0m2FQ1GeqmYp2vBbDvtMfG
X5N26FB+DnGVAxZnfBkjIu/tnaqss4DbAecv5wbzHhdXpNcpprP2L8DS39fgYH6Sw318mpdtd8gV
RUdly13Qluaxiuy0i8AVAk59Ea74FjnOtceA6AnsvQHiaJA948wlmGgPYkM+RN6rTxxKYHufjM3A
JHex6SyZ3HfxpGguJJHeXhnTOpnifMz6uG+5bwQb9brfjvqM1beF0FKJr1rwE3+8TCB4mHe7I3Ib
NCt1iNpHW30cNYvH9GQhv0QfkS+6xhV2UR9YcT5GlV1FPDwCrCRPZ7mnfX12jUB0u4rKpPfH5pCD
MkU0azMB5Tx063GsPM8xocKyNdRAzrF4je8pjpm/h1MibRzTNOImkf8WcmLw/iaTJIBOHnz/21/E
D4Em+7PuJixHAW4HR8KKyedVwHTarJszGjU6PA1UYo5o+Nyn9PfKPZm/LGIhK1OzBXjCuc/FmiXp
1gNOrlv6NIm6Yo4PR2H+Sb+1Fzek8PggfuBjIIwV9U5+pugjWYLAkWRQqUuWS0VczXljdRuqla3s
ZnynFo9+BWOnEUoVIFnLuXQQVKHVAgeKEJl/PjpnQvBLiPa0oEt6dvDvZADbrYpsUj0Fx172J880
AMXP9LXd+MdV2wNjrqYX6Da59L+MWRRzoFpiVhf2ecvRY7E4dbA4Vso3hqKLGSnLo6yjmpfzS6PJ
tGbHmPJLIRmC74NJDsdT+f12eeMkVJvdg1cX211dM/o8Fp+wa+s6N/JYeOITP7guQyUhQnlx41jF
7JLZFtEq4rMdYE+TtW1HGKeXqKbR7l+NFT/kB8mpPyD6Ism45Ksbcp1KusC4YKyv/RevVab9ujL2
0C1Nujm4NuyR0SqTVDx9l0CUcy65XyrLs4WRo0OSaqrbzee7E0fq2tbJtd4InWIjkPkmdKfn/TmF
24PkUzJZ5x/1IAq5BITnVnKQN8t8hXbV876mtRubjE16SgRDBf1q5FmOJHqKfeDmc3kn18nNl/NR
4/7UdbmVgX7oq8HkVogiBvx4H/5zYZ9fc2Vpm88kSziI8VPz/FLP22Zax65vbDdt6A1kdWWFmh4K
PsL6x5saWJ3waGyDqTDINevMsv5enLRzwcu1FgJ5oXeTKKUIfZhZxVUcd4Akx8nz5jBYyVRWJ5Is
0++n4GL7VBOgdgrvkQSTmEp625dALbmk9MS/5BlScncHYtrU/p1xzwiqxVYjsE2t+bo9nax1SwbG
Tm9pEo/ilZemLX3IKd9x+Kn6zD0mBDFWLdqNsSSprwniEzvBu4Bd4nUSK1Fd/CcixOpnDEvwRdM8
tnPzvFj6Z7iR3Q1qJTVHATMIT7SWX4S4hDivanS+dj+z0N69Fwrl69tLQvU0asNoeLZNwh9g0AGe
6uHepn9if2O4izFvOYaZDWyRXO1XFdXVWqemqz74yIl/XYnvkK0D85mX+hdPU3Q+m8epJfjqYKE3
xJTcostKL3akiiJwIDQQD3fNP2F9oH+M2Dj6mAWsL/5PlcAhoqQSL9XOcYrsJZti3qR8cx+qijTF
CIxsZyYA/C6Xm1hcioWZpDf9RKjxaefw8fMuhXKWnZQ5WmrZBbh4EmAn3EWHPhtm6OPuaJE50XWF
2jfiWNIf6RN6pWtA3OoQBI7Q5IfHgsM5KzdFI11RGXADAjlQ6cTceIyfsxjxkDZ2MjueQiSvNuzP
pwG3LCgzyeiI60U2NCZIc+0gnnARFZPkbeUTpg7F7+Np2RyFaRc78KghKfIfG52MBU36SHj6hehz
+ofshAkrbEkTi8gsoQqWxDEm17UlYT15Q3BklCQvpFP7bA5pSHsTZHeYdOBOVgMV5bfas98GAK03
AhdOX0iWJkxPHlL7siS0O13QEu1+b+Jmh8CS7q1VcfIStzg6zBUY2nfvR8XhWmnCHjdPFIBly6jL
P/5cdO8h1tsxA6UMt8e7iUo9ubKvBrNouKdKhHmWrJf2vM9P59X/jROqp3g5phME4JYnYNBmBIeC
Ms1MHwnYvEeli3kIcpbLf1I34KCAxdNXw6cHVC557pGKmT/uRQipRgL9kRrsT0muRecMCsJZ8gEp
ovKrV3x4T8mTgzKpAjBpvJAHc99mpuhoKKxHJ/WlaPrOj5t4UwXLQh4DCXGT8SkTr8AMzpdLfW3n
mvlNSEudXo25xXiHeC1erj8yjGXeAwNFz5xtF4egcvZodhKYm2ZB4UPaL5LqWnLwLec+wdSKdcbg
s9UTF6pgzo96Pkz46MtD8UNUjVwhaC34h+cgJgY0MFhslbQKoeTVI6sdjvYu2Q5M9JJxjG+tjZyu
ZdusmmUy48l+LG1a3rH7DeTDutFZMtr3J2pycDalZUCja35T7sRaqvRvsodnbXXoedbu6YYw46vh
JKQHUrBo8pJWTQepoHHiSoTHiKuF364jo49WzPZMiEybIiDKLKKNsLeAlEzFo+xLamAcNPr3Bk5n
uF/NYqJ6xfyVv/EM/ZUqB25J1l9RDl0F1c8MQa57Ebvihy/bf5de3VmHbMgmS4v5PSXIKvlu0ATc
bL8SmT/PxQdTFehSmYELpwmUslWZoFtLmNDth85L0H05bpifebKRkmHIo10n1lRlNXPSLorCGelT
4wbclN2adf1y4Oq/fIszI0gYpSkMjY0SKoMSmLmmI32W+ONnSlv5GNdldCNP4BLuG1O66ToIXOpd
iHEpkc/spLLzgFL4gSvsMDE+2obzjiHHu+hX4TeMRRGIZNf3++jwIENd0mpmpoFitAoMskoPrw6N
RE19BZtufayYzHxg5qn6vci3KaKLtaNn47jECrIkFiPWdIEevPIgOOXeTrM5u3zfymf4hhxSejJv
mLbXODTgXxsboInz+nvTvcpZcOiN6OCpPiSu4l8SeCxjTgB4pm2ARqYI1M7U9ZNdl6ABxiXnbQe+
hoM4jjSmAi2j4fNsDrnLurDT468wRS7qvHVovFsbawjqD7qpC/+gu/gBv7GTJIAg+yhv9t/EgshJ
C7N29OXrbgBR4W7jGMV6fZQtwHhwOaZIY3DOh2WspCjqxC7d3X7NsSBhXwe76EIX557Gtdc3Kbq0
8c19W5bafWrsqmpA2Oc/RIJQy0o7Q7nTe8MZYyKkEbFDRbzMCCJHropoz8LSJOd2//s6iYJw1GyU
zt7g2EmMW0i7dSCB3svGWsB2nU4eaPEOwGGPiDjDiKjDKcxgGGNop8Z0yZQvNjxTQ4HtKR2nsikT
z7Q8vDPz8oGFyjZ8MTsYEw22XkqjitEv2W9NF6AK1JJ5jbwTjroAuxtJER6CP5bcKaQYJe2lAzme
yXc61h9JkUSe13KrmcD9IjSpAKx3oD6ZM/Oo9ql911qLRcJ804d/zso3CtleeH/SJBPxRD9VXM+P
d2ScsdrSxs1eMDPXqNNsSfO2XdDvj/mdEW4EfTohx2aFR+0dfT6LxSwlRr2LzyqRbNtdwRjaLCnl
pI57qrUzXiMHmzpFPu7NJrtWksUyJ6r77sYSQv+K68C3FBHB/ci062nL8scXXi5Iy6HJ4eDPJ/KC
7GcNzgJpmSLIzpJd2XNK0weQs90L5DMgZKWQUVBaJbCVggxqMG5GwAov0l2gzZi9LljaR+fwiHdq
H2DI9vrzTFDL+/4MXJua8hpF+PTqOISuaUE334tZBbjZp+C5XOJFIIayL8kVe7AJJh6HMRWuxR1s
1tNgNpnjdk6xRohHo18Hc+W6BXH+DnbE0EaEJhTahl6mu7HVS98l1G4F8SkQSZthcs7vYl26yOPX
Y0niuoOL8yjotoH+p2QhascV0WkK8RWSvkWc/yaZazEI61eB+zkmTHhcz9abEZCIx7kPTOdLUBb2
fKVjiZWF91tLsOzMGUtv3EQAfmoxOpTm+FfHRPQ3wrdexiRdp+LUi8qpSlQ+h3rQKqd9VkBVHAAK
+lVhmuT6LytGkQsir0cyDPn+1m32V4bx9Yw85PWRPJ8NfpBgOXdl1jiz1SdDnnhEICS+6U+x3Blw
LzRThqfH2lb4Zt/JjSX9Ed7srvSDb/yCX+l32Oz4bRpN62K344LyNjwMScTqsGO61f5b2T36mVgJ
mHCkl253EYCElrdwrnfCSSMgHEE6cSlwB5zreTsqU1MOU8aEwkLwqqF0wcMs34eFSMK6Cswutm3M
ExaSaifD5jxOmMtjOmN02DVVPUHwwZuWHkzDG9S3qX/hhGKA9HRVz0duDy46tknYMKSqlIjz/pCa
j9hWMqq6L8NIx0Xa6Pbninmmy2s1LEOfO/ASPyepyoRtr24ENX/fC/9NQy+d5YFYjZ0nKiaZrV7f
NQzOZQCBEP9RV1cjXpcbApJz70O3gp3Ta/OP3hx/qvxRaizH/7Yf607vZ1F9IS1kAH6GKpbjJ7a3
kT69CAVQtB6AzV6eIFX/u1vciRh5LaChmwD1UPt6+787YNx00i9WdqimXwrVA6wQBYgrKszFgwVq
lf+5azzGHi8BkYoLryw53HOVm9/mOt/iKtREbd9LTBOHtPa1md7oATJHjGDCHsQswXxLZX3mMYZK
rbsrk9bIT4c4Ak/Y8aqBk4U5W+z6j55t9BFNN5ajsN40UtjbFSDt+DtFLWrhbuBXSDO1/z9O6LHV
70ejOylxjCFn4XrsNCOnvaMMIy6KkKi6lzuykNoPMu3b0tZmiiQMJEFGF4axNTtp4EeGBL4pxABl
FFkf7GTFhp9TaXTiAvRgUhuM9Ex6SHXf2nEAXC93cCciNzND5maomL+BhDd86ZU0C01dUIi+PWPk
KCkShhuu89i9B+QxMEmyydHVbAbuvl18Rt7Fm7Yp2bnMMW53JXR1rEe4nmdd+V8SxNoYOimYbuDf
jZ4dkljKsw1b4+nbF3/5YWKjvTuY6TsWKdbXgRIK8ZhcA5HbCsL0AOEdc2pk7DCukW/ey42ylMPQ
P5d8FNKUCWvFLFMgwK2lalrRiHzj+v4gFzA900EF64L6cI0mSGhbtdqWHxzpTkC3KPmmAOnutoWZ
/DExmzGTEkcyYN7NPTK9vW6PPKEHpLTAnM6hbEDMLUClAaqMHWG2So0KK8zBvPEDS64JIyMLiS34
eVOpS6ccBu62TiDnblJRZwLOzO0oK7uS+YEnr5KWxASUS/jSrTjZE8Ble2hrbi7z1cVsAxjH4tth
gKcI+SqVGNHOSWU5uanlOhuGCPpWLSiZQ7FduYH4bUs39MS6g+tlpuzOaQN3/r3Cg/7Aj5lhfVjr
O2rbQSf9IyIG3MGSuI2zm7HvlW4NrAHfG5M20oD4uDl3/xZACDi9JCayvuh3U8atwLMO/FfU2TwC
ytKikxRI1ucdXCdaKDHwb7qvsJsfFdn5Ldmiv19avDf++gKEJRhv8zUefcPVQsD4vxalIBV1gRDN
lpu4a60DCVyGd0akH/cmJ796ubJCX8pi7HY6j0+FCuF79NU91HxSsdD4iAUHe1BqI/AH4VM3q0fa
8EBo/EOrLhHuNN2SLcY3lXor2td09wnd9XaSMVB8uNgYpHjWtMk0VZfLWYgSH3AoR4xPTup6eOnM
353caSAeshGUwto58+L72VPnCywHv/jCkn8wNtuw+JryDei9die9N0u3wrpK1727CvCDTmcv3jCR
yhh3/TNrxln0r3JyARhmL0WPsYANQdmgLJEQD88S9/Ce32COXAn7CaNZOX6QZSZC9/Ie5pyCXkWo
5LqbCozthyOYh/MojcoDXP5MMkkD+JQY5Uwf41iwrxvpXWeNmNBI0lSoCuDDyAKCQ5he5qnrxCIP
JAvMRVvDgPKVZWbiGJnLrIubQAvKbpCbkI5WTN8UmOJ8HulQOTZSGnWQSQTVbgJEkpNjMb9k+y3m
vJnIH7Q/KoHNIBJYyjJaR0WPY4vdwsnM+ZdBsPGElUDd0SP3rL1Srh2kl3I+wwn4YuzLX09QY33l
lTv8BcYb9Q9PpMAvcLBhhbQIHI8DCLavqBha9BcUWFx4rguYIf0YMq/10D5frkc4G48WCqJAXIBX
eRf4KBzfrT677oqKIxzndYPNQLtN/YfKPb10BIur2txqOxRkGWbWpvntxPev1GHysQcdacxFLy7q
Nu3F8zQ3R4PAxxZ8VqPLXUSvlLDgnwuHu8ggHbcttpXjw0aM0adUvRSXxWaPS/8wqL6ZS3zG2VA6
JCREjoZfuanvuiGM0zv0yWBVS9gZtubOZE5si8OHUdMX9AVLErGeTGIkNAjqd0F1AuiR6t97Wne+
6itSIC/uVaqyDp8x4AeB8wnfwsLKsvdYSqHX78flPJrDXmhGEPlDCKLxe7FKsvP9ywaWlsnTKTUC
AODvlbyTTACYVNFCZcpNJL+a5D1/EAJFoGvgmgwfQAmHTmRxhx5Y6DzY6QFjXEH07l3spHSywbYu
XN4CQ5lxY3Fo/+n6Iys1ZhMzb0M7MvWi4U2BO0A1bBL/oPcTFM33dQV/qBihL9EjFf9NqOppP0QD
AVVNnRYL+FtajjEOn6H6FrRN9XGSpWM9lWvZVL7qPj1S80uiD9iGdJLILb/29wo+GKtIaHQxupT9
C031FUYnuiFD8Q/BrXm/wjkUmmUM2+O8aVBLse+XkShBpHxlBYKH+juFjUaL+NULwyrI/YTWBpAm
FU+LY5QlvvmMCmfUYH0IWLAViFS8Rz7S2geGSjLRDpLpgkzonVa0fWtGsru5is9fvyEXuSN//AVQ
ngW7kOfcplbV7pi5Hcm9TvC92rcOeNZlYh/OJ9BrvRdkhn5XHW7g7dHyUcZ2Hc9N72DsdluNcVMY
4cqV8m+Hx413SiYNGsD07vwqojQ0aqmuoBalP0LGUNrXFCG1oTR78nWh5mwU9FuWGOjbIwhKtlOL
ieWjtfn5MXD7rxKtMTp2C/CghwkZOLPDV2BHWoKEXU3f0hZmRBAfb1qQyVDRVOJSDXVyrrRNj04j
tkfzU5Njm/bC+CKgbBPLPpOkFol7qgk8uDz0lGP/mG7CojG6JsXibN5EEeQvXVqmgzCzfMRLMyTH
g7dvtJZRjiE6pSuRspjWTFT9f6su9/GzYmrk10QPL3CVYoFGDPCcR8vL4aE7fWHhQj9W7h1X/YLN
fGSaXp+Py+Bfg5FVJP7GhzDuinH+K92yBTiiWKcwFhVFGfvZe4aTlMlzIBndEbigoaerE6lwoIHg
WnpPN9IeK+PVYwcFU6uP1vyBsVNoU7FLo91DL+Gv9+aNuYgkFwX/KtG7C/x1+8qDJ2FVlWqOxymb
di39A6BN/zBPVRCns6Q71mWoaxdflMPxzPXFiwrJsxq6ociNH+fYNyIFaUcPEbJpFMJ58f/4XBJd
+FbmcLPDpekhItiC00b/uMpLFtnD9eMFzfFsYScb+MKt7DMy0WZjT4cBPwaDf9y6AEQWEqQu4cx6
p3peqnH1Y8fSc+0yhAWqrVasCEIU0u9KuL0Q4rERPVKJVXgHmruKZDKMk2lz6z5WhpIG601GgtKm
/rFJotibDvuBw4Z77EAqzCE4n6iKn68XmvRUcrFfNJv7ivP9+MTCT3pLpo17yUnCAyS+efKeOIC0
g11DI1ckt/N2uMQcUwHiSnEPGtW1YUeBGhkg+3LZRvWcNtwKaXKt2nyFctWW0FJq1P9AGxEp+3Ds
iqS9MbTFOxnZ26do0SemPZ2JIHK+7Q6UxWUW2G6Jgj1kpTx1g/5CPXSBNFyUG0IMhZXJmJnQIZxk
Iqc3BC6Q7Ewm5TnWBWr7zWIZA9MCXVCyYZdKZW6fkFrrx82m/tq5yXpPGyxecR711j4i381pQV3/
tHl4RSfDA/S54NUFGZvVnfcZppGKnaeS7yCImnKEdsghkfhbUBKG6CYQFeiVwevgiK6boYJo39q3
UNqANKtrZ95O23WGlc4OYMHX5dVTLabYNG+EQ82z6xgAPSLXvoeaX8RmojZAb9ejgcjhKK4Lsv8/
9XAjOKBugn2/vVXb3X9kX4nv7hr4R42DKfifpA4dOcvh9wssLd85Su6MHTN3QlLl8P0okcYoIKbs
n5qhPGtBTafzBHa/a2xbdC8J+CphLLU66WcGn6kSroMRCbDBVnbtGmS51uTX6mt/Yu59IPpSmHkk
S9OBXZjky+Zs8zUw91AiZPqdVVQjaVGHtUSmxviYiQa3lCMqNRvMHGlrkUWwv+a8opiA31lQLBe7
EHtzX4m1ZiTD3qQXcexbAEmEXluOuh/P3RUZkhJCrZ+8mVr4OqyaNxCjF0ESPyeD+RcrncXSjImS
Cc5lNVX4Humx/pBSE0d+NUM9wgyvyIy1GFpQmVqh4wbTf7CmZzLvh92WTcezJkZVEZzudiDVmn8s
nGq1CDG4yyD2BOT0jU10IDsfmiRYjibV2lkwFL1kmie0csoGd6Jt6rE8d7Z9XW9ltQj3DtbRuaQQ
ncjCQFBOZ5P12z3MBgYkBEpDA7hFRvmj9Vp9O9hmKCKvZpnaIeHzi5JVfRa4t7Clmo90vzGx34mu
xLBYDAZTWDtwMXYytqjfaWEoYhpTtmaV+ZT/ZNJ75/oh2xXK0tU88CrP20oP9eQUTcHXVbDxw0GG
Au5eJi814mJqYZ62lEqoF39P8NwWHMrlF+gvfjSbWyFOfwAeCXVZKbz6Q5MqQEOeEZSH6m6sGcY4
5Tec10CYQgFX7k2bLcsJgMThyAM9zM8cUFekocEkiZnMdugfA14g8oNxcbgPMnpzp0C9/qQccyth
RpRVUQ70qxWg75IIzURInix+e4g+yGohNR2d320pBkcMXXiTkT2OJd2/Fn5oDu314y0nu81hSp3Z
FVS969ci7m7hp6KNu4IjXHA7GyGtTBogRWlgAD3Mhn+v9dNIYGx7oNPJ91M6aPUj3bUeTYFWAb5o
Tg3K82eJx0x2EMfe6CC8WJO8/c75zd8MkOK8vF2NkKv0Hgw4/vorsV0aWD5O/emkAJ5De9vt2aPs
sRsLYoRJNtvJZhohK/k4k7SqFDUC2xanz7Aw8cBGoIakEraeRooZzAPXwa9K6jrfX1ft9X2WO8qe
zSc9pH0jVygovMAWlEu4luMdwWT/zQOWI1yt7eS7/5TJGyPvsG/MBbesd+Hp7MGuR/oXn31ZyQuQ
iLiEZL+qvmLaBaS9KDctKtdIue8K7yybHX4U7Z4Qqj7t8rFWoLZKtpxYgyUyWnzvR1K3DKJM0BkY
10Q8O/i9d9QiYBDg70GXQClUhOct3pQdnLPQJY6tsuI21683Nv0UM7+hLDirQJ6Qgr9YDHdRal1Q
/CmSZ07jSZIVNTDnWwHqXMYI1myulvb3WjI+uxwBlhtymaWpkWUrup9x0SECZa/vt4XWVcFulf+J
wDnIQeNpc9TVwrLtytvTtDDKBKiomHlMb6Fmz0mA8EswHsCyTPraeziwvRj+gNVTHYgk88xQS7tA
FQmrLQEX4wVqz0GukLDqt7lDQgu2Z0z6d2UzNtkpVtTWEQ5IjnlF8wqq6VsuqfBOGNTgnUM/GNED
erGYgcrcmwYns7xo4Ln9mheHDSZ/cJMhaehWFz4gx9amQbbnqAUuMU7HRY4zAdIw/nExXv6UcUkE
poN6fyoJrKr8YJvRscuITgo1DHCytUqgp+skoQ5cETFALZ9TNes2oDJRBwp3ua0fMoCJGyDtyUMh
ZquBEcrjOuJW3sKS6iEs8quqqPXjExSmIhzvrr9SNH4fy7fbznDMnNzUKqlqb18kxJjAKqFuSBxv
FfhzUMFXptEb3irK5kQjez/r6b/jBh/B2g/3uhoK2IclugaiyxHjGZslzIy5VKzyoJ8kCBykc21F
fz+WUsMjWEm6Vcp9j43jGSMDUMQXFhaltSFvIbwJVq1zqh1KccxUv+8sQmROclCX0EnzewsZDiy7
c9EezkoHwMjkzWb+dTNrTXXhIX3mnyqhwOGT3jPdPC9H5m3xyd8P3VcEqp7HcoqT2rpGK5sdhUuV
B+Hd3MvvF73LqBM9S+NZezOn6JBKfvTXz8zBlDJwVHJVU57l123t9gTi2jBs+sKpWQW1x6Jd8z8c
4+Z88MMpHh9q9P9xDJ0IsbcxKUV9nwAADLUwlY2+TYsgVf/mC5F9v49fnbYDNiGBoM5kx5XbNCEb
FdhO+VhODia5dunNp9jnDybBs1BwMW56p++pOGKzxbRVLB0gtqcYscdDZ9parm1IJ2EJOebxnCTs
v5YPx7EjgSGThxPtx+dngdF+kW8TPG0kb+tvmxiqhQ/CvvEI4FtVS1KJSd46ibgcixym4i+bZPKk
TvcAnY0bp1kPKse8rYeArtAW72QPdq230jzY688ZfqVHFw1IHZizxm60lJazR4tF8/tA47R801kH
B8Z1rv+gNxxJEww4zF9E2js8FSDvJt+8IL1ugXz4NZx/hE8XGJxjUGg4xc7/AbydniIU6T9MwsE1
o6tp5q/i6SaCO1pdUWr6jO3BZMuEOxPHEGbT4TXz9zfNu9etY8U31DYMy9RrmNSRAsTUo6UI3V97
a+AZW+TkHKROHRpG3JqgNlfyeQtjqjsQgwEh2i7v6/C7CQ94xNVOipoqNdAfWOyiBlTUUmD9h5GW
pUGf1vrKz9TGMT1K0xvrQfe04MBjyRpjW8FkIU3cg3Ts1VG2+bg5jJMdb6Gda/DV5DGEqG6ngAxi
hxKpO8JapUAoiVxKqc8ivAFksnlT0TTHRI60pwAjNfB6926HMGwzKiTCIB7ggneYEhpeSl88CkXl
ctXEp1mC0oagU5W3PNTp6fFy4x1MDXDbSC3CD71BtB4CG0E9ERdtFz2lV4KVi7JTuhrPZaOXfV52
5RQywsUWwc5eYDGuVq0KxLJ2MxZGXjFzj0uwxz8IHOYpaIEeBtJFLKsHJDPIYRhLe+ZCs+htjGz2
tHZU7kF6YzDTqvTxecBQlPA0nVMvbw3ZOmO3czXmGsJr1pvQJP7nX1OPXZEPItT4pWc9iWmaQzzf
IY+16owdLXMdcgNkAuIpDaegz0UIVZgZF0LkKU1eOZWK62BcfRAei34STrwRuyxqTHOjyXMToTsv
TQJZAdaKHnBV83el2iSv1RimxziiExNVeLA2xCO96zbk4cLJOVQ85teHrYOeznyUdOWM0dZ2GklB
biiswukW/LDv8jXz5iJxYyGFxFkPdxODaLEcxlWIzyYzhcKEn3FqfnccM7VoEhsAV5My7paPiJdP
D//k448Nye+GVKrFaWIj1o6gmqW3J+hn7x75jEiZqNZK1UpH5PVmhcZiTQcducJjgEkLuaEQoW20
iCKM048tTJ4sNqi4O24yx5LeOMQuIf29FpQhnIW6MHerPZhboVtqSZY6muHeZRQBaAjpikKshtk3
JLff2JDjbEK2mMd91jF2X3cKjy5yrZ/U1JMsfTkc1u7p4UStqgUdB9zMakyysI7sLr7YJ7Emhy3Y
YhwIuRFQmdxlr87sCYH4PXkS5IEkjgH2Ai1zX/orjEmQ7rCVIV6gVBM2UTA9yGtBozN+2idQG3k6
mUMSgenIXKZf2kKS11sV/yk2RsSgIlRDijssxVRwYvaH04hgOXNcbWEf81zfb/6vd194YCXe0MnS
CsWEEBwyZpFjL9AGsfht18X4d8KtOXy23A/ySSEeoSIdJGnV5E1U5AHfqGWx4hBE7f5jlxBFHgR+
JJdR23WyNuH/rs3wnsRBwkA2fYo4NA6ntY8uY/dDNvBW/U3F257GfLmUaqkAHBsXxfE/Oi6PbTLA
NSRxqrMoRMXHT1Fdnniw05TutHjL73Swwgl+03j0S9zkBKL5o4/oIW+vSFFPHtQA9/TlJnlcamvs
hnlwgkUy0MlPkRBLY/08hXXHUAQDdI2Fq9muomljS5Yp+ac1PGaBa/yeWJmJKeNGo3P2O/6w4sSk
wode9qs2c9oI0HoD7gYy+hnHQp0005wP6JLJJQ0JlO0Lnr7REf4RHBE3Rdo0nfS2OZBZNPSlabj4
9sXkDJUNFLF5LcvaVzsEgN1blSapXOuouf/LC+QPK6T6ReyXGnSUiYVshZKMakM3jFqhKpdZlk17
0a/1DSX2eDDhO8EwkE4kALnq3Kg3nhrcLxt7qAdOrU0CTQ/S5dpXUKRx9zjThhT+0JhE+MiQC87L
OVQcpZoyqgBwqTc2F1KwQnhPG3a/EjIHTZBTpXl2ae/q5NzLgTtH4eZ8C/pJXN+ZM3UD4m6ulGEp
jXyp6BULSHvUbHYW+f+7sq7jvUJrN11z02b4sKnCkTJDsQW623UngmqG/nd5sykt0IaWUTiYnnLQ
BHj0OnJaxgRoyNBQHQIQd/vkzJkgW5qWom0A9kM40IDLO5hL6iTizQOq4bEW6SWM+iWOH2dUkIQD
hg/ZGB8eVDQ2Vwb5ojUaliuhimR3H+QBRZ6AFe+cxUcmj3rmbzmIt9sRcIaxPCXUVwjudTpLnUOH
wTnzQHb2TaCGmCgKgSLEpE/mq/QoXr3s2XYmyV9Xe0qm05pmTsW9UyxmVy9VHwio+M1S35b+mJoM
lHWN5jsFr57XHxRQv13l5o5veIKEjqDH5MVfqmjl668bVkkX9jKQTXdGfq+1oP1V6PG49jjdCQup
ovI5gOSAJ0XGL/RPjcvubEmZ4YeqvPoIFFB1WfQbMCCLk1eyi4cxe+P7hp1jNBDnY29QsEErv4My
I4W3mz4SOuNsr+geXIKXS5VD8PuJsIM8Uknb/WZIpm8qYuN/yqmMowKSClzhJG3wV9Gi53zoevbo
JjHNqHRwKcmwBP/dk9iI3X12qcTGqYfPSGvE5r9cWOZya9sB7HLmKqBYKWoj3wZFOaAPQm3kWSp1
rzZn3VdEHNYgRTrbaUIcJX8aQca+QBtwUQHJFELiyPLCdXSl3pvuTh6fZsNFoXbVHgYQ9sBHPVDG
cxfJNjy8R4YP9FBAYJu9ot3rWFzM4AfYdwOfeaYkm4J6haY0ibR/imT2tYETbH+NHsvOD2AsuEJd
PdbM9yjAakxggWPflzsyKgh0dXycrZ1k+iPpv+s5PvsVteSh+EC6INdzLdUK/o2Z1OvU/IBb40kZ
1awdXpsROjCtXHoKGsmkZt8NzYS3tOskk7bhg5oEFr2bvn3EsH1s8pyp5w9fnVNrKd7ckWkBlXZm
cQclDuNRhWNsHKqj0j65YlyXCmgkIRoAETfGP4n1iTn9ZKzQBarigaQWNgelh2C1k562bcMS+8+w
3tSlxhombq7wTMpfjou5W3A7ox1jKq0BPjnnfEochbEj9L3rZ+fi4hISvnmESeyZWXp6fbP8E8ZM
KbiDBTPFUSN0iIdpIagODzM94G1CdOtZKeVzwYVlVCAGJOliLMALMYDsw3aCrzTiZZ9SlymfAKDM
SVcl1UQQ/59THlYHZusD9OROtwlNR1wQqCbEB4IusaDVM4JJf4TF1xgUU5u7X4CWG36qlM+Ktdi6
7+YKUFTjYNwElI+rtjLKXtzXtUE9wQYXkzkQn5x90pPjRvkoaicLBrYoojs8LGkcc0AR7PyRWEfc
smKtWtNWHZki8c1+ChpLa2kfXVTqwWaOibedQj9e9I5nUMPSz/9wwD61YsKJ0JqkUVCMGfddILd2
mT1vFJ2hEkzd4cV4j35t+DlzQJ9gWV3pKG/9vV5hA2uc0iVqFtr2e9kT5kv34PxNZmgBHsns1Jk2
Ek+FZYbxXz6M3hqWjAP3+BVVANaOzG4Sqm20QALawxJlNmKhVhRFqDrqYEzD4bt7HsmDOHmPFq43
bzmviIw5ffBx7vI9HUOTjtw+PvvjrpTYsiwdsVRVQEP8q/SaBodUFuI9XDZv50l1dlq7qn4OX6Sp
+ep6FNj9SnR5BPKvqm/d0Mufr7RVtmEk4i02HXPeSrOrnZ4g5NFn07qBKfatmAWxI8Rd7zQ4BfHZ
YawOtI+cXod/1Jc31ChIJw2hhDvHOJ2egDNEVWCSLcPl+cAxWzJ4RJ/7DAMJ/NhQDDUxX5AIMYHq
fjGZuev36UQ64fPjFK900T2l+Ub/ZUXGNe0FFh9toZysK5Vcx85a8ByClTFJSVDbxZuOsd81k7CE
TVeAE19VPJBFgn0TP3jZ1FmLFgrG7kWLAkY/g9glmre5XQ8+nen7adteBR15/2iuKQYo1P6oKOby
1idUiaLBVKmlpv7Z5LMAcNXxtGvzZYzHBQSD20GDs1DjwF+l2mGKnL4PdT3bBobPLS8MOnwcsZjQ
zBtSr6LEbgUjd18O05wDon2r8BknEHpSGplL2YNP3jhuIih2LQQ1KawPQOESY0C+UR8430XuYFFg
pIDSPJMkQ8uPL+xaxp+lIEafy78pXXyMacJQ75Q3OKW0yHAADGhIgg401Vn9VdU/rAsljryr1b9I
aUHrFNGzu/aGbI8cZ9Cfgj5zOfQ06FJyTjbG732jbRi2MTwSkfCOdFqIEeZcGN6178CPwEK8cNNG
wtUyBGUgBC1iuBGsLXF8M57LFOdUriHPjpyM9fJYG+Rd5X8WsG83yjjTuw0Bv7uFmbqVC4PnRVLz
VJUkB6rpSiXf60uO/oqdKSGnSheOIkDX65uD5rdVQe/6yH3JFu3NSTez48DFHXSgcnVRpOqmn6+c
XxGUGZYcTuI9xYOOiLCWHZ+ugrPU2B0I7RaEnfbFjffp+MYlmNUM5mHt9SeENHSIQbYA5DpAolFW
XDXjSnAWSXDPcNBWMw8NOjQYbrdDKjF9iVS3wtiyjKwUyD9qMOYOIPS78f9ZjKhT3WLeWbUoPoNp
Kzx3bvNAGOEuX0Iadd8ws9WUEyftmugUo/v9UVrhhtPq+isggX/NJK7yAhy15AEj7jHOmeVul8nK
iAferIcawil6RcHi4HIjIxTn1IiaiLyIOaUkutrkb2w4TV4fXNJrR6/Q/xhLt8FNcCSxs3Htstdt
6LCviHDkm80FROAP30tAtiEkXm9J+5NZZ5e8Rj8hIittjAihG8KJPwHY46tKCsAJHFznnM48620w
T865Q2nPPjOMunde8NfOsV6tlqV9KYywgRAel667/iiON1IivkUNOAcYyhZMV7r9kgAQR08cp6IU
PWqNzl2aXy3QSvgNu+S1aLf1KAo05RNjjc1b5fxfB171QmeQdwnaM3Bg2JDn/aZe4K4UdUHMYi6J
d4L3EDHSwTkHdDiaRRtHhKlEDrEa6wyqNISd5dJo4wI1XNdpD/U3F2TuzYVR+MZSCaytdIJiu7wh
ioesQQvo2WVq6lGwL6NlVVnMOaFvIhaUAzuPTCjeC0iGtbpqbCtpR9NOygdAMupNQ/1KyDR8iJ2k
sqOWuC/mETK0T/jZ5B0hrc8pl6bVE57jTktWW/zb3rP86Dmk4w9ToZuLUhZwX7pOMuI7jA1/cMMX
W35LFQPT3alcIkoZYgOb9x2S/NtQ5FDJqyzFzEzw4RnVzJyDRtl5iLyW/qxayUIFx8AZt5Gyc7vw
St6rb45B0D+XwU6tcCLH5RVymtDEBLF0T56cgrMJWjLFt6iFq2ljmHrhmWXYvYn40nhaa5mNemzC
QU7Xg22V2Ey6HA37cbWuNXFR/d9tj+cDQ/t6zelPk5+Ya4hEV2EpMYr9+5eshnQmRpGwO0JDyQC0
WR/RFTGkbYG0nNEMRoOCOyl9Tc3UITBD0IIL9HwJIEaMgMM3RWw9+HCKcEJo2am1ZwNSpu0V6htS
eToQFBImCWTBaZhUOrWWIG0d2u0dkuTN0iQpd0+DomTbr/qPc4eLx7XoXZNBkZjjUU8KvdmGmtfM
i/q96G8R5YANg2ONMAhO/NYq8YBFctnQZFW/ONubBSksnUXATkd8qzkMC3mxA1drJf2cgr/E2Kyz
XGHK0xlwJxoQ1WcDh6Otto1l/E3+l1oEOl4oog8YoLkkNZsdOTmEE8/apun3zq7eunaVw1rvXqVX
gkPt8V2IaXXUt3ZGsJ1hZ0/HS0qIak35+JnzIN0zz9YXtV4yC4YNnsEVUN7Jc2YyuptYw0qg8OtT
yJ5L5dzmiW56Ljto2hadpo/zdNTto0GJQu4GDFTeq66im955S+WfwAOGYadTUX1SwpPXHu10r///
e3l6SOJZLXaqIygttpmlLL2C31vkQDOcnpQvmHIhkpo3FGEpMn0T0UvUDb7qOU9/IwIpfiwwCQdR
0Rj9JEEzvk/9VPqnx2CupmmHmKQiRxfjH7g1ecmCsxdcqp19UJpf92T+nTMFacb7b81X49646hXm
Z5uDGViAHmnndN5jdMiqrVjySvBk1vG3FPIVu/ggcgO7InAirESCOSREbRwNKJOKgO/YPLRn5ZCd
/3DQ0lZMf6/Zsjpd/ObNCO4zXQLQU1Gf1tnsz3ts84IfC0eNhdWqwinRxKX+6hlgiUIor65bL5Ki
oknmJWRuZ5rnlmqqOQprWWhpEgKyAxsPiWunmESbdePpknz5/z/RCkHMp/Yj/YmQtKACMPopPHNX
cAXnpjRfz1h00Z2wP6R47kU0E4/lV04l1sVFT2qczFO5ATWrHlp9E+zgieYpbQI1fZIufpPazrSn
8KkK+wtTyDCcvaLnlnP4p9TTS2nU7jnQEyQjkCwXgbMWXH4bW1XVlfIFj/FujYO0QaDKCkff4lLm
s0zdnbXLCXJy0847UR7YQA3sdkdV0Rye4dURwdvUTEjIfRACY42oM0N1YNuU/teu0Be7mMIS1Zra
EBe249NRxrA8NB9lWSGRIZwtSkMbcM1vBiefTj/ITa/C7XswK/MuhLZRtF07FDp1X4PoAHuUoPOk
zVbPd8wbjw/mW+TSBkD1LJuR5U+HqNJQQtBgWPyMnW9A36aTsHoYcFYmR5u+9UKruY2Zzet22sA9
JGZBeJYI6eE69l3IaaSPjzyiDeLLtNTTAcIV4OKdzM8tCWJ5tbC9b58jC0seOofix2sm38asCQed
+sbToZ60jLynz6W6aZMEV3rmTopvpzAS0AhiGkg8y0skcS7YS2hOvHEsqf/kBDDVSjD/l1FR3dqA
eni4RfIAcNmeCLu6EW2i0XGnOvUsGF7lNjFoWAj3ilIu7OWsUpco8X/iJtGh+vIEq4i6GTW7V15x
/niQO9J5LNFBr0uR+cNdni+kSId5EmQ5KIPMU3e4rEV0lUjadHhU0GmBtLbh2H1gjQGRdHvpZdew
Rn1x/QIQZNX81tg4+8EPa5GncAplO6ZMLmbHugIsqrCVH/NmECuKxm4DCB2Yx4sPZBuaDONdHjX1
HDC0Psw4TWPLiNMU1p+FJD/v1gN4V1vqZBAfvzWi86WXVuLnPJ9sGFWoz/1xy9sxgdSrzCCQgvOo
RTUPN5Akkx7mCC87F/cEmOcicjI98faaGmiIUMvGTNxtxdEpCGtVdY3wSdsmqqztoWxeYgJjigvJ
l6/91isIlYoaJCIWPTQsuYK+4rhw4O2SebYthD3GgDIf2MzcmSsR/UgBdu3yIHagsrVmxUFGQWlK
t1W7/iYtLNIrEG2kKLvKFY4EOQOa0Rsgc4ur7h48Yg6JwbzRXQzyqrgNqLdcr0PmQlTAMp3s6pHH
PQGoMQU+8wvQbkDFZ/A2raJQNdAonAOpvOelweEPqech3xSStQU25RzoZLTZloAt4drWuqJwVwHx
Qjml598fPJS6heqjxJ+URoUdU8KxeQXrFXhcWQeHmAaP9/dmKTVXPpcRmStLXquYNVJkrVVUI+VO
a98X3RYrvLHdW1M/8dwH4zpKZ4i3shCQ0Yo419khBNzQbDHw7hzba6f4/BVafbku7zaFSv9UDWKw
oQgdQWbegdhY7FVed/zLN6TRi9nacVp+0vxelLxiQhWURfgWTfV2gZDQ5myZB6krT9pNA5i5md67
ga2OBldMjG51xqcflY1Cru/dEI5JQKB7cn5DAualsAJvisrhQIJ44/S8SouFF01ttSJKkJXxvFyz
h9pEqpc5iVEQa4n6vCWa3NmIOjDIwa/ye/x7gaNe1WkmGSMWKSaa8BvI7d4K5pGwjxFzhsI6pN9g
39Iy94sWLqED9E/nfyXQp74JbQKilxEDXtUxdQZM3H8HN/CSykajjTTMSkNMaFiOicypCOu47vCF
Kz4oBRvoaEF3n0xQvw0W8vzspwNWz3mbEuIXuyhCE8fvd5ERPb9C8lsZR9eQtTycWxgi/Gn+TK6C
62lG8kVLgAkqv+7jLUnqG0mye5DzhDamI8Q1clZ5o8Q741K4U8ptwfup/AG82YzElbjiiOjHurmk
4lcK5iZnm3tjLjOvBJgk85g8y3lOs+yJ1cfso3lowuwahK/2l8kdZ7k+ZUDIUZ+dsIJakfYdot63
Bypg9tGzQYscPv/9nef4uWe+nahnUjUIfAHTaF+hOHAM7TgzW6MkRX6Qu1lsIF6esEh1+kWCKitQ
mhyF9V4qjCxVZsK3u8CtwImb1Ixe1lVamWD4s3ey99SKsYjulGI9PE9mqLbG0zHJrs5KlaoKzPpY
7KK4G0kwXoXUamRO0g3ENlbl8Xw8gsw+8h+fA87ApuSZRd6oA4Rhz0K8kuxrTrFJ/FeKHwzIYjGY
eYZYCacwY514XpfbYYiUu2KfSHkwsgeTholHItxpx0Qwg6YGvShKnaVbaPUVY3GKGAOzmzOb89Yr
Z8mqf0qSNIbKubZWQJ/WVqkxvYfrcu/dUikpuYCoueNLvIHGSS9x0MuoKLT9L5LuuzMFhkmdTNQ+
G2n0M1thOCRri8bUUXSMiIQqxinMD4cdiCXzW1DIKsCKQYq2Ntm20YJW1jNwtK4vwXfE3GesMFeM
j3Ev9nifLzUv1yi3fMMIYIaXZYLiWtt2Mb/5ayznLjyVHFc6JnBms7ZvpMnf4Ma/OrFIbjZi6FKb
ffpHOhVPRHmn3xjTx48nNb42RirM35Tyxnc+CCL0DRpnEUD2tnu/pPuq+pYJ4QGmdLH5iWy0BeVT
H04RpeheojSuLCHPzYXDu54ffYRLP7SkMgfdWSKyYiBbXgBmbiTpSGQOZTpy+e20RszTi8yXb6jO
tiJTW+srjdTNv/K8H2E1P4UrlfUdrCSfgJCu1amvFjAmsVgg3VOzbXarF5sGCiyt5XOX8TRe1wAS
jNzDrALmB9vbCb4YrTjy9bxQZz4Zxtnl7Nyd30kUkN1l1d+jC7BFdOi/IqIoC+R7h2vnnZldiJ0x
SNKhNyPADrRZdcM+mq6l5G0qKP0n7CCU5Ur7+luCmUhMfukt+O78VMObDUEolTlIOoxWmlEtZFg1
0qySnFPqQiGaicnYi/327Yz8WxtkeNTkQLKDmfXPUFOpTIXqPQ6JTLwHG0EeiHLNi3lGGMESU03P
U5Y2ax8/LpvVO5LpCz+FpsCHB+SBJZYqX1uFb3DnestuSPE+hHw4xJxqNH7uJd6HSSgeFSANgz5/
JI+JH3Dz6BmMXLoetAWG4kcydFmUmvJ1N/HMbkHDCwS4OowEHKS6l2zSnbpWKDXxyteO5ZB5TtjF
NPrw/8hERuRFq5ujqId8R4KWM5EDeh3g4gt4E/yOPoNF0JRxohdPov7APPzOJyWor3BeIlbXIw5V
HHHXNOwGFL/ChIVVVHfZPobCXbooVq6zWB5ci9ew7I0mU7QD44bRuEFwjX+qoJy4Q+DO8nEr11ng
r6iwNkD4CS0Ni6spLonrKwRbNwrYYSQoqasbMaOaKel/QbjYD9fOUaRQ4JRVU7KaTD+s54zoiKn3
VGr7l8k+0NxEe5YeJzpHxJPmpInvSdGSZ48K0IWc91G+6HqvupyZgG+XJxF0mooRYVG5rX5MdgoL
/G66Y+Uq7WYUnOiXKit+13qrHh/kJCQWxsyH179MSRM49vBBS03FS0r1WrDX6tdS5NMJ++wk9+Bf
DNTDilra+t4zj9AELiMii0/XYEbGqskHVgjxxx9fuA13DTot6qjZiwbOqMaL0kHcAKz6ipSFuno1
NH8q0H9jYTQIMMmir2WMA+uUKHGIyIPokln5Rv+VK22soyZvOU97hxJuVWCX1W/BfNkixeIc2hmB
8/ZUtrqswe0+r0/ny9+gwnxb6XKHENzewcMOirjYVK9STDkv3Lwqex0kJsBVJap9aXNXpOA4+d/3
CHzCkRHgvEe4CM332+ylbV7dvNsZVUa3dBEA+WAGGkCO4616Lq6I5A3ueEXNJu4ZJ+VnyApJEC3u
XEDyDvZDoSNVHe3yAek5sVWUKBJ3bVEVY2JVRSSB6fC+LL/6c8hUmAuhAcLJoOTv44NPjvAqeEQT
GtSWyBwXUyuGmhoR6MJ/b90/5fal44Xo1A4L6pSqQy9OHLk5D7AqsyGu07U4sTEdDcZLx4YUlWS/
6HCK7L2AmzdTPJH2OGxUCoQfvLRRSWkvxouoJODJs2JacetVb3yStP+i29V0xhdyoFRv3HOkbeGF
zMRr5v2XoKJaI/9FgTX1On67yq3iVKDBCzue+GJIvyfOuFYDfGAqxZSe46s2H3Nh9jmdXc926brU
7SbtyOychyTjiP8kkirwd6tLSg7p8Xie67zLyoZWpqiOVJdUlS1hLkG06BvZ8GNMKPJW3Hq9qcOA
5U3nBoVSSuLRLfQ/gbkypiN9uf1+/kmyc701tHZURkny84w+5hatxZ1t6Z9VCIPSkT4lrAcWHnCZ
pVrkcYhvKOfRBe94faXvfHVtUieEi3XjkrQCKCbIOKAqTIl6jBiifJTSHfnhm5jNy1lXlqvUu8y2
Mc7Wa87Ra14AnzZHTDp8IiIijc+1/gRTGyaL/JgHVBh6OPaosabpWnreyhGq7e12d3ULf7z0pP13
LiQK3kxXZ4TxThwkpY0cSvmoAkGsaYn1tcaL1Yq92QWb9v7Kxrn60cM2vs51LJrp67lKTQJQ8ae4
swdc6bZ00RaPN6AzdilCiu60g8ttEKH8V7vZr2BE1b4OLEjCkXvvPJHmObGPO0okuJy7Yv0mikln
+IDhCXHldXEkbX5JjP3wwBZssntucVP1pfzu/UbMKiyfeBww8G67B3HHCgsndF1ht6LC9KKq/yQB
5XxO43mBKwnUymUpqTanJNXGOgdFfnjmO91WWDNDDr3ljjbE9HXTDo3Rxvi3FpFH2xJXFFrUBbGQ
P3joFJZay4GyPBPyHeFasb/3AnSNcT8NCPV5RYmaDqK4BX13A7QHe6zTUuRcxpuU4VGwU38n4T0B
T07KTOARyZqTRybSaH/5tf4QVI9hsaQMs3Ob69IwPoaM57VI17+DrfeK/JyWLhe71AxYQoLx0Tvg
/0h+llBrai3K5Y2DAb7rMbB0AGoQc8li32TfpfjuTxTDzUn0f/2BoS5ec7dbI5TisWd9O5Nlhk5R
0pKAVDa+uflQLfvWG7Ea1IvgLGBSbEMDbTYO78xKJRbFhN+Isav5NpPOBK9quVtVZj0V7dE6gXx8
2spJKEz5uvuon8wSWAqcHkys856GJwOeyPmLLYyr9PRc2H2XCQ9K4RfRI3inXcklQqKsZD7HEeue
XWiVzVgmW+tAy/hXxLQypOBat+QUKcmTC2HQ9rqU21jVJqOQztnLDu7nyATH6DANDSrYTeHWa63I
SawqAFHSFJk1pVmIiC5URND/q1cQXY4VRahZLzpnlXxMr5I4zMp4QdIf13wnSi5zuZNoijidz7A2
h9eveUqEEfOyuP3hXJBAvkT+dMcLD0Jug7H657huSyihT99qiFQoTbAwxrCKE+DAGCqCFwhOJEvp
E7kKBDSKkGYRNIkKRpIp1fx6wZ5UegCrpnxhj+GTKRebYUtAoOzGE6ZjhmNOGjufaDfeCMtHox1m
Xi9HKQzefgmPNTBQDeDg4q4pMcWY1s10fPfRUF6wnAeJO1GhlVI535Vu+3tfV4ZrM8Dd8zf7tZw6
SJIAq88akjAMgoRVk6mr0pbPpYwBO/5oGtBAPNBOqzOife2aePTGQnGzstQbfKX4973M/SF7Bgc6
m6YtMRWwiW7iIWEeVHwF02lIwqs61GhBh8v/VXofWPR/Em+DpZz5welVa/zCz6Eh03TU1uPfPBk/
Yu7OIyiPqxq0pY0RRetoWwehEcIXqiWzz68+irEtP2nTbXnyPFNkgdW6BhcFtXxirNx8rV2ecXHy
1RpGY8tNFSCQ1jxYv6tw0iY3IqdkA7NZ7fsCBSFjabtcDPQeoCJn7ZHEh9+ZupgOTs33sy0L4q8n
XKo0nt2xMFgTJ0YxGyf2yShrrDkYCtj13KCNSc3N7JhqDmxVV7ay3+zZY1XFCuJvRsnu5vvj5+eB
C3WQVnbeFQCez7k4ytAPqHJ3a+Rtxgv/HVp9w6B7Xv54yDWVdmfUkqqD7zpW/AUtIKrAATCx/C9n
HMEYCjZlAuMQc8iGRQhitkRQeWdV+RJ3rsLrsUzC9oLJkVP2mJ/JqBJouAVkB+kswz87Rqtoiaw7
+Rt1+V6szUN9BULiAuxUS4UU6aJiK9XrIGWnUUKpsWjCCXnnJ0gWvT7ES4tHSlne04EGE3dxomHo
sXvwDgmq9J7vTHuWNt7hL246ClOs2yfK0hEc5JnfZbQBcev0dnBKbxCinVGE+C6oHgLcMKwE/BEs
pTOQMePxnWCjVJtrsfugsUMePZxV0MNosFspioF1tIpDWf++7SsQFcxNvTEhgSS8j+PKs8IfKoIa
LN3tLJwyRvEQTvzI8O4K0aW45HolG3rXsAPe1mPYXfQ2RF9wu6rvqkYeOM0dxZORqOXgl3+84rwn
HWBkyRipWAPoHeoYaqg8QUvADCM3INEQxV5xfktp+hYpmL+TPZiMuZ8mSN3UmiCKZ5yV3dvCAWsY
fKEWH7N1gi6wDiHB89ZXI8BLtjWw+e1+IZb5dcVbN6FkqxdsTtsWjyBXZFE8t09OA8ZNB48HL+WA
PYHBrpcUy7x+2vvNfzgGy/RofCynIcMwqjmL8cNcoRx6tPNq91vMiPbPf+AyBSMr8enzBkRs99lN
LeP3RjXWaeibxKRDdWJyXICirGyRmRf9T8UiqkiOpZ1zpqdzRhwdizJvne6VqzEGFKnglvMGRjJh
T2KXSSS5ve5H0URmPyUX+WAymP0QUh38u1fjPA4tboXFHm8yNLW4R4B1V3uFAW9BZdkR0UXDMs8a
qIijKWxw04dLfLm853RlK9qNE6PO9M+d9XJ6LnxDKxPkIJLBjlazHzA8r2TDLSiBU+EsNvYsDUhZ
8SZzwOdsyEsDy+JKTZRrKZxegL9to1yuML9Zti74mLHDn7z/qiNngIJXIDVd0NInw8hA8afnw0Eo
Iu0vTLw0jKpKIhvUYnSWgLbO0cKqSIy8+GZ7GK+l/7lLJsmV91ChK/kWWHpz49ycL2KvLPqnTnGc
Hh8DBM+sZChwd2/qSLYb4G5NmlqwWm2IxcRd5LS5fpl3xEhmFxMtSgzKO2Mz7Wjg7KD5/Oeb0fbt
HIqAbZRGTsEACV5bQjm/fTu/g3+xN+rZVQeL6rE93diEuEv/7/5egdtFhRGR9CWB1X3T9meuFGMn
eBNwMmmqVZMGbmY4J3yfSgfPkoToO8cyGQlLE8UPAJk0hue90aJ+Cam5SrDpMfNogMCkC7zNMbuz
VVYm4pZEwVrRQN7gt6FGGpbPqGBf6ZBLrsWRuvZMQtPzaXw3dS6PPPyWj43S1f5hiMd0PDk9RDPo
NktOiYXx1fsX1/Yr9sscGNUdVZ3vSPKJgnTKgfcaI8BPNKH6BvcGPETpGbFhcJ7RJgDGYdiGY6Kp
kL5EG9y5L47NmnYSlKS0pFz9aAH+UUYx6JIS6PdsvKp+7DZgn4mOEtUWT+oZAm5dmH6zktGtTJ2g
FrVb3Rx8+zEaGf/rVqpNO4AFTcZH0M80c2vaPNUM2UpRXXGEPlXrbtY7hSayM2i/73W5Vn/lohd3
wdkO49o9S5lneG2ei/L12levAHmrG7jEjDr1yL/kZnxyiLlcJtUGOz8qNIAy5KF/jQib+iZDmuOB
xPu9LJNc66iCluo8s5NHufB/oDkcOaVk9sTxVZi2l/ww8DON9X4YqlCC0/hxdVNYQjyRgPgE9cvT
e2h38Fe9qpyTUQmauoGteNlYOwSsgutBoevxyvzn5GgHPUgvuaFXqXj+vJ/JzMB6kGfmOGMRzXOt
AOoyB2l5aY2N/m9eDd4kGURByEzA6nWhB2tvgsG8E5kbuK6Qhjs3Ut2eRn0LLqXKjOeSEy5IpeVo
fuL4WtegePS8WqZgBzW3HThZwYZIxMwjOIBpqZenw9xRtNdxY6Ou4mEJ6rr+EqA/Gop/ugeBYaxf
Pw6KPOyqB1Ttl05LJ2J86684Z9XnPLqLD3xp2wKlqSOvzOUZDgZ2aFKj1t0t4Mz2IwHNDONLWKG/
zWRmaprgN8+ffyas0c7Ac7tbKbasbnfv3S9o0HviS86Sf2vfYQqvkQgDc7g/OGkv/4iKj80sjkTN
doXvCPBSRJ7zLgWz4RmjeeZmVnm3LhHh2WnUiJBRU1Geu3kzvhMU5W96l+Y8POLJjHWqIEHAuLgM
/dNLtFjXo2SYvvE6vtwW9XQ4p1uEy+o9p3youAnGV6Q+KLHw/hOZWu2M+qzQyZInj6HhuMYNzoCb
CfKlixk/TSe1NFP5qgVjU7svNiNNj7Bu7/XmlfzoUYp1Dt9QJxpHyivrrGIMpy6f0LOfVkEU/2rX
IqFcOs0yykV+UhVxy6iBE/fy/xTN+5YLHI0iTYCbZbzssSc/8hfgwd1BUU/5xeD+++EqyWqvaRro
a/sjUD3DvRkz6vrLkXgtvQ3W6h4sQ2FhY+ShwqBKCKZdT8mJZa6LjrdLV/xMfH0c4irGdr6HBSC3
AqIeHxHMKPnX8GnZ8CF//RA1meuarXynNGuTOGUNYVYOjMyQmevbHzBxnFKiM03UGTfO1umdqP2j
Q5btA2yeeqmqT/Tu3/FdcqL0u1cE2XBiW/I75H17fX2BowPoBjs+Q1g3LNCkXneCqPTVHJt+IYsQ
aBAO5t6VAelf3WuNXF99Emw4GCG78ZNpNj9fATXI29zJkZJZTROpukDhXTjHqc7KN7HAQ61A85yf
saMaTSDwchoNOx24YxAwf1LXTCOzbLY5BSHxuzu0PkjlSqnrAT59EEuhExRA+QC4zqtKs81FwcYf
xkFvTL3WaomJd36+7qJJV1sntHB+5xTgWZMtIZZVf0R5fQLrggoYgxlQ8QLTxg18pEW7Vc9fkhVW
BTGXYNTK3BenJ1MCBlAGEEA2dBBsRcG3sUKkMQ5KzeLbaUNkxvL3i+A2tambHj3S66bcDcXuRQWb
P6+BmtuC3Xc4RfElIJWyenHvbrfnAvP3Q5ZP3T3nCiPwM7TnrOX8kf4c/RZH3HbPcWDM+3RyCRun
MSrltY/KwxK3CK21hTTTIE2+w2Gnr0JlWCDO8P2k1MagTUrBf5JMvHo1xOqnE/tZ74PBU6ZpFxyu
fUQj60WEkBaI/je47goSzlvPb1QBxgBK4MOE9JYcR2X7/+37fsvEC/7BvJ1KXr/GROrmP+zZNtGP
g1qEYbdf7bMuOegOyzogN0PzT052CFkeGY2IdBpAsGpA63kKz+u3j1Bgap2mDimdXA6YR48fYJEk
X3aEmysqRJf8HQgZecbb8xemQwIZSP8LqHS1QrEJTvkz1jDszKZysAZyU9G4pL3Ru8mRz1pFNM01
4Fc3u92FmpGVg1/FyMR20DVR7zvPvcEDVIo+BP7KYSzl9BKumrysWnYAZknBmrMuBOKzcdOfvVm7
047c0I1BT0CYydB0Mtv/aJkNTzKiLvtOHYpAYhPcBGpnHakC1JLWFf69bSzKOVx4DfndN2+anjDH
pwdnI73CHEGODm/TmeID5j5jW6oPOgl0SPArgE/Y6s91JjeYk6g1UUQdo4iiNym/PTSUNZCfAwss
Bm0IkgfMdvRdbDq7DnvYBC8G2w1OdGwZOG6dWjwyO+DfyrJuN3VGtZYZNlbna/hyzZNL14KqKdAa
dsNDQY2qeu0U0jTeK6P+Qk7OJIKzspoFAGRoFOqGFXePoV3YEZmji7c6X8OIefR90kfipiZYUK0u
OcdxDKiXchlsc3yVClYVM9Wi6ZA7fOLKYYUCq+9lY6ttvJO0e5zCTp4pWr7xTz5sDWqlHT+xUC7E
pBTVm5YvhKwezbzBXbD3rXwI9b8HbKSYhf1YRgnVI+kBVsRwqQxBSor7Mn35NSC8jKwgm2Udr0TP
OwEDiCsYDQm1efSEqfwXZH8tXuTT9GkgDuMVUhDeDG+w270tg7u+jUNflAOS2dAg9mKR1+CwqInw
7aHC8RA6P7I/g5fMRXnR/ajo7jGVo3yNC14/RiKw81s/5gllmtOeTv8h5Ej0zaq9fK23CuVwLrbH
c7MxKpixtc0bNe2BDcL0p85vSQty6LXxTb4NCelO4KfYoYkdl+9L5hn0AYznuw680fVASB3/D23r
ObvpHlegI+7tiM3c6xkot36t+NvZk7xy/CRUAfEfHmdmzsgWO4O2fLfjbIpSXwX/wdPrgHWGhhk6
Kcf5N/4BPOILCei8lPwML/Uvx//XWfumFkech7KY8X009BAdGv4U9KzRCwiurvLkNEA1KE1pw0lZ
AD7toM0hBz1TAC4HX4tBaADx2crv0YUUIGUGI0QOwYGBfYgyB6V5haLfdCZBJpL7FzezpSd/lQ8b
hD+fxFN8vv1OO8b9PFzHIO7PMnfTSE6r7VR+s3J0dN+eo3E8nB2onSEoARUFpwHCCDsFlyPq9kgx
feyb3W+EfX4nmXdCkKuihMHepnVvQpCju485G7iPzCVsNY5zNuq6Zz/GNmHt8GTgBcZJX63mpHSJ
FRCMOtRAPyyzErOqqPFt7G3596Yk6hz21p+uRX+ygsI+RHrs7btZTriGjZvkqUBwOoizFZtA2wLG
dTdBI/X+iE/9KoUUwIqHk84rESkOCMptAcQmyYIu0NTyTisBKXqJBLj3xJ0ywThsaWs1U+06VCPg
NuLIYk2UEluA0zuriyq4xPnNPCTZNS7iF4P2mXk9Wyn9KYEAORz6+iquOaOeMuZ98qhRizgELA/7
wrPfkvDVoNm1nSENVj25AaKXwr1BIRjSsPXuKHpWDQ3tnPwvvS0Zog5HU2k0cl/hjUptSxqrNAC8
f0zq40CwyyfRgQgwbQ3HAhP6+++ufIC2dDNglfDBqdbxRnc9KrcQ2WudaYuST7/iE5T6aXGJY1nu
RvB3QScfyXVR592xLcwI2oxBGYeYLhcNoj0zxefT/QPW2wsoLbvoTAgJttfj48aaNesFOU4Uyj3C
94hGoT8JeiqPWfUNTmaq1Vu0lsMVP3C20fXyHLVYlA3IZO4oiNM6w/w3WK9mH9iCQKEthBzKwxbZ
UhMwdorvcp4M0QGTv4r9PTJXY3P7mv+LWeDOdI8W+LTUeE/o2l+w02pmWOCfz+UThz0S69tpUgvv
fzprt/klNOH9Ahxhx3pwFF9NAMMSlgL/jHKsOQspVIwoSFsHyBg0NcAQ+UR+90wtJINh4d0tKhEq
XXrnnrFiiNw2Y2Z94Hs45chlp1t/mq+x0IdnqSa9HA/vrzABXTp7mGUdHZy4TcnOhwat4AcfFupX
Dv1cM/GxFwHvwQcySLzIfeA2S7skzI/XOkTVZX9FuCxSfFqAQ0nbX2GxRylFafInxw3n7ADDAtiH
XT50D03CyqCA3rPQC2hsOWdbIdi8wSmsLnvsliSH03/n6OPT5aqphwE7fzZLPaC7ZeWWcX8Wr7rl
DJHk/SmofBN0zdi8qPJ0i0SMvT+GNT/Wjaclj4KwBkHZXDK12Rx2PoMShJ7BoLh/kKmyyXYz8Uz7
Y69tDAKfEvmko7cZLeJ1Td1mTbThBr87n2V9rk5VgabGNwXtmuatssrgcXTI2KPzI6nxHq4jEJV8
vWbYBZofvTvSAn9rLEcNhkzjQP3laeMXCC/vjSJly2z9/fIP23SKvWyO4xmxA3m+cwOkQgyriymI
eJ9tmQSCk/QhRHWf8K63HVP16WXwHe613NHtN9qwhEUWDKiEcHmacCJ4fi6AS5GmYj/J8/CKGtTo
2gO/H1P4Mf64u7WAcD0nsgPaC1lpk8AtRbr0PX4LOxyNQTrx8STKut/TrdlMCBwozMJUFWf6pqd+
0nDHRPq7+kyBJEpqGobnyi1radMx2B2Mmg1S9VehJUHWsJ/sqZJEYrpXP5FGnTslSUniMdiqgPNX
2EFbGQRHYnfw7CS1OUOx8nSfZI/UhuTD7zWLWamSXtUO7jTmOIpRiFIdkgX2Ly+o3fbL0frZu00U
vRP2G+9qhDiURtE5oYGSDnVv4uGGAcK0nMN4cCxaAWkl7xCxdDshBAJ6ic3dis5u6OK5MsL5mvBV
JtUzB70OVq2oqPfmSHgfnc6gg/y2DZsjP/pnOLFZeSdjZ3fPeJ6z342iaKQMV2s/7PyC950nb8QV
GRetsA6s3OK49CYG2BmrCnir6++ZeS4K3o1K4CJWp/Wp1EhhhuU9KU/FJA2F/Rq8A6ysD1QoRs9B
AVGWwyzKBF87DyX/rSBX6svhO3cvfMDRvF41GZdgvfblqqyqgYOXc+O2by4mgwmjkr1UJjLSoLFM
wJlzAf5CzK4brjRh+3jZigWH0Ei6tmBxveP+06XaRctdcNR3FiJHMfCyHprdD8poNILsGlGMggcZ
9GflI/6WD6IuKfk9WPWGOqmSVsGqMYDa75Mb0oWI0wSTLfS5T+sjP02B1NjHVUv0ocheFK9UNqDw
qWaln3Zps9VvlBDsRb8PTVhRqBoacLEekJcKOWSQqrGU/51lzjrgt/KB/k9iiLnX1amQ4LTs5e7g
RrmmH9PWcFSJhiXkDEf6hL8Rn2oyRgAXynxJ4DmzkQ4tSbwnAw+MoQWiKa4DbSlioaiX5eq2rax7
fjw6FF5kZc9d6J/11Wn42RX+Hh7NWmbyi+hff5U2damkEzVgRbZyeL4QVC1/fyAOQ66PT33zryMV
WeSynpx53JgczDCA1hR+jy+jHG5RS3kEjh8LDFa7TuEZ3e4WUDSwyOapQ35bedfBeSqYz3knC87t
fCcFCfn34hfVkKIGuPknojM4Nu5i4bxLWoTuir9Thk5Sz4DiezOgE+w4Fs/bq1El0jvZfpo/3vxt
O/arPAgAsO8WTpwFVwsnBQNI0WumYm7oD5tbOs3by61zxIUxq80frKsJFJd7MSKr+eqq2kEw1BkL
rEqo3psNV0gCuhCMfHSSx4Iv1Z45Ys0bQ2MBkR05Z0ckyTnU5kMAkIQiUc0f9UAGUUW1XVhvDpET
oZ1t22DEqBw3lEaXdys6d7HJg7EGDa6m0uL11wbtN/4xJKsdHX6s90QtYjRrGzvTeo2yu+aZh6NQ
2aoHc5s+edzbmMX4Vv+l3hChqmurDvBwToF1V4f0zdDELH7GU60O1wRL4R5wjeX6YKZO85u/EX3g
efRbPvk2wFNdUw/vkOBMgYtfUccR+Ed+F7eNKeGenktec3v6PfhlACJ2ZOvXOOWYGRabFWGR/PAo
nUT9A+5hky2pGDcDXbGppVMfMtbrSVYHdqjfyYA3k1lQkS0+LifErCley5a5Dthhhh2mIAjaEb77
oFGyVaLCcM4vO16v8YJHwoKUdmyeyDaehaSU+vUS/xxB8h5+246FtIgsQdC1TIBP+0DmVyJVi5BE
xYh5m7Sle2mHcVOkRgel8Y4eF3qrMg+jT6HPlHtW+fbPq3E7HE9+SQqnRczZZifT5s6CV/GttdQu
oFa9VWZlK+u/4QrlLTlJT5fhlvJVMLhgNkZArK2vpiZTa9qF3jBW8qIyndzrPBxX1+oa71udzAS2
v34gtcZ3yYEcV5iZQfBIO+LA1Vmct1Q+YFlmIF+8ylLy+ylh3C207/R76zbpucHj9hYu3q2AzO7D
rPt4WY/HRhfSOikhQR8cHQ4YyvNaG62vOLI3ruUKhbN/hxT2QmQ/ihLFLdIqnBFiJU4ccrrebZLx
bZ3W7NAEj+btyp3b8ZJDRS4vnNUn860ah0rxLZuN0Brno1txBShks0RUvzsrtn8gydA6t5oKbHoO
xjk09jQzskOUgz4WspBt1QHpqsGJdsosc2FwqyVJy3DLza8AKLOoAZbHWsRuyRZ7JQJaV2EU9dgE
bbQ6N0hqM8rv2qHUP+XDwPAdtp93R5x0KPauJWgwwZuISL2S4EFqRQn++HuEUlCdZuSt0DmYXic7
jI45KTo5Zp70EiNVlc2kdLKmjRGhEgjDNHpH3dhpX0wI/TJ1lFdIw9Zt1HI4MMf8oMychAXtTNko
3ROSP2gmKaRl5jWWSyb7/P3Bw1YU9uwYUmulsuCXlRq/2Q2DST5N1lfpIETtfwe2ixuknYgxxdHI
4dh6BHfzFunNOJDeHwm1jWaUohkU2V0ic1w1SkUnpGg5akqCUXN6cqOtkz2eWkreaTYOxQ1U/cQ6
Zsb1xZ/4RzVGXOj8kodDPEeM7SNPBJClfiKSvJWY+eWIPV0hiYW54TwLE90PLzTyinz2DAxgP4us
nA1wr1quEzlldQXL8m5QO9oaLZEbAUOaCZCcXjbiYoKtc1srhJ7BCa0Qd5C8haHmMOQTSm3eqSuF
iRqYQ82TVOlHgv5y01EtYX31bHjknJaDzJosQGhTHdzcxE2goJOIpz7XVhFrOCSvU9Eg25vEKMV2
2JyYflcajLHA78fl043m7E9+meFjCI4bDvq7OWb4Mnb1qhwQh8L1BR95bbz/z66bXGZ5ho9ekuaC
PTKqiT9NHe5tDLFwIbnPjWS/JtzP23PMTNpNRZXW5YUiaUUUJ3dtqVF9TGOFS0M7r8FoAnF2Iy1J
yGZKyH/ci8l5eBU0n3FWgi9HubFjRoh+EWwhz5ZwywUofWjpzvxRnzMLHDhSw98gl3zBfUi37BVc
xP0XdkPEQtGWrHy921DXl4lvmwyNqNmnO9HzSjDlgB1Vxj1N5YuLdQ74cLtEQLy9/BcAcgAyB1Vd
TraG71+xYdebkWCK2KUqOXe6BIydiJLrujEUfjSvQxLi6csuMMTUdK/OD/Y5jCFzH6pcmspMPVEA
ec8qgmYz8TyIb88VdFvfdB/634QNKJutmbUeG6023BQIs3KxeDfRjYosqxuu1ZA4WwX9a3rU3MBk
Sgu/dkxNK7EJYk0d0NIKFUfT8nNaqV/sG9l1BIVA6qmHGv0tWQVV/qH0c+eYEEQrynENMXxpawFR
bu+Y8IKp4JsbhbtzBZaddL64K5QpHLU5NhBXgG4VXVZQwr3XT5QH6FcpRRvJhyRnfN2y7O1eYC0a
9s6rESkYeI9gQZE3k1AQW5KcLrk3cCkPx1TS8NGgbXX6yaqmYTBUC5dB7gJ+/CWZNzm7JPsghmXh
I/cGqbYAg7hAWRRcHak9qgoWBQ2k4XVMULIQZL/v6zOzdZsDQ4qwMoc01wKM3t0FeftiwMQnZsYj
OruCfi/eV3r4+KoYO+i5Ukxt0Uy+v1baxNltf+QFLW9ys+IrUJ1S20OT+OPtJOQpdSGASNTFIy7L
26FRQpqEraJKHBe2/NfbiT4RDWc0nm400FKez/XYY1KOYBCZj3RBjApO7/W95oOuHzhEMbFneuEZ
YcXvhVy9fjFhMbmnsfyWLlFZl63HzAUveM5ctALH91Gsx5xatmbZLD3Z2mLJWrMe4wW2nJUbSnwV
I/K+utm6M5u3GkgAwym1BTfafp+IRvGzYhbzc2/4J3uLNWqbmHKQ5kZURVie+iCRGJXv5oZZjWih
+TQyJnLvEAszIlbC3tqT2MY73aIg0pvfIr/ZJem7nTYdTGtvyXIEF9YRyLkY0zIp4szQPPezovoA
Nli40CfIVomiY83tCwhFJ8Mt0wcuW/RVc0vCkLimnpAyeGngqX+Idh8Clet3RwLe5HbOcaz1fyb5
Y7CgUvryS9SX393O07fRrI1zvOZnDMxFYVl5MKoCV/9SJKMd8ScPZnGDbXfurTD2zdCzZnueb+d1
TNFvJctOZMVbqvKXXPEXlCkEf3C8ahwoqiXGPN4JXmH8/pN7/nXNWhT0YAGnNqt7n+n4ZAp0B534
WaZ2TdmRyRX49GLCyzi1F6lOg2oKiDmLm+Jrev8b8tqXMeZP4pXUyX9S528BkCiMU7MYx30nJu8w
BAl1WmxCflGGqMflJxQ3F8iREGWuacV/D8SK2GwSPXugZuYhXCbZVcGFh7Frhh3v4vVcQBx06VHB
9hJcRSeHmiJ4l46MZnWvhj/tZ/SgUPA3M2kBCdlmGMbEWLdXAlWJvuGNx04WPMeMvwa6qxILIFCE
wC186p57GXbXKDTga8esQrk00TJcqsF+zBHco1pU4UkalZXgqw33yur6x2el0V0jDnDMrsoAY/3T
KiYpu5iIGKCj/TUN5sZIK0GCioVmk6PcgrWuNg9o0VEwQVr1zQ7MKLCofLZsE8g+5+FAdxbmNZGl
q6K4Oiv47u3TER0E2BFQHH5pwE96ugZn1dihjo+hZ411Eod60wGk5dPVOpHjNzosn2GChnhukZuP
HmRy0yqwMKepQQK8a3jYuxF54pm+kkjbmS1drD0joDxN55Lowftjwu9ClmZF45ThnvGRQBMbXo+z
COI6Sci6KFTR4tEyVPLgaUE3bPewVU1m+tD5hHsgZVe1TLyjI+be7nJWa4aSsZ46goLG96MetE83
OLXGwb/To5HYjDGkJwmnK0R70yv79RFdWaOl61t+93pRikeIM3lMoruhD55cPFUSrkCuaG3IzC4C
kzHRbVP6QlWN5oBgy1/3q4598XtozYckBmXMkQcgBCwHS8+lQZZfjNjfF5Rd8Kq8hP2A2mwT+qsB
kDfm9vF3wntzCYQjCOGDtRqQL3rI9G6Z/CMxl0DmVoPzh0UphfG+tfUwDo3YQSGAqzf+OWcs6kbw
wXHUCjH/iYh2vPUElh0LoS919PJPoC8HmrP8v4axn6AcnTYOEi3H6H82/fo4Zz1xS1uuNGG0ubi0
WsmaUGaCbFI6yxYWoYNOC768Su6h71lmX9dJvUOYBcrRce99eQ4o8iFc6naz0n8TecnFPAM5BNBy
sVtAoJEXVluSk4pSXxz96zGo154qDLg/rtnD20dQPqQh2nt6hRY+HxuJH5NxnTmHMYCjoCK6cKmx
crID0qGr4desJBG4NJjOAs5S/UXQHeKMpLZCA7JZ3uTsKPfwKayM3nDg1pT1yMxHlVK9Kfww7zq0
otW7jn9+aYhC94LTE4AEm3Ha9dC8w8qFW8rnaShnpm/5Emv1MwLR1rGCSKm8g3N/8Jz8x/inJzud
MZKwHVO7Bq55/S6gG3OTvj8GZXmzyDuixqV90/7YX8aPUIllV49OQuI2L1g2C6GlBCgcavtznJK9
u0RD2EBdrCO8L0pOAwxGW1v1jFeCGh41GloOBJhgAcvw7yf7Yf6Vc4r+kIlh1ZIc9LRE+7v4M3oU
Lp+DHShsX6aAQvJdnNXxo8dxhjZVQLKXKDsEEvNeT5uT6o+slChj1tPHBItNhMQ/0qoNQ/VAbXxT
0NQ8M6PK80ZwpeKqKpSjm4+ykyJzqymQyWCr/kjuesFp7NtuvQ76x6eC1jIRvafRHHhVPzfbeJd8
9jvVm4M3JK235HgRkWL9cuKEtu5X4eGCH5rD2W1BKBKgOw17iZ0w8WWEQ2V65Kel4piAWrjoO3Oh
6/2QfB0fBMIltnBmvsP+Cluz5BfDQpHV6a0qgcQEB0S39GGYiPptO/1HH3WFTgBOuMVnj8zHFare
1qQW7dailUen0AvNwBoLju1mMI/Ru0sT0mOd2fb9FWAe4snQZqBABqfl6tRMdgwR/n0Vu4Xi6JVo
3/wgskCcem1j5k3muOlNKSefhEGNY7zE58njgfWtJjyHze8GS56ne5CbwmxoITeyCknyssAkw7EB
0y6zJfJnMtj4x9tT25A4tC1IlAtfToskgp/1Iuk/Rt6WI1rk8CKR/EJenz+WqxkarvMEA4OpB7PR
g3vSa0yDOZGEO/jwHzbX0Gq44n4IMZc/zTxKMCpxy+5oqzjjpG2u2JBJpnxgDwbGnLDj8TdOIPtX
X+T3w/jUaHWzCPwDIwWOy442/ktzSRymfoIC0158xMGlItSzbEL7LtRf9qZJw5GV9Utb+nQkDB/z
moldOscXjmz88YCxKOj0USwq6plUVmOpKb0/W1GobFcykDEJdS0tCndB8jua9NtjVxQdTJWfpnr0
ntI5rsr1ZmK5nZH2Wm4+J7nmydMh/y5dHoKxJJni+wOizqaH0dLvoBs1vJkIndNkbgnqgiMD0EDC
0iE/967hHIT+VIxYFH7qnex7+wRO7TDE8XnCFJDXMo0kEQ7V0s0dI8NugklaXLWVjgru6IS9cqUl
is3pLZTFVyfmqFjHMfMhafdT9rcdpt4SP2PwYiMIiSuimzFcfZnWchvLBAkdlzSJnlDb4h1k18t8
iF4f3xxXn4zZIdPD+xXueBiCdsO8iji3zhkcBZ/qgUoU4VciDSUTAkJZS6TvZAtn4gADFqZZ2/rS
F3pA3gRCzF/g64jeuyE7yAbiT27cAUdtiyXQXB/MliIp3S7ibmNVVhUSpwWityH7XMj7VA0RdzkB
8y9RPwZ2N4if2hLjhmk15WKkVuQtNwpOzQzs7NUOLPL05/0FI8FaZphE4iygt0SgLLnksAJ3zizs
pokm9dsRymKMQWUnFDeU1oHKCIaqY3vj0qUSeOEJCdivHMBtU8PYD3zbUZOEcMY0FYrXVvRXvala
c0KXH58ZMoZufYU8Ad81W0Rp+1Rtg2XRyPEE00eY8NwpLRYRKEcmMw3NFlue/S0YZgf44z5Rss7h
99t6jonTAewGD13T9O2m5UpqWxDslHVROIr13qI4W7qFTvWjc97Upu4pBkHJKJGI4r2q/QwstxIX
tWHVlc6aMCoPxRJWQlQE37D9A/CZEE4KRGyJki3xKjuFlCo8OpvA93LkZ5ZLvROWOKGIZ+8Pa7gW
T3ndk8ht/Uf8+jO7YjsLPm+aJfaFjolwWocjYBiF8JvHe0sKlNUmCPH+zuUiujR9Xb963IbG4vRq
ldHFMHhGB4gBXwgL0diQiY2+IEPGD4AE6aI/aBNmSEdarV7+tujc4o6882jAEylJ3BJD8RRtpsqc
ishjwwFA1rR5hLtNeffUol/tm+aPq7Rt4b7lZFqDACEP/MoPpbcO2E9wu6OHBMXea1YUkexiCnDw
lYND8njY1TAcuDq4P4Q4c1i2SxucBGC+vW2zpCjWgAjEz2D9UJmlI0BEn6DdZDZvEHmJqDPslgAY
HdxRDnMNwYsYnlufPdt8cNVsObBpF6wpNm9tGGfHm5Jxp1zmmAK6u5ToAqda4giLrYk3LQYy+kfD
yEX+GhiBxayt4xVk5vfzitmx/GfxPnmQmSXzRyo71dl5ahdlKZo+uIlixXeX8hyjNDwzq/4Fu2Eg
2Jakxfpbr28v/U3nwToQmnkPlITQyf4nZ/ec6ikw0Bbb7YJ8SAXKoDD/04K34BjiC8MlGBUuirkr
YRSha31K/+WZQHxK24XZl472B1l3zQtPYNkrQbTJPvNzO1G8NQoih8LYFOZqm/CRy6p9XGckfNU4
2K9KgN+lB2berKmb2vNhhlgYM23IJyvW6TulUehOfUksPvP+YHR0UPJz9ZZYWhbcLqXD3vuebU2s
BXNbuRTPJ/euvk9IPhT8u3o0SSFWfJvHlDUoHEiip4N6q1JIKzLlF50G7vzl6QRaj/H1PK3dJDjq
R8/aFIjy661RQc+y+Rh64HqwEWfo2/kRYfqu6gRnvcaqw1s0jD+JQFtVszVmdZUNHaLobCv+35Cn
sFWol56PjPiRQSvMSftILlsTb+l7w3VAxO0acNX2MBW845ntSBJ+K/OfG7YW4syYWzejR132worO
xdmW/diu9S6GmrBwzh0IJCHma50tVBu4tum4Q5TrwSLVk3cU7XK4cQjnHOCnDlnZCJRiORBGQq5n
4VgmaL8biioIv1SITY4RNbQK21cuULvTKXl4M15QDcX2aS3jgcR1YelQntu1f9N0duTontALyd77
r2iw/Ph1eiNbukcZ3NY1hjgM+NZbxRXKPRaXTXXV2Tgzxl+ygk9s7lRDQR6UScUzagC/CKbIOngN
rjbPNWJ1NQWSVOTraFJaiIT8/kiD+FSSAQWBUrlz08Uw1ORuQhUSF+jmzsa1J0PohBvDAYns5HHM
YbaXq475WgK1lvuJ2N8PdW+GO6Jf9B2VHeQMKMqF8oJjm7Mno5MveFrH19BizLvSg8qOiESUiwwQ
fW/r7aqNbU1OVHdgYc7HvnSz76K0yrNwIdsGzfxq3S4ocVYTiWMCTVTis15dHn9qxH+b1d9EPCTx
yNI2mOxe50tBVQ3i5UjTfnGsHmh9pHwzMyay5vFe2Hoy94zvoZsSCtEUebNAUtCAXnNfQRHl/oe5
cD+WCuIgk8oVSJ53uzVLrK9vJzZxdL5GEV6NNutn3gYUreEBt5JQr0uJKt3IoONEih7yg8jHYztj
Lzg+EH7L0rvmFRqLlW0edFc40Av+z7ipNaQEC0Ko7yTedM+6S0ZkGD70gM/59K1mXvGbsZ7KdF5W
A+e00sd7fDXLQr/hHgrWvQljGwhctMRWYuIsuEs1xzpGXm9RWYhlJsfp/kTNdEm7xPpYLT6NkscH
NsMlZ0MIMr8xcIQfudOWmjAjivqjmiB16JrZTI92EPOi1kTtYH7W0CfzWcCOk3lmqefc0jrl6k1f
HAI8iQHaOQeN2OPc04JK6EeAoL3NhxXd/w1oGpqrfJmx0Hh6Yr0omW2sEjt8oxxihQN/MaY9QmPb
F1bUCqYeX5RVsfI4rnlqGQ/tWwRtJgg0SdJu5Ptk4BdT2hLsR0N/Jf6qLfYEOlPf5+MfGV8/MPlw
El3msteYKN2wnp/i3GGgtNM5R7Q8NF193qDNvNrXZyuqnksRYS1z1hBKzsjIE4QdERwE8yRc6DkY
Dt/ADmWPqFAwBkUpCiwIjnyBrNX6uyn7mW7kAKZlLruRJ2DNTKpRUgFr+25k4kYrJHwIzowZ6bYX
RgkrJKePVJrVcI3xE5IU0mWXbPjzmCtP3KMrdm2ukwVwvzEcWHPJX+npegIo0gegnJuY36Epq9Pg
g1zAnRkGhQJ0U6ycb8Wh2jUiG0HeT0jqYwCuM/u8CY/xIeL8L6eLnGCa2s9qJDII+dxGeVPjGXlr
fdkwKXt8sWsbAlQhnqGE9NNceUM1lKYaI0rg6r37mpqSZ7gJK9Xu5cUI5QD8HeySX52+t5rDwoZZ
QKS7UgS26WTBBV9nEmff5rrAMdaN3Yi+42A+npsEXMZcK1XL/AZqQJ9AUmhjHibD7/T5YsHSrGKM
+jPMvg4FtSHI+OfW0GSVsIvzJ9QdMimsW+CaffyJUsnumWUMr5UhVF5Ztq//0uxcEE1IWVnfQ38g
Ui2UbQ5x2lNjnlBSuKjdS4JhxB57Eizbot8YtTlI0ROgkVTmww08Ytn4O8ZrTPLk56JH04k7R+mx
fURK79gXvwc6eMQ3EAuCARCap/d6wh4uieQVJY0mb4xiPwTnYp415Fk9WppWHeUZZ6viy7zp9Tsp
oe4IctvU9tLOpk5xv2aI9/UoSC0wGzxkpjMl6wOQsKpddxYEARDhjRghqQu+r2P0yvSPaBeacfQF
Jl0snYi5GQhpV+Z1+SA6L/3Rw1cZY1WHHSUjooCuHCHYxfKkc/+UM1mnl3quRICN95+akRTOG0ZT
IkGBoq68WUSTpTyC3DRA3XWvGtH2kJHxISutJ4vlco0E5UK/drJMHHED/UyhtyAN5lmxvAVsxvc/
safsyoVZNKlXavGNUF+p8z4jqrObssiqN+zo0X5P9UEQQ6CHJi7Z1dCYGfpsQawoPy2oHpvtV7Gg
YQli8BNTCxcTkLJqgqFgrGbAc7eQzQDJuzY0cxWR1jbaHTkzD/a29gkhcJ1bdFhHf/PKAh7d1dY6
0nltvh+2OGG3dmCFb0FEBQ25KMYV1hlG/fTpwr7vnxdeo2eIV71+eQBOGGgiTx3iSAMloCXh6N/G
SkJmOEiUTWTQnkG2JYV799a6F/EibVjGvXuregO6JpWS7AOz/H+Zw94OhG4Phj77a1S9bbeErmVQ
3xNPBqa4zD72n2XN2SgIOF3pWf2xKkIBp2vgmgKDVco3sL1ipqySJGgsD84zuxCAyOBP6BjmqQVN
tmHuu/Au8kAENVLT8jtbCmkD7YpCHrnTcUsNKzGrOrkrGtBp75i9eg29mdJUSwMW3VsA7OIzmblr
0rWhR1XB4fggCYwsRRj4fLLoD57zu8ojPCY6sGkR8vtXJJKxXF247FbLc0kRbJKudCpMOz1vgiSp
p+MTiFAutgVn2Dwzx7VbNR8IuUKDYHO+al38jlE6AiD7LIOUcRyMXMiTwgiyubu1tdqXOYlxxTo6
ZvX/0WAomfu7NFRjkBTEjWhnX1jqTyK/0aj4vG6sMFEvYYItyfL0XQFDUd62HIL6hbgRZ1MhKZqd
e815kSF+mSRXj2FVY4YbBATo/rx8sAA0S0wicMwYlC4+t4yXGDV8BPf3Stl3ifqvFl3yGgY34mwv
p0ye/tseFx5m+oq5FWj+W5H4VY95aLU4OkVlHCThQL7iZ4kfLc+yGuwi5QnNbh9fpYnN8DDRjWk4
83NfVgSCsX6rHglf6oFhef5WupHiZc5ts3tDTQeOSiFOibehXyUDjK/m6KoVV6f9wraz/DPWu6A6
2ZYfrXavsrFD2R6JYCcOiJsEuK+TJXi01G+rxo3JSBysoWzTR+ujek4ROMK9nFrVFyFtvi8PIyGG
XK+F1OeOeBwxz/+6YCMO/1iTDPgoELjUugNVoVXo+Mads9hsUcisRevWALPwxhD76TPR51rqdDp/
zxEqEG9QoVrMWOUUdB3x3TuM41FiYV2t13U7da50K/QD5agWhuLIbvUVOcBT8jddMdimb5iz8Axr
pjtmc8IkKSU89kKWRf8p5WcEAUHyI3xPsEejriWkdCN8lBwqo5KjIx3+dgYJ0Iwy8U4XTPOA3DuB
7S0G8SpqYNh022biCsdwKiOrLMuh6YnJQnH+MCHuUfAY3VTZrDL1OdFxt44+E+rDjsLQuLDrxsVp
5EEakvsY9HjiahHw/kp8bWdZbd77YHAhlu4FcuszEsM1KnmRrv7Td66F430TFYXA4oG3KuVIgm6v
XQqJWeDnDpuqO/fPG//9lLFMglhKZyYi8wBC8fAgyXbeKPCO2GUR9Zs1yDx91yIvhg+0fMKq861V
hc5VHFrQOaT/wDkmcySOTQGVdUx6zZXbQLoyV4dbLu6cmK2WmBwi55c+RPRzWooRFuxhsWSp6QAn
t5DDemSdJ0+sUJOv/gM4BZgDTEDgekXMFP60/11eQ22vGHnG2/WhRnCTLkd6hFiE/zLXMkd7HzWT
hETh9/bGX/+UUeZ8mKNhceOHywaaw/fU3/VFpYtcb2Dhz4HEPRnaTUeCjChV+de3pGWPL21y1SNZ
wjPy63qv+SkU6aTi0L2LwXmXJKdLckYekR0xNL+xBPZWfcbYKxRlM2hq8EeyWoAcVaQMJUtuYBlv
FYrMMminAfSiE1I3iP1ckMvIgv0nEphTzdncjCzT7kX8QcoO34sClsFPGoYJyuS0HGdGAyLEujZ0
3blpTGA66xCY5cAQlFREpAK/sFDY1+Mkncsz2XzCpsS6Pl0xcBljs7u1D9KURvQbLNyHBgFjAd8B
1PQObT1ej7T6Eg/FGtXIeMDV8BPl0iufyVE9EkX+Fu+lKndvc3jFX4RsDKbH+1bkcnauEzbt22nn
6sTUHg6/FoUJ2cCkLYAyDDi5eAnZ7755D/VVpCZ/iConC0HYXtShIRTVwUdDhKLnT0tEn8FlbQNI
ACchgwDEfmfFtvSdAHPYTL66wznktj+ln4acrRRSoS8+rtled3/QH03X/UB4Z0m4iZRNa/PsV+WS
qSLEHIW7ytU7JfTW8azvF32pR9hyaMxc6et1MgAfq21eD+ihrFJz4DbOblySRIxaZZ5aUX+sQg2K
yDQNmqLRe9RmuDToyP1oG/6kuu4Xi11ae1xKU8WrduhNHKTIGakQwr5g8vYs/9arvhlE65rb5G5n
czmlunVuhU4mQMOe0VsCCt/3+BAuC8yUMjaZ8VTsXpnKc0jEG4PN628EJ33q4san/uk9Z1gnMkrp
E1WA/kSw0ncNAbiEwzZ62xIEsLOdBKM5EZ9lEG5STaDSnylt9+T2YWhNWpxHC3RDa2yM465Uz6je
N4UENLa4fo2fpX30S4XlcyqVfqql9GmFAm4xUv6aUfhrZMtSL9sqtth/noKgsGZAqYENBQZt3WFa
U0NwSBbj9ukS0ZtBflFu0MHcjkxtnlt0Vj24GzaWoCBMGNZ7YX7jwbN1Bb0Hv3wxlt+9q4G5mWOz
/8kNHJQiNJBpjP5XoWAzU29Yn7OPJ+Gx8HF7hOxWIPdGWQpaGhq1RZUiST00TDtg3xFVvmWTGEP8
JhQIjobDX3NsRhYAIMEzMMCVODquO39QWMMtZ5fMjGzH6m0dKIMmkA2N9CwIC3Q3at3XcUPHOIeo
hKyLBhvfWrwAwtfvvGk499N+OSY/y3hzQq2K3qcmXQuX4Ylz3kYVTXtdPmbR05StFG2sMAo6mTSm
mTN0jelgqgFt8fbg0K7u3hJ8cr77YDAmxG1DMD7V2m9z2Ctkpndjvw5QXPdRVSBPoUgnAqLwqc1p
83JkoSyC/WJeqFLzhAZwlbvvFz8P1hRbwiexnCnkh0ch67W6urlsrY34t4og6o9gn0TvfudirNqy
vr3m/FmNjy1YMmQE7MFRDRXTEYpvIX/cqCOIsqAb/U2o6u31h3f8XNL0I+lDDRt2zgiCBdbhVyzu
ffuWn8JhYnajr6VW1tBEsV01XJh5+oUgI08RA6fr5pWwsMUgH6NfmfqZiO2d1RCLzOXGRNxbwgj3
PtjuhpiL47VV3ryl4CgNUKHJlxg2fxt2UjJKe8dppLtSee0EKBdl5dQ90okvbQ/516tOR04McSev
SByfrrJb5Jc4Vt7e/6zt315OBpewLWn2EWS1RYPS41MxHubJeywW6mD4T8QdM2hX6Iqg1N1cSuF1
J7sWe+Quf4DYtU2O//01f9E7l1K1hh3G0HWnVbkMDT53bdT74XkqSzdpKC0tPzKbyTvKgVDxFpNE
eUPD1gIaQJOi79MGfdfk9nvuVISSQdSJciFGi8TE7cljPMPoT9RbgTML5849KUv5VoRywU8Y9Dat
/rTFAGoG8/rnivxAUCFtvAKHIGsWVFZt8nY66OItI33mZ74QDxLZgyMysccNJhEVgH7nqnbenxQr
9sELtzIXhMPh13iGJhzjH2wigDELaei2ZxBvEZgKk8fIkKZvTGEjynKpGdtHYRX9R33Lsoh7EMqA
GIbiMPO7MhhVSm+0GrKcUCoq2Jn+E8C83uKgeYlzlR7Fe0cykh6TD5ZQvvDhUf5hZzo+GHXjEY3S
kiuq4lOv89aX0bthWh50mNf4VHx3MpuZi4u3/ASI4QFtUDSs5L+NM3QgJf0Pkszo10amNAhIop5K
cb1sElk8PbHyWCrYS8ofoYLuMlddwGif0kKt3oHeibDYmh861MHQxoEUJxv+cVYiRx4Ps0mKrD4+
fMF/gLwE2Js8F38TEkWkptn7K1470XsZDmkQkpABhNV1R0VZRUJxCyGTSLSQjVcprp4/+cwSBHg9
PGL5dbo+MhoIsffZihVUdppQe0gkmYfvIWebLNa/KrIIvKtYY89ZJr+iafbGQv0Rcf0A6bxZWJKP
5bsJmexhl4Vphy1N5sX2FPjSSy9b/94u6tOx5ziT5eiCVT+RuK/UEgSyLlG2llikpdrQsJCsxIFk
kJv8pdUJ1/E2XUs79BZMYVqyKs6Vo44scO+ONkcNqMowk7Ib8PnujxAFa4Qn1SjSjqOldDC8k2uj
7wIgaEakMk8w/pgrwEJxfDR85MJ95208siWiQdununawyXO8PXImhsPdqo7l06lMkjO4A6Gw5/Zn
/b4rpsJRurnmrAwsCKV1yzObJdTgu5vQJidI5gDs3aP1aeMJnk3pUA+WEK7QDzg6ZBAU6L0z6t49
bVCge4RvB+T07J3uCbT9JPiQhPb8EcqcC9uo0oBUJRbBDxaFRDt3JyTAlYJ3jqHFMm8qjn155MPc
vsmKZ+sk7kNKinqVLkpR+FL4ZEKWqFd9reFcVDDpDUP76SHY2Q/cdpdQ+pUygWTyyvSbGzfdDnGO
RqtR2JXMLh9F9IGkmKghCB7iVNwqo0rXtuRT+k6w3L42jXtWhbC/dkMFrKlRkXsQ5vHZeX7oD501
NrJEw8XYgdwzpHjRALFhrE0396KPnA+s7EWE1FckpAmRmbzpqMbv2gt9/qfhjWGJ6esh6cxou+iV
eiUMOGaBhojPJLm5FauM0QoPbUrsK/QOl3CEt/Uvl8eGNSbmZE6De+XBRXbzXw3EUZQdQ+Sh5Ies
ndZj0u7KM8FXlWIUFQTgB969MPhk9XXFec906e6NhHn7fWet/fdAeBF5Mhie5WRbbUS4e6PaLYBu
W4u5VZ995pMBQz7Vp/IhoFZz2TRg6e5V/bFzlepCRwSLDyT0Fh/g/5Hz0zIfKLun8AU7VqR/Hd+d
Or/hYruySh+iK5dZ9GVqdwFZGme2s4FJ0hXMb5t+nFyvAGIWbNf8c1kaPwDhz/9R9+hpd/o//8uw
7yYQBTxxDtQLrc07bYUJtKMZOq5tgoPQDrBnfRyc2AhaxwvKC4oDfLujLoul1PeWFvW2GO1HI2kV
1v/SvpJuI3Y/Ab5txzq9/dVei3+8m9V/NQRu2WAATvgFpWn92RlPDKS+vbm4tu2dQEZbCr0X+hvq
MDZQT4WSom+VO+K4Wp621hI8zcERL8dDwKzylTOm0l08Vl3xDOWksBjszHKSnJ86nQdB8iad3UYv
VkwPChapnCV3BRr+vZoLLHToBNORNrh0EWtz+2vtV76nk715WRqmvNal15jUK0amAmeAWrQqlYO+
qGyQdPVlT5t9CTDn1ZfXI+F+49FhjXzAMfH1r7TEzcu+koNE4v98DFOnL9LkCFBAD7QOfvPBboVM
qrBDFSlGFsX82JM5Gc6BwQTqtHjgCE5dUMibxaWSajdFrXEX4xTm0UQnzWcUPCQWHKYwAIzFWpTW
uM5i9WRedMIR4ezq0bwIBnehM+mMKCEEvP/CZ0pFnLGq0UhWr79s2LzpeIGcasdF8PFXmDztY2fP
eN2XHpHcWIsxJCy6QkMGXmeghkKzCSsYL4bUh0uk0Gf8FQ5SMqpiG+/PQdglg3yWRZHu4pTGMLZA
JmXnjoTqlaW0tgrb4/JosErIpK/E8fPVmnNEhYbSisjxT/GRCH7Yn2MW8b1UFHw/KW3xuqc/Thye
OvVoCWdxl3HrWS7Prl368QLg2lRYIr+cxliEV8CpJNX+wO8N+QVPN+JTImMlmgCQtR8LeGgfM1p0
tESlU1eTe5y5fTH9lB6GGDn69PgMR22Ls01kTfX2GyP6AYd79X654FWbNREITwK/fMK/GgBprcg2
jnxmgY1d3hw31Q9MNqF2NkwsZIDhQ+X5Vjcj0kQiC+eGfhHbxYuGECKUE/5oQIPI4Fj8Lg5CO2rs
SYIl9MBdBq+n8kQGhKbIWSvfaZv65Bqot/0ko9JS5PXzQPqZnsPG5dKBUnLEELBbfbem6JmaudIq
otkBnVKgpmJw1GRjJy9u+YJhK6AO29EGk6tCSK+Jw1oAFjGj24KPbxhuftzDLmHIF3Dpm0YOJ2br
e1hFm0N7eUy4Jg2u8vwcNVLIyB/j33CAqfOj33auSo/yZmr6G+BWy5vzE+S+NyixQy1zgRNZvdJV
iURH9wrTGrVDMyxoTsABGBm+aH5QkH+rdAWiHSTEwsQYnMSbWqKUdrQ3TDsiiZRvuSyPF3MK8+1n
elWirKRBdPhPtaKHuPzuLrGoOJBSaxUv+p6MGda6axKuZy22xYKLpLy9wlJxSwxUaHOSaXytenRW
Cj/qJ/O9iUfXrQEMy7pAOFwZEEyH0E2eo1YNP0uxg0IqCi8lfMkphDBoitlbnZTtLrgp2PFey7vW
XhbRovhhny7bW5orXeyH7/Aca5DTO1ZF1lSdrf17yzdWzoDjF/2H01GTBymWoGJGP/RcpinQiRIE
dYrKZ9XSzy8ggEhCixL8DQf4gG89FuDPZ1L5G+TaGVzGk7NHJ55aPR7ulEGycZ8uym5vZbzokMXU
ZD33Qbmk69xFMdJ1AzzeWBcnjgFiUTUaZlAjC3S6+HukbcnZyBfXwgY6mYL/8/6x4CFQHD5S8/tu
1PF4lsAIU9IlkqqqGNeuPGyDW4TmU9uqfRRBpvKyxGHirxZkWkHb2Rzj2yItU+EH9rQ4Zy58BBJE
8h5o7iu4orKDu9umtDJabF06JYvRvneFWt+6T7lSDctOxRYmEtOncCC68j7GnRaF3dLsFLfOXhMs
hXgmoXTo9eMFVoK+oNYi43f1v/KvtC8CNHySze9Hv7ww1hb3fj878F4rRz15YZDeAKGdL7Cwuhks
9AMVxCHOwBoxLXL1JpzMNhN2JISyNf87mUi9mCFb5ukfoywS6IstGnNX7MVu1P+N9EeW9h3jVBDa
DVCJjdrLprhIBh759V9AgibWR3TFTTNSHCjbn6JBwehF0On1DlcLCiyHzA88fOcqGa3S8KFEK9pD
+8u5qe9E1O80FN77ReIaBv1fgcBCUWVIYEq7SKK+OOMf0zBav2N3yLVERRdhUuacxGOx5AQsn5sd
OiSPuBxXwsLCZPd1qXIUn4wUzKaM6xXGQySTUUNCcfbyhFYjjEBLst4WAEXm1RBvINzIivSaQEV5
4sI3y5GWAqvZDp76FmtmSQ4xlgxpXElT4mj6epY3Y1PkxMWHhmAMYPGYuXYtDbLjp2PhifNb54y4
7Hojg+jxbaon4yoJhILxcGsRU6zsgL1jAe5+k/M9Ye9OaKDRJGgEM4quuACc5N7DzHs+JLeaCFiP
z+msnisOISF8tS1NDsYjZbvfmOFLwUvbrBFJ1GEp05BEmWl/eEU5X7ixnUxXYUHW8OX2BECwKjWY
O2y00sGcMbI16cjjCOaggw/brxiekg5OTwAfI7NaOHWXFBOlxV53h163wi8mvXT3d4UwgjLEIjN9
LbRdTxglmSrFdtG4L9kby1yd8ltDsBnnIsTuW1RxhP4c0OnHTNhTPvFl2ydbXVBSBgtleUa3279N
QY4GiH/CtCqhHxtFfii6kW5F5WRkGwObXPJYqAf44rrXMoSRv6/LLrbh8YIRVTH3jSoJGM0k0UYU
PdX5VKYdYM/XEE9i+HUQnhSpWCiueKue8KEWG3YA6hQ30i54y3MB7vSAPMrpZw9XLlPCYRu0unoJ
AZUB50H5K2k4PaDlR6Iv5aKQusZR3wyeV187VQHTphtw2l2zcLvdXFHtGKvkRHfRguonWPmaoDnN
FpmWKD4X1up+DJs16YOgSQwMEmEZkp5VL6IavqHkEOKoS5mHExW5F0VXM6RxFQxXSUW1zQ4PiZr2
wECBoncbf/otn6z21L1TrNCftFCImi+g9vgEwgAk8Udw1ivcKEYXQSGPoYBS18un6jvwPmwN8FYS
sYeI5n2ACyjOQrWZPWXMWurPmkMDOosFGfMYtNJRcoO/sj4U0MAWzOialFFDFy4x6LdsTjSQwbwf
bLHwthVwe3z2zpgk3yNWYZMuyLrv5431BJnY74qFvSC2Z0+blhNkIz7jYsdjY6+MMZFwFgL5NhG8
QXnmVTv2HK6xjOvPjlxC2ihqTUl4CUhM/EvKv7ldSU4F77VW5NhBoIOiN26mJILdfsULtvvF+x+M
2AOp0718IU0FThQkMX47UH91P0D05ikLZhRB7+3QU3WbDIJm3UoG/Q5oHRtvDGAwSjTDpPOv3316
Xlvi+8Vjae/VXdkE/7LSYVf6qQCkDkSxXqRYAJR+w2w5XLGosvCKsJQJ6b5NyDXbeH9B1Gf7SJqv
l7vPs3d1LUrSrne5WXgyEOfg9BkRB0cu3f+ORtGbBQGErUKZ1P6QocQmh1EHd0++qbhHf6znD3eU
ghj/rYXLvOYx/AnAjOgIOfw5rRbHOodjH9b9GTumoPFJMZqr1rLzaVXFug7sIHz54PQF24yui75L
JVyIyony89pKfcr/AHiljgFWS/sRonKCHVVZUG8X2mURqydkvMSMLHuRaQC94iS/jwrL/mvTsKEz
wJzYMz967MhjGpIG/ycXN7IOzvHsO+cFQUI8keqxuw6qwKGKB82DKAlHp5MtI6HBJ7RLQpVmkU+G
QmZFE5bkYVaIWVpOuIsyboSgLxN/NimSDdpUhVPSEvaydaytp7t/qNQH8hAu61EanjSO8hmnVcGC
DYeenik6M/1NUdYd2setYYRkpO4u23DVKxQwRL42cE3rIN7a4+vE0AgYkd4c5KcSL58ZG6sBQiBf
o8LGtrR5CIHWE+6MXN+x4gfhxWZH189rv2jlx05ckH667efWNueFcTflQe059A1PW21h71a19NWL
V9jtavNScGNK7lgJ9K99GZQflnpETOySlVA1VNK1n5eSTYRBFCYFHfmzponkog+rthleFlqgxou1
+cme3tpI3nzFazJflCUWQiJ8TwF03QlOwN3froV5HrTPEwrWS8RphRv8iTlSOeQ7FGRK24v15OSs
QYHKks2Kv12q6Ene392Qn2DvKYnwE4ZzuxjqYK3Q2TTSao4PAFY2AD1jUFnl6Tqvu+GEF017lWz9
/cFXp2/uEDMYmvBuMTVq32KjqGzVqwFcf5EydERIq8zLpTOlbsyb3o7/D/M3D7Yl/3oESPATkvrs
5nm8XsJg5pcp0boInVZH76oVgMwY7a4kZ0CRBhg7gRkP9+bCYipS51bOQZ0yfJJMRGDJYW+etbUd
CsMI2/Fvili2vcEDYkEzm0gCxoMZNLrNPLyPPLsBQBR+EvhbLN4gmHLt/hesMhszL4fBL04BcQxk
7/Tab9SDiwWqoPdIppkUAR+5EZRZV5v2EFdichqPNpVeonK0AfYlLg8SLvW6ejtvvhfOgSgP/FRK
QxvSmnDLJIKrqdpzQbnZjI3vvL3/Y7Pq9yZKK2BAnNwT6x8PcY4QxRb1oqcy0Y9Wr3kVylh5dIXl
dOnv3/be2FVtn50/ljyopCwfKzUQTi0DQAL/Py2QBPh+XjBvcVMt+bIPnn4I6Cioh1xyHyvA3QtM
ozNi1ff/4RiYKlCI+UsDQNmDVEVjyxou/F6KEzuq1j8CJJ4gv3xkFrxgMQrrLUmMJ6D11oH+e+WP
6vRbREHDLhI9o9upMOmGyj9EbUajVDvvFAzpJoW+aeHMnsh8wS7BoERn9dhE5J3EGEt3n5XtLfDD
V3I1cxKXvnldX+Yk0kfJ72Nm1hGEIbNUWuGFA4FtlLZQ2rQL/AIAuAzOlJQe6lH3nZ1UESX6BNn6
h/jnZPGPv1CqQYe5jCj+mpAqXZZSZGjjCn7FwdhvjJTf4TKZY5LUT63BOQK9FEoAjylKgC2ZF50D
bBzEcd2SY/Jg9D2yt4zvRqrgllI69ZnUYDJGDc6aCLUIMFcib3FZ1WG8wuUoPH/ln6zdWdyzJZ71
sKYwi7Lln7eXi3GVvlskDGFLKymkhhGTa6TEGnAHk1UcjhM7ohMAWq6scBqSfvwgoB1Chz5hWfVa
xwZgTPP9RLRPH/XOn4K3QaP3Fgm+PI2mdLhISff0ecAlbyKKHKWAxrk6iB9zHpLQbBgK+F68F7sb
VYaimDsuWqGkZ29uChfwF5756iaNVosdfWQ3iLzUBct92bxqLobdrlBvDq0/gihBA+dFXAi4qFtX
+y1DY4ajc1NKpgT5V9xHOovTt95OYgYoNhdlj+fkzxnN4uQiVNkjdqEsu6gFbOe/PbkndlN0mNEY
Ad5kMYSa3FRqOImqJMBuZETl/jgRFnxuGkgRCif2ScY+HX+Ob0f7FzdXGugWmvhMmwQc1ytlEgSt
Ohb1Mj8FngSo01u+jTeIC12LbYTQ+CkCmVbfz8mzzEk5T8JBMh1VZBmuMBjQVKLg+42aOnn+gRDT
Ta652z8YW9Y32B0Vs+rB68+kNP4kBWOSGMYo+lj439Nx/ihFmemtSDJuq4X98wJ0tsd/3bea7flj
30I+VDyz0lO9qGcGDVvXuALoEl5cSal1bWPH3HUBLMpjtmog94SepqnnpGXYvXX0sArd9HCef5i3
Y6RbM33VOTJzGwjzgGkRrwX+fJSE2cnbb+UZqK51ibxGUkA55yhvdEY8dXyl/n0mKDjIePBszQT3
kS7IRXlGr18PBHtuEgqeOMLHpXVM4tXCT+sraSdkPccs6tQKhrZFbQOximWtvGD6wyjG9aTe75G3
8reQt3x46/0bXzgD6vGlLFZnLuSG+Iyc0C2YygLYV79dv3gJTuVwdG3TY6mUCA8YNZ3llm0ft8P6
8MyZSCliLREnWDyZRmsVPw9rcsjY1DSzbjbvmOc4qjJo1EqzT2mgXSf1bqMvayytvZlKsoQPprBj
A6KGawr2CBgaNfEuDLFD7nGuKZo2SpVqUlKuabvvjCIlpCjiwkksQZx/W21d9bmuKfYOsvM2Jz0L
UnibHyAxTgbaJh7rVAQ+DcJBQhYvqiFLixfe4UIVfiRvTj2OwCv6lk0kxFhlenWxCetQmA5geSGH
E0rHzKDwBQngWlFbfNxZP/I0nppEDVXpnLTc/eDUL+IDNifHFhG/JGI3wTgj7gg5Y/K2AUpeKl4G
Dp2hPuHiIUvmnQ672tPFrue2NNxT0pGdwzgngCM8u8eg7n+Eb+7Vr+3BNDJpqjx8t7kJ+GCZAo7U
2UEEJNytjAiRvlhl972HZSdeb8vk6o07U5tgbdavWAR369rliNjN9b0iYmlguB3n4g1kKUvfwQJB
AGpf4FNbMFzx5KdXKcpe4dvuFK+pPiv1H3yi0VGtl0pIFiS+8HGLVw5gvF0kwCcWEIWFHpLu30fs
ucyZHtyfTPanGkUnUzMj21g0Gy2VbaBTaG4h4AA3JMR6wVI6Tflry+5OPrfo2X7eYdGO86L1E4Sz
gVnmBJgtOQhElG661umGb2ktiBOZAHHuQZ09mM7D57kHRNaH8G3SFV/j7yaUOisH1fmF0ig1j4Yt
1TzrFDeg9Pcb/klbYVzphlP3D4EEWdHLRgb8WNLnhj86P6kTYbMQCBNjlViA/uw9L/KCyC2l2ew2
WJ0mBSXdwpKD5a0o2zFsL/SSvLoElGzzdGIF3MDPVllAN0/SZem6Tdy3th7Ru+Dcd8QgqO9/4YDQ
mNR/ymdmit3kgLbOtrj405uO0wfjwrjq/Rb3tDu/WyJo5OfTNWHMaZQ5ccZ+ch2kr3iIm4NnxHpb
w9Yn2bNOtq2X/RSZ2lWAgd+2oelnDOm5Hoi65tG92VAq8oKqUwZHJFYmw8BVv6L6O1gGaTWI7ddJ
pMnyCikxTiVwPmtZOfRYvY4RlRAf98lFYeV3w4zzGsRCWmxXDm29ARzRAnuyuIpp2g0m83MG6gGq
1zxpsraiW1U6fJN1GG6k9D+hmN+MDK+pqondzRkkMOWKiAuCDvcG7BhpGQmFxvbzG+b5Py1Aair6
ZCyCwGMRvGVPMh2mV/unaBKtdqzxZGoBN7jwNFxGLEOff35rzOg1mR4z3mulAhlEFXby2HcZ1prg
LccsvsR8PphpEuihAhoT04xnbNbEaDqiXD/ZVLvYysX7vxeGm2CQtOmQZFr8hm2r+pBXAGJMsrHP
El0RWTZIuPWRUXbQ/etEhoPl2flRy+1vteM1EuFan4p26SwQ02HzJxfNTKH46NGnGsTLv3rSQkBV
ZtOcu6pQEiA8YS9JmODJYzLtSZkoCCE7RbVjQ/fC6kM3HmNsUWF+bXZx0ai5sO6viJBAhMaz93yV
cQvRJxzYEL5Dit1CffpjNCSoyNMzD6PZ8GGW2SamdkC/8oKDb1n00tAv+BZRulHZSIjTczoWlNqA
9ghVKD0kwfCJIArwDatf6w/JzXfH9kpDXQXjr3t1PQXrHTrYL/o9H1rMhoUlP/idxlT328rnR0Vm
kU4vYhFKMn5wbeYq9dGbm9K5cbnCAsb/d49elas4SD1dTbiVcoApBMKrNQg1AIQjhxVRpSypfgNO
PDlC8V6Csn/+dbLC9bz7n4W7C8TEO0+ketTClvmS+NZj4MBgI7cE6DcMnIVZwj7wtwWlWYwindXg
pBwSQAlQRZEiH92u7uYaLvo6DMk5b7UvHTdxG/RagQfrI00iki6GK1EiltZZ8dLZ1P3sgzpkkZWU
kiW/yE9qMIF4nJIj3rZi3QsJUFTybX3Dlbvg28+gvawJPZxuNjbNQ2hDMFp/dUfayRjp4cmFJNdo
ewQazsfo3+XSQRSB+3rthEtsmtccteJU5ImXUwqm1tTC/ljaniJENIcEW2hBGj9hYLSh0pMEq0NF
nO0EfkfW2h6tboyqQ5l67CnvMyr2dVBbhjJFvA9FZBjEL9iQFMScm0ES6Jvg1d6d280qla+z4E9y
4GtDDvUGc+p6PoQBvt5e2ZD1/8o6FK4L17ANUcpVzoSSZ7aG4eb0DRRwvxAQuWAQcNHD2JBfdD2q
izVmATs6bOHozBFw5GBHUE9341JmBRSoNxBvlPgk3i1KeEFa1TU/RrtoHQrsLEhY4RoJHkvL7Es8
cqXGHidQm17p6MewNqOg1q5MY0oEYBvgjY17boZp+7qK6jqpY+Aqw8Let5KOGA2c60Jnv7iMRsCL
dC32S96hdpjNSXpkzsi0XW6aKOLIxbkwmcIPToePJmEnNaeMG0nPNNGtzHhwHLqEc4SdZ+wzhIO3
FGGWiIgTAr1bNAWkMdGX5qPYNkLkxagrsw6B/WApd35o7wZXRrD/Ar6wY1s8XfZIJs+TaU9kRBAM
pDL0wGXxpcnNTPKNpdVr45CE9CjDYVDN0OChbou4DIYbSVq7FAZ9ApJ6SSWDxG0Y31550gRJnh+N
PjRslJW+vGRftpI2nSq98VRkDfHpgvBfX0ZcJLWf55mwM+FldONBaFarpK5B/5SGF+a4zLbZRHzr
bojbX+lgQgIOfwcdwNdqbiODAMzi4zjvAG4kKlTijzyrG3VJtyF8F1uH+zJ6IMY0oGmVyTim82yU
ryMsfIAcneo+aTcw+9DDs0el5IAfzAO/ANgFL5qMZqYgaZHdNfKeHW41lQeUdC1iiEHgsnyK4+Ud
rLKTv79bAWZ1Z+BdVytYBKKEQysoe77X+D6QUfQO37/s8Ki5Paqu+/RZGbUudEvwJmhQJoz+6mHh
th1qD+eSDtUGYbJi8njYkpPf3LarRjty+NrfG3Yk813bPyV/SsHaVUloXzQYInqKd3ZTfUxmUBkq
wC4j132ObeEolQ7Whp2joy7AhyOIu6WasRliFFcGijxI8MMRQQ88lewJaR9D3Q7rAkgPWGkU8nOv
bSqBQwdAh83dUxQus4GjnhM0VLqcAb7Ly4PsbcjjnSK2O8HZd6vqJQn48/Xwxe5z3O7IYJcmP7It
LIoahcGidiLCYLAAbv3aVygAbcjTf/lpFuFh0bWo6dGXby07138jAUbb2OL0LZdUTaeNrx/yj5VE
++/FWZ9CQFnqH+ynK1XmOLdy48eQGYv8tptVdJVWaX+/DnYJtd4hilnJ7nhT7JiyjYyg5VbZQBKt
M5cHlUktSfdLQGpdAR7H7yRu/7iiZx6ejuLzZWFW+lP3MSLV59q/LBFPkAyWtyrjQQkIJ2CGNlJc
r426FF/S7QxWaJJ8KEpICWA3Qz3cNWNivSEz+7otFEu99AiRLGTCfHylxXNGePTo9GaKGoIivBvA
G8P45pQdAyF/Bo5ZjPM4ufYX4xBKMtEFrE4ppTBUlx2h7fgxj/1pmiWmltDTAr+xGZejYX2s5ew1
/HTihVVnyVoPhh8QKaV4jTEsU1X80vtSRpT3NIro1qIxioIHlIeQMqGpdaXzfLU0wedC5gS1ETuQ
vmfizY6A+fg7rLeVwkUqKq3oE0HxpmWZQwLwqzADOSzWTMJuhqzKtcYd2Vx4BD4t1aRsPxfQFQDV
qEBWC5A8tMuZTbfTkKenpVfluLZwcuyM2HEBpKIbdGWvOPxPTm1yoVWr/+waeJObIK67YDfrYO1x
bJXY4hOpEHbCRohchDJ8AJ9Pg9Vz1M9ZMfhmavQzIXUIxWHpD4id/oz/rwpg+g8KMGGy+HSluQQ/
BEcomKpQWRpfhbjpQ+FmJHNrv2ND3dlHYbRHXw2ibzu2EXVKjK/Zvg28RS1vLZHHsX14oF7TCoWR
Du3w34N7Vvl7qZ646kxzxEEMVmvrhITHQ+/4HeO/FUA6bOPnjePewj1/etnpWHDW0vu4YyBe6odh
+oDslO9MC2zr137MzgHEId4ftrB7hKvTiQp8NNrpMT2z7qwrRm97FqWgpqA/0rMWRgaG3uu0jRGY
i9cKmjfC0jBBxphYsTdJKZtgv4H8tgCpcssnpY9J0jGsd8PPwmkLf8ARJVYHz4OsqUfSEq3S9JMq
JidWGuZrYlEFimZ/O4RkTConUp6zCJr8tkgxWnvKLOxa2cvNI4Q5wCryYCquXEgZ4sXNNZvAI4kH
IHz/ZOogVn8Munc3PbCDBPhVGNG/xe7wq1VrgWxigpUOn71uPh4d9UhM0Q0miOO36Q7o40SzQxQd
fq7VLRnBbqDOPQyfHsGHqrGhkgVeJQSpUAxJVt7huwZ/w+0gsYvFOpKY4PhNXpdtz2YRwuSwUfv4
Lkf6gviV5jVz/VAaZtazMK2GAJgwfuJ+CJZ7//k9MMlbIhsWr3GCYFV0rf5wiJzOQNgOUpnXsLJo
m/6uL1nZrpuTXs6OO3woQW7esoUGKldy49yPwu7dOMblPhRNxn5deTlomtSRE6SuY3ALw6QJpKHs
tPMtzdyPI1AARem+oGbVLRQxMm+E8gtUkhMmLrCF5UXTTHDuEK+uAUc6tD7OkLlgQ+xzRDbnBH1V
ZGn+qKpb4jgQedTadcpzCKCP6E29WfJeH30i+RhGmfIqMLAHLT/ZjCNK403im7/aQ3AzydIGOD1K
BD3MBPO2NsE7iCis6LB9QWqQZezghKwOsQcfRwX5l536fh5gPLd1QlQLrEQN7HHZV2zOk9duexsC
/kLXlJgdDAzbfXPoQ0qumb9eSlyzPFfWV7zOYJ7yyjILimx4FGIePe2klDQI1yY+DUB/TCYApRfh
3b4/n/AOLEmfCxyvE82yaS9QT6PeffQhYILKKyyVmisBMlDXldY1nsvJYXOiiqT8XSyLSSjSJMFI
Bt+joaaWPOtfda7sHCFb/sk1dgvHSjaayfaosqHO+jmt5tUPQitjUM43HiN1ts3SbtTYeO5bSgf3
xH0Yh/ddvUNFSFv8cpHdp/rHtwofM2AiMELeyTrsIdkQVpbfbPYLBlhnzqv4TPMiS8CymFpXO/ZZ
gaYRLI93v1OfFUB2XhdhdB/kFisepRYf5bJ855WG6wHmdG5RrTQdr0sN6v+XW2vhxiywNhk0JGRn
gCG56NP23gPDsg5AJCFXtm/NeVdskdW8tvs5grsu7K44sVaXjgPCyncPFksJBwJl9kCgD9zLSj54
KwiElJhtGu3zELCdAP7y7oO3Vqo0mhKlWqFgcVONQ2NawkTBTAy+FFf+i8eE5GKmFQ8NsFQ4LPIE
W9w6ogmMFMoH4nk+e8hk21rxlstoF7AHcNs1buxwhk2t9tQDAtjvvh267S6yJtcnst6MsvYdBTyF
UAHncsKVsIdOH6WKxHgy6MdXSH/zWGkIBdvN3AAX6wzT6Z+0vuNYh4qInJkyHymyyAQhJevJuJ7x
iyd8AKigubIeibz4jQJkGBhOc7o4L4hRXvKRsqDG1BKidRq2qGo6Auwxx165UoBL0BAGwPdBMJeG
ThEAfFySdg5TmRUr3Jh1D5qJx3b06DcKeq8FVXMUyYrQB3/WI1eTVTvHScL6KWnQT5UJsJpIiNc0
S7pT/HC2bK/GYDcFiG3DXOuOVGUCt+Q3eR1OD+xCaCrnBK2ZPHzpeI4zuT3eK3itAbvke86PcccA
Mpmw87oUiJweqHXCgN0BUIdXA96uNiurgRRPV9CFN12bdR2tQax05vd9IBjrdYJJX252O9wTr6b+
77gNFv6o+tv0Ps20sWMm6+/K7MebJ3v34jiwsA8eFPXw/6Lg9MFozlg66R6D28Wl9jw7+pxLHID7
JdoYT3lFVyge+bsNsnBc7dnLbRrtK2tK55Cw6mf/f2vHVr0cunvt4DKpzTOReksCVQv9zv0Le1Zw
U6G/YrYF2pP4zlmXKjCI0NeRaOwm49lOhQ6blMbj3T0EhstoDg6p8NFuh4TAp81e5GBmyTmfNkRB
Md+cYCBdvr7HfMVKNGWhoig8br2zwqUCpuU9CN/4fGFcBUoDSSHipnXWbVXZ/1GVX9MlVOjYU4MD
ZXeYIaenhErbT72jBaywyYPeJsJY58MqDHNAIwnEgzv7dY4vHDb8LVToRDTtAZS5ZceARBRFIoy+
e76ZjqxNrMdKAhMcFQlTVsF1hCHYCZTUWV0XfS4Fzrg8L1cqBLVJwStsc/RTabWJ6XBrBBTfszNR
mtBkWdbdhy21hT3lHHckixkSVu9NG4CzzOm9fMyxzMaUac3A2iNMzZ/8inYbx65dAC9WN5Yz1ADX
UqpcAgFH4/pNDipMQ9w2UGw/n7VVpk9ymjnOVLheNqMKkbmC5VH+EziyPqPoG22r2UIkJC0U2Gbo
Y5Aw+ur8qAuF0k18ujl7oGGgUmcfH8RFl6PRWIx1GewtTqrjuDAhRBdnxS/n/H0mfU1rLmQMoBYD
n8iprknEQT2ShojUS15lkpTa/1aGnyBIiz9TgcYhjeYYkipQo+W60/GCABznvMpTpqD+Om6RGQol
ULm5X6R73t0n5IMZk35g7rX7mMxq8bJwa02DaLyXT66Sw1vRwc5+YlwUofdpy9QKwW6m4408K1/g
lu/ls1eI9VDUIp/bV4L3cQc5K7ThArmvdqJLMk0gKPLy967aGTtSXqSM0tgwssVvrxnaOW1rnZaA
yBXDVjA44XQ02NevaWQNHGRSB/yvUYKVehe3gEytxBJli6VR6x4u9SyhlayOo6aFd7S66fPu50DH
gLOGrE9IKvNkTUF6y4JX7NkhMsSX/KJcno3COLpPmr/YAHU5qj1fxhCv5XfBrRMOZ8e8x4v/yD4g
noPtsONw3r3KVfAGt8U6eSWMYfxe98pWOynsn9LVlmJHZSoATwNfwJrN7Zl8gygY3B8OJf7+098P
+dezu5p0l/ZK3LxzA4wG2n+A671VpPJ2okCNBlqBQqHI1Cp/eiR7xGAlN2nNCQORR8SoI5DHebPc
AbcRcihqcOlGUOSywH+5RSVt/4lJIoxGThoXzVTxTlpjCtM510IFTwzLG4ePrNJZnPppz8AIYvCL
UyjJwhXDy+EMAH3xVVbbSU+hg/anba7EmdSwgZvdlmO2SEeEXNl2CkWuQhxfYGNqrfewVxiIS41J
ewploDzxjpKufFqTTTYRHuTRJ265tH8t2vHcI4JFZ+pCdKGHjjAtRjX4y/zCHk+NQr3u0tPeJ5bM
R2z6NxgccQC2gfDbBGopNF4f4hW7KfW6qlFx2E15IMkvQvXDjPByHDqUrGtByKrODhWYcqeYYuke
ch0dPNzlvFhGQ71t23kZ6jA5wH3MvgauGQKWW1mgE+J5SmCOdEn0DC7My4LqE/38UhXVP5EL2/kl
Az12TNkcV6Im6DkpVI0wRnNDx0dBu0cu5leN/prACbNWWuj9PPlS3W+t68HfreHVsRV808wfl0zb
1DEnCPzYv9tNIG38sz/3KfGj3Sj6UJU4UFPirzRtBEPx6t70IcZSwH8ncXuJQJL4SAF00Tmy2Yps
z4yCAt2zvwad0InoGs9daTWI5UMJhVy3ZREn5hKbmeik44fOhFqsAo647Kk7HLrliTNgY+ucPwlU
W8mBhwEf/XDSGFoYuiW3Kd4O8KKK5FqCNKRTDQXvaDf2MzRqNxdYtJlbcr5c7Ole/POPNOBYSEeo
MAdfkJ5ewqTN04BCL8oVlBSxKxyPhnjEdNSqqlYW3DAOJjxDD2imxnUDkXgpxo/kGKEbwUCAcVpZ
EZrdp5bPdF6qozq1sruiDnIba04yLOhufTIjjY89H+bBpIDu1Xt62RkFF+ZqB3Aua1ARsGSLGqqH
21VN8rXjiPDae3uL7yLxLPrFomGVmHUbfBiGJtd9wYeR6hke6NuI7afwmMdgmJxiLcd/w5vLNoCn
yJdzMbof5gJkku6Df6q1yAl2nWjzGH7shQshdEI8j7lQeIuKhG2fn3Etsrw24N3xSiLeo8nHDrxc
pnNSZH56CLUA2/X4a2DuCLQFzlXfGURZU4XQFr8XFXFHHvJwftHhz9dzv9hWbL8MWMfPLJfe8kke
WYLBVOHZlT1r0/9ZutjjCRoS/GRR3xQittATU/xqxiohz/Y9y5A53vlMf1LZjFXaDJIbqUBxtyC7
sZABqLxRAQEwv/mpJh0Bq7qBHRwItX4koFMJG8ASVBxZa6Oyizpe811YcRpKcrgBPlR1e32NGU2c
3FxIyBfcZMEO5EVne5k2hY8ZmX6z7+/Rm9GpreteJ5pRzI3lmqGphm+kAxyK0PPmHL+2h1aqsoUC
/0MXzeW2KT7YJGYp/bXijSb5iyZ9hMUIdsdSHFwTQnjKHzEOEJiz5m6JbAfFXVYLyHMNF35NWJQv
c7iDO0+5gb6G+p61zgbr59dRDtQ8YU1eA5h/PZgnpq1C0awJuQdVyWNgQJ+l+yR2D8j/7YY04aSL
hMg/L43FqsbPiIUf0NOHKwBrwn/Io/sT+AFkxHwGycrqigQuvQN6iTf5ggnxMVntcw/uvUMgo+ph
es+853BB8kc7wxJiDCWNug5Nhy9WFYUey22cCxluli+RjoIU2eYgKFW0w7NzyDMxY+zxUABah5bl
tw+0/KCQc0NAbDqIR4n1oMlFXs5rWpLsTK7TmsKFs6JClyQw4WPQImKabcg6ioUl/jaksxZxyPKD
l3xNHj/S3V+MmGeaWnPohnAn9NPsFLsJ4RXXMxfZFSGlBz5hmXg2oAyMxHQvjubLROimpLXov75Z
dZcgL0bgnWrSZOFmPWLhDmZk/jg4PTrVWQirPx9dvdoZrWrQUne23dZKTzUgrCjETNBrTV0G+epE
0SI8v69Pk4KaNBdrfaGRQ6c3kKWGKbhcU5jsc9QarA8UtrPrsZAYsxPROo+a5/kaOEDv91qI9O3b
ighOM/FYMu6TNvDknOXNWWKVts2n0SQGoBHKzkd6jJ5bbujpOxLQCc1ozhb1JwOBbukAU04t3A49
dZUL1x+1dwAT0ciypgcUSIzCGfOjj9nYCqVNgOJ/XacHhkhi889e9fkjngjPjB+2+G4RxKS8rN4A
3PmA3uRA3Y4fISMm2seoKnNmcAUNaX+H7xhlrGJWxEOReWVTF+HU2XYnqA8FkXqVNpOxqkD4RVM+
Mpa2YtyRA5mGvyAMEO2mSX78mPVmzOMaiukGG5X0tROP4wXeeUvsp5MZRDxYeXJpo3DM1r90Jund
PL72rXnQLLMXC2I0CW5dLlDavSvt7AV/hp+XnQks5O6LGSQCcQE4rPh5JovRLDRbLxR1o1ai1hQI
4K+zEyfzteTJgC4UJTcDZB8zJiZUl1s/kxh78AOgynYQjRgQE+6tlZ9E4RlFwFMrEWRiMLiIX3LK
16r7yqT7KgflRiWIcrGwt17i2FBJzm/CSrjaptWl1XYMNY6Tt3PTaEELzbJj1TgwRCtb5Gkkvfhj
wgxL+t4RLW5JsdPTHpOsiynR9nBF8mA9aKYlz+/SNwwJOgzj2CtQ2jbLKbsqK+K2HTz5pgx6zIvg
YqvJQt5/ekbhxvt4pAeolHB8aRIO0Y5yCNURMbX25wtm0caehG/au1g34coAEFel/MkEiXuCrEm6
yBkAHAFd5LeI8Zp9s9HBIO+1uT3EmfOnlpHKifCvsk/9ZqJ1Tj4o/Q+3VkRQ9NDi05k5MR4aS/kO
KEooE8AWolN6Wo+QyDSboM9SB9xO0+S0ZkXTAyi/j6aj5oVZZ7dlX6NN/BCiAGRJl1AMOfbV3rLH
Rq7DJ5ceL4fdXDlzGTjD6jnIX+NS+MdUfS3TequUll3Lu39LZV0/Hlis4bs6J3RRgkOfITvaqKf/
6K3Qw5TLwyiIqMP9A/vDHq9m959i+G142mY6VwjmAfFm3/trAzJTte/SF/Z5pUVsUN9Ebvtxu1r6
0GRN1KeAw2AnyhJIOhRw3Z0Y6h3D2ZZyD7fkvWJUQs0P56Hh3hBYhbsNTYYtfWzD8I9Pj5MXzdEh
Dq5Z57osoR8jxprFxLO/uzRiudnjKHozpElhtG3tX++RL6iowx+c92rUhgHMHemCoacONFsMn6wD
OFKNXHHHgX3ws/GWY580cPSV8djU8d24P4Xy6B7GviRsjX3E6bMqnHd+80o1uB6+Z9oNkEZD0InG
DKYsBVr8XAEKu4cRJkiHX2Z5vJzSPhBocYA7GCCQ0RG3mKVIp/Q4a8RVdeDadbzuDYdvatLM3dea
mWrcKvnYv0Lk1grIXyuoNWiuPwROeRPwX7P4E7njdINbiBO0XA/CFVNTNzP0Uow2eVf3BtKFd9yX
H9ukQVdUufU3HnkuPXaWdr/HQisRClhjNSO/d8s6pO2rlWUkpOZqYXI4fCwNPqrnm+VsNWp7QiCn
T8c7yDG4Toj0xF4Q21/UiuNF4h3tc+62z0B1mEABmaG4CSHRtXnT6j/88WucwAktWE4MmWP6HNA4
vFWI7ILcyFMCJxHX9jiTRKMuZHGXz4OMXecFgoi9YRRfuHWYLWPUwCBhP7ywQOnKP7Dvhwp18ka2
cmaqbqMBwrfI0I/+qkoI1CLMK9bjp1/wFaU7dr7gFOZcMPudyjK/ELgPYvOmkpBOoJRXZS7BzAX0
+6/vY/Emjk3GhfOqtqmL67REU/8Op/1gGsRWLxY5BqYQkq1Bj5L46JvGoe8O1+gtn4XUd1dI3tOw
TASYv7GfmLwCUD1/rMWeOkBK/fvAfYfei7yvTqiXT+S3LfuF/TzYRidr4agDWOEXubeaWPAXJpfh
Uf+4Zqayb6Y9OIHCbnRVlnnKbFXtl6AhFzyCJ6ZS6QYMsUKMXPwAZHNv5rhtLf+A3DShwBYLLbKq
bp9RlL4HjNGo9fPxcVSYzw4Oq1mbhk5dT+H4GIziTLXL+QbQDi+oOLS5V3hwyQOF7LYptu9Pa5db
abx3Mh3/8H0Cno/FGQqnewHY0jebx2P6Ef9jVgpehKGeMl+UPzHbDRPu3F5lnN9XP2c+AgNPfu/p
kI7Pz2VJX25f/s6o976H620kU3L/pMP2l66byPn1xl0pO0DphgcTwgb0YQPpjyLCHyzIETptPb11
/UYnpT08038dTSM8+Y3+hgYteeo5vdapGGkVu6ZF1uTAPRPZJw+n0SrENfBJtlq19EV0HuFKuuEN
XCqrIAvQ8KUKafnIt0QWej5DNl3+XWTSEJuCJdvG8laN27jRRcCeF1R36Qhyv4jN78wxG4KwcbmB
9aDWDrKxfolBpNxxzYFyFI5LMSF+xFNf/GTDpOYKVzTii1KpXP/yxaR+v0+oRGtK/EZHDeVHmy8Z
Zkp+bDZU7L440DlGBZUjl07b4Gd2Gkkcx4ooPp04PgXcsmAuQ3uQ9r9tbpSilXHgkCXDSQzqjOPq
jPpbENsI9G6qjpMwvZxDZYv1NNZ6qb5WHoPQgkQeGxvKjISYtL97Ty9RakMBTTs2bvyU/R7lOWrt
Cvh8KM5ypHdpjFDp9Z62txRtl2FZezE2F+UqeEgNoIy0TMcJ2xlvL5T8lzbYNMbK31uvkHIveKMS
SBziUxev0kp5KT5HSPIxC8XvGdHyiYQ3NFSbKo/WmjdBhoioMcvMG15g6CpwhwguBF+Eg0IhQj7M
B//qWwOkH33zunodzexCwErG4QMpVNc7p3gVu7R3b9U6KGwbJBABYjb83OskqUk+M8Pv3SmgFLJ7
Qo4M7pURZWRbqrljc4UER3VfzEOItFrRf2TGsmXE3YSUBJRzDkNKoJt+3VN4Z5Y2wASx51/1penB
k2enLCywjgj7ebD8r66sL/lzpFi+FPs2gqVVkKXZUScIulUweFIGXKbaFvgoUd7JJWQpTdBqikOP
uKBOmAKiVd8p724frSm3YGt80Q0UF+JHssseQthv1SB3+XcjPLTR6bctuMngT7emOp8qVOKFDBGN
vlgKcAyvhHN3VkLlb7gCpFTCBythnndU1ao5e3kQ9o8roqsPwCIkPRab6BPhtYDMF9XxcpoQ63zz
lgHkhIc0O+k395+tB16s6iRz1jxljNIpI+XETXfjEBZdEFz785906bsb3177dnoMcRABcV0tX0/k
2//fXLuWz8Khsm+2j8tV4Hpculo7XQRpxQ0ygNu/7b5hSf1X5iZfWdnCZSxcUTT+ewxtv/8s7Ppf
6Qopj/4e0dPBc5sSJoAfxvWP8WTY5IB8f1HOIewlJZLZWdqVwSacqxjtGzsVLnqr5VYhysm9EzX/
miAtqgbN7Gu/4P9Z5kM+PG2KDqqHqIndqfTYNIYirIxfF4tElSxbVFIa+Efn4tulSk/4DWB/QQuE
56j9lTxbzTAnN49Dq2/PR8fCxU/AUuF62wxlB4frgUuFz755E4lbU4JBG9qIP07Rvlbci6WzshZx
uCq8iRRPb4EGRHy1DwLPiqIeIgywTfzAtICX8sv/+exVNmywB8F1Ub6pnKvYNil7kfBo7vafE+eC
W72NKHjOT2bVlYiSvounaNO8gT190mDz9H8OyfiQUImwRexIxwyBVqwDPGbMFnYgJLzlYG9nNZ5U
KzttSZ0lJYq4sD2F5nnj/QlzUPxycqo2TlwacFo6l67/DX5ncB1t0lXUFaZmeOWLBeYpaayWRb8k
ltl0GQ/g+WG7tL/FFKrXaGameP1KBRCpp42fRazToTsAR62/1Y5ZO38Kujwm23zOetPtB/For+50
ZGxGzfdSg4Bn/6eDfQH0AhgdmUTBqtjYbMeOnhZSscC9RjlUE/24S+eMBalJl0QkfsUA8MUEspcB
OxT7Mei2riF5CggEGHoU0SkZb6UWUj6GZlhjDFesuZ4hbs+Tp62U7hTKQNo0qGUd3bFD1y60sRE5
EoqixroK7ykkk2LD7cao+sVLJnPstQv7f5I8DrAnP0Ka4qm2kbtRECqmZ4cI1/3x8EF7FfcUS/gR
8SC2cZkEy/AEieozLtUl+yiOqD+9aYQ9Fs0qpDRtPexAnS4PTZNXaLmPe+7lKqaV0QaLWVg7g8BB
qigeZCYzBbL7zQCKuMNQ+Y5QRxn5A6Nu71KBmTXjmiKb+eY4nz73JnypgSHPHhl0OXqigfOFkz56
8gc0nq/cgGM9AQXFwg2+qdvMNNV29ABCQoMpFwziuLW0PT2oSb7Go5ZIRGt9kEa6MyDq38gnuAJL
zc/NFkdYPUHsf0qk+mkSc3FaYLy22DRtaBI2YURhW+tEslgtY9oQjOizAJAw8Ia/4ZrQZTzS2F2u
H/Rz/UiTq9UKp+2/3DY70fnZrOi14rcwNCVB11UQVbVgemjc6oKnfskBezdsk8Z8NpLp+prh9aDD
A3lQOPwvNANoMyLACt/FY0Xil7vvI240apnuPwy19XjxjHdZs+JqOBfMS5vogAsizV+gxxVZz+19
atAErv05bQvlKscHLqfHI+b2WfofPipztwe1uFnwfNtLRJo3bH/M1c4/rpOc5XM0+NYm0KGcU/8Q
xks2w2nQZVq2umPl5xEUDf72SYEgtZwPzb6wB9qoxaGfWn/gS1Isx0oPj0F6wdWinnVEzD5i3HNf
UjFVKzV0iV7V6fVntjnxxN0Pd2Xh6+XseAai4IGvtCvcVyk42lZPACWAS6qL2aSfOsT4KvZfiM2N
imRfR2vpK8Z5gCAwB93E4mU8N2MklrhPoHwpxhHFN2DwjV4tMjHoeLJtvo2jTbsQqaq+Hvory0yC
m7FvnFvjwhhq0xHMIebwkZGncUyDlsdEKcyUMFEgQFzybA48yW7nKm2R0f+WO8W0Rnx0rq8XMNZP
GIX+mjABVyMdETYoq1QcFWH3DUBbBTepWCuPaIhyRVRvQdEMm77YdLuTWeONzzrMNb4P4T5UO3wC
7ToCsRAp8OaxOZSiK07tYv+HDcTs9G0z5vylSRN4KhhVfOorDy1k/C7giNxTTP3+Ds3aHFQEFb7t
6oG3JZXDMKFJorJAac11YbE37O7Wtk/AcFxDrwuehsBNR0M8Tn68/iqbWm6hSNrsbnhpNhBTEWYH
VOPp5wa5AjCck5cY6Krg0RrKX+4r19HipcI78Xz9e2yFzqfNdrmVGJNP7KLQEkwJF1m2u/L3nPUg
je5Cyq7T8EfRwGO4r6+iTATEOAUvETnLNasgieVWojtd1sQ3TyZKGYUtyGCa8TFBBpznHXvhyy0c
zifJNb0CZXRig0xf1GNUTqu05uxj0wGKSLYwWdwxdfkL+I+NqhLHomuzbH1HJ6sWjO/xdmwxZU43
d29aUMExHNDRdt+QIhAS5/AtO5w2ip0X5riZ3PPrgvvDSLqkVZFIeLYrE+KUi8twxpSHcREbz3EA
mMH94VsBtXVMvNcbnrKVO8RDPIkCDFmBF6nMAMhY1puD9KD0ERePjeD38BjuI6vO9gocNujgJxBc
asTvfsjZ6TjQYsW5PJIGm55Zlbc6m+lxxNtXuDsv9Y470t98PZ/5ye3+U3P8InPsFqAVAaRgemEk
EXscEaag5YUKHRc7txUXYIvpRIVKEFhAN2fS3vqeDpgA1NPqjJ8IKsKhiLLUJ8mI7js6Z4e+uvNs
/j5AAcO0C9oYWnma+2s55pGlg5JB1uoOgGZ093rD5grKZ6fvy9f//s738ArGhZrLddYwDCVxY11I
OydJxxi3jsbajxKWRQRkJOQo1JgSSQ082jQPLDbbvwqEuPY1JkUpOBmIcXAqdxsnmj8sDYikdAiW
2XHKtickinGRGWBnoic5loKAkCsFl3NDfmFiStmW+QSLdUDLBUMCNwEWqltmOdseJR0wqzUyUQJw
3N8KDaCX5dFASF2G+3afo3wAWhxMIxnKDZ7JnPbFRnA4P49JM0rsZaId/vu9e+BO2lNXG1do2EKC
ZZNOct5Hqkm4nkSr7UQ9RtaZ3ZSzWTbl75nAdxQSwnrFO8OYKpwRFNbY3GCjwOuoX50bZcZlzfiq
kHz3rlkEIjtAtoArAi81k2NmWK0H+WLe+VKidti672AWWfe+XobtWuRpEoFBQGO0Yr+4b7wKqoUQ
JG3ZeY8D+q0o6spqth67fyr92HSqOIo0qJWWhUySeAKCQyDgWct8KqCWVY4pZ0y2Gqs1IKEArBOy
Yw4844ee6OwNffNQV8EqkTM1Azobmf/SI3GmWXdZ5Gj4nAmWnOMNxqCuxU3DlurQil9VBkDGdhN7
HH5UfLgTxmLfL3oE/puG35QfQLH4VJRugO3D6w1pG284PhDPTTxBXr4fun3nQE3V9U4VDh6R1Mn4
grh54i1yTUov8qajTlMcTQQmysdziGL7fKb6VPw58dnA7xk45MtnNin2PgFTFi9U9NIs3QdjCGos
Arei4tPp6Bs/mMWi3D/VvMsWoZ3OG3T0rwapjaIJSmVUD7r/BfIjevsAH8QhVXxttfawe09cHgKn
a8aseg9xMOcJJGBBT6ELGQcrC2C3nqk3G4XTjuzqEfpcHb4BOc7090SNdDDxrS9NrvyyyJzR3fBY
KLSwplMtjjorL+jLg+pG9rlXP2YdsatozuHk1+axVIBA1RSy2Iy7vICWPbQa1Y3aHSr98TLV5O4T
NFbQLKtsThROoxiMSV5/zZxleXP2s2UeWoeioLWjs6Gns2bBfnQMFoGrUnNvVW5hJDgi1/Jx+0GJ
RDDemK26OQQMcMA91FumXVmX/H74iIo2uHhdwYkMUyIZ/cShntWz/kAGeDCo7VpynLZHWQGVV0nh
EW8F2OpfOT9PKlY5nWhViiMy1xo/qQD4yam4KcDjx5MfNfdYKzdivPn+lcnT1Co/uMW9pDFUoyAy
WFVT3WUmBOmbbdi2looSSU87rIds8xkffSd3zI4KAmNtscHwuKEgpMxwGAKTH7rmI0wOIuxsQje6
0PRI7AKBeC6o8lf4TQXOITGhTuH0UP5p5gfjWczabek/72DAL7/tVCWrD24Ny20rc7bmCQMPKAO6
GiKTh8oTdN3WVnuoaZRNQF1vZiC/FqSW4hn7UxTRIlWcT1e3e0/lCWU7hYDRs7Cv1mxASc74gZXJ
zrf/3zRNF0aExorDT1gjZOcG8Z+Cp5V68BRL+FEcfUQbqcgMwTGjXa92dNVd3d23hA/DXHP8GsO8
BPYxtB9WOg7IgR5JtKQTdFrqoOWbKRFc7MheAkKe1K+J2HmtdD6jWp1/MjRHvcSOz3y0O34t2nv0
GtLEhaXhr1Z5Jc/t1/ULDVkVweNt0vDxco5kpL7VtRiTHp2Q911Bxf5IonS7xOkeN+mycZbcheh0
2O829yQU8F97gHkfratnmMOUPUT27N5CNhVH6xlemw/eo5beKFD6pvyfp/TM7uzBne6yzRYpQhSg
461anLnoNhuPNnWo0pbpBtXib8l1wYSQ78ucorJ8gG6jRsT5BTEgdYIjEcGOCCjOY/cL95sAsP9B
mrQL+ReLP8lSij+BDRPpsRSSTnM84nJK280xtXrhOrii76tf28x+VXHc119uVW/gKuh49uu66UXs
MtQwi1MnQu7chb04Jm7f4Pf0GQfM+wCnq3mKKYHxFjgy9fhbsmQE+draS94yqOYW6aWHViq3uTNZ
EMwgQj4FeD5zwvO5Hv5IPULa5Y4AU02yRFFnRqdBKFed68pAWCgkTTEvo56D3xTnGUMjgrm64MsP
TbxP2p+8KiG4NG8ho9VO1KzP7W+6TQKhptCLLsqSen+b80NZ1I3PSfBpF1pmZdNRlZHwcbvwpZiW
lxrcmHoN0oynQa5VsUXbx3QQt6FZVpl0hysVNIxm9M1OVLi18erUZxOhW6r3mjp6fH0RlhSSUxLj
gthYHKsdGZPWVWHDEOUtmMdMvtNcVAGNbdoOgsPLwuYtZBWJ4t0z0WUcrhAltElQRdtiIk5xxN21
x1OFCYO4KNNIW83JlPj5CLTR8Fwzw/Qtd35sXjQrF7jzW7+AgpXFDxI6yI+vNc/5vkGdTeY62bau
s9IbbShxfP2/03KEv1IMSWw5a2yMcbJrZrOI5kpcjnVCcYoluZb4q6VKJw2Z5TI9wCBMf6WIk/z7
0iZttpd9PAOYnJPod5I3gmSZKl0b3c0fdSkzTPkAbabglO+b6MfSB5KDNzJeL3b1bv5fZS/4THtp
xjBXFVWlikxqF5hmbEhxtNQFI4L6w5RRF40mqt2KdKOQyv16d+8ifDWdRo+5G0SN0dNkpiJfZCI/
EJvCNy3fgvj7knjXEtlavoIYTdlKBY9fBVfHLI/owoAcznmufJI85OBRn8n+LqbY8aJ5ghKHJAhM
yUvg7rnFxQL0UbNIz6oqShHqFgbx1YvmKL4sBowRC3mhJEXebG1hZEBAUbklgz1csKUGzpfPPJ6t
ToXLqGCji04qgg0UgN3qdBYveQPF4bKMDoNhDWF0vwhWnUM1gqQAdTpAAsIGRDYIIkPrPx8cnEpZ
4vLMN1elazh7psWInjmCVDrk7Yu8O9/lOOsWkvzhjN17weXL22gLqdsnEtlroY8OUy0+pJXodbLY
iLiXa029mJebyC4/WFu4pMQKIneyUNRKAzUurpAh9DcXoKSlXVvJMs0rj2HRD4zmVYWQSQUN8tbj
jSWlLrE2kK/mdjm5z20McL8/ppVs/WoQX/49HuPX3I6qvsEt3/pH18EPkk39YtBRVnzmeyRtCRsY
ASPMuXGAbA79iPiEE9EgHuUhZPJfFQWEQLcbQJgFOP/2+1U1+JA12NDdnljzfgL1V7Y0yJ6xtrWm
bKfSmT8ooXtA9WoECiL6StYD0lc/60zCdC3eXCa5Olkwex9DKlveqUT7TJxS0jvkILJlugWq8aU7
EdZgUGtXkA9AYta7F2PSowa6SCnLdthK1gZ/Cafjw2OWs+ZfZlsbPvwvl+ILiVMIiVcXW+tNNGAV
9uJ1obYfJkTWU7l/IhWmmOtmXwJX9E3ra/47EJx7mZ8mF/AQAJn22EZyE31Qg2pEKBBaRhHhyYVB
ONpsErloke+/uvWUx4IMSjr9KEk/pCapEeWHQOoc4qsMR1huVeQzNoaekcn4nwSvSYQeErJCRst8
hr8KsTTixapM0IXjS02uBlKJVKEiCok63Df8jy61nXHw+liY3UTzeEkdR7NGZ+aXbIxmlT3w+763
bENrRj+TLEM6vMVeltGGI6eCZ9fR3eaEVa+Ar+3vvxqr6Dewy9JzqhanVIgr740yYtm/saEj0eCS
dXhblLHrN0d5bnbQZ+S71oj8wtj74cyfUfsZIwf6b5ueP/+mJaFu/433lfNqPAdDcaIKyeadxXyY
1egFdzSyjbBRnzP8njQngStojUxAn1lbLCyJcHGSWbthaJBWGoMulapLa51AQqT/tP/36Dz/9ELS
8ahaBQ87BM93OGo/TSWfKD8HwmEwVyzBS1aiq54ahs/flMzTYGXXdZARrNnbug3tO5hSJDW7FnYl
eu2qdSxS9ArQhKsRCyWpNFlVVolF0G7G6Hj7QX2H6a5qO4ckJDwXLZgok9goreM0Aq+deEItuaxe
QjiQW9p1GdPDfxCVvSy8QPGp27IPg9ftEiKRM91h/vRHPO8FmBuYnILEKNoGwlawWsdW9H/7HXay
g6DyWreySYCnSKytcnDx37ECA5aLGyz+4td2bWOlcE2AbmZx8josFqqT1ZhEpQK8c2ewd+lWkl0u
jYEK3wSKV9kJtrXTFzC6TrvdpLLgztNuDdemyE+opIs62S4Zor8sNtyi9Q+w5lcujlukYhaXmVdy
hos2cw1rIev52QkWEt+XQumgQW3fbtcBpD+sfpY0xxuGToOz5fnAZaKKnIwXcvkRBSTQm/TbwvkV
18VAb47yoR7pOF3zPTYT6JuvX0xRNOnL7WxKeepX6Yxu86kBu2ytWMAb5Ka3SS/fJjwd2QOVvPiT
Ih4aDXFR7WGe25CiM1PpX9/vIrWJ8pXOMeJiyWH0Qv8MEyJ/HMLYjg3KDygczg1q1rN6CqZYQjA4
RSW484YPnvjHN53tDFlEQw6BoffYgMTkGAndm+xBBfa0+qigAJ88tdrWoUZkTbdsr5lvl1dNsFB/
0DB2deXVAkXgFYwgdG3mSvVp3puaCq8TSP60Bok+aKD7T8g20lJDKwsy0J+tkiL6yWkrjw9x4b5P
CqIJW4cKPjMLHpoNp6Y1LxCXRI78hCxdHuGroVX93elDgbau0n+VkO9CLaL8nObt7RGokZi55gVX
3sVgg1Zz+aPvCtI2KrVfUeRYESxygYbV45ubyRXWNwYIJBOnGEK9vcCT7ZL3Lp4HTI/0H1RXG7Tp
D4b6GauLgsoqK2jQpmRuwuXU74C2P4vxEuQoLcw17yq4RzVuaiD7slnfP7GeOEl3WP5kKRBGAoLr
Pqa9n1BeLaSAyP4oAr+mqI5f7ZKeK7+BDmb/+5ugqCJ3XrWqoq4dZ7YOAAfiPf9cPLqWDkK6yyey
61I+3LdztbKKi1pFKXoMNXoKNE5CQewFM17zeBvPeTELo92UXRI/39vDO1EsvJcPzGOkUsvXDHs3
dQ4gEShgtPmLw0ayV5yw6zP1wVrEk6cOZBgOCpnKTSC7BLXASIFdw6jV4H+xx82A0DOgPYUTziqe
+yxM4FcUoIMei+E9peMz1SrsJkNuJoBe3DvkJ7YH4i7s4Nde1lzTsGPDvrBOdntpLh/D6nj9HEHf
o2HxEEHZixl8tJFFGAi9Rqe1jAwLmCYQ6lFj9FjYN0yY2RBxxN/gspsAe31TodZn+S397yjY9YDx
CRM3lHDduCyratGSuoSm3YtEwI+axZajKWNxW0jApLsGp06RrdtwzXfSno0IYGTfK1cxX/eUJn+8
7axQa5xipTkCSZ/w6d173ZjGYkkkp45XhuWDUqY+BX7V71qXn+2SJnMXyWZMXSVXATUBnAegOJ91
wYnIn7NmTjf4m47xncD2g15C0ZviAWmHUzz7HqU5Az3ja0AQSEFtwA8PAaFFn1wz3aS/+dpmpVqt
s4/sgfvv86foR+TUZFtDJ3H7BDNcekRqVEZhlAYU3lDSs1dkvpYbcUcVHHUrKtWOumQyEK92deVZ
gYyZm4P0FzB0vbUxR07upjiCSnQW3SPUc+T4a0S6tZcz9MKru0R03eDy7F2tlVl56rjTIM24pp4x
afrZ+pgh4BjgreM+HtOGULIkibhd/mGqZGPpZyePVorL4HMwo8JPPqFDotZ1PIA3GdRSVwcuN8LB
D7w81kDSO64r0FUdKxM6/jVSi0ovmLEyKvgJf4Hm4DQHqhaiGYPwnLmjAbvUaRh2mMKqnQNccmW9
bY3p8oGa8s/ISW9rDsJvBaakEcmIO5zhKdXQImfQ6BewwCqJHGv2kKr7vl1gWlf2DWEV7MJBkfkz
Ned4HoShPdwL59TwK4F4MDl0o4p3I/uDxxVa2EGQ49As1Z0+bpCbnh+P2AcRC8jxfSM7L+8nlPc1
T8/Xcck1MjaikKDTGokYnYRgoO4SFLMwZW5qJBj1+wsNttUDMNR+La6/EINUMIZlJJAmSlZs08Q2
cIgF/MT1HKjMXpHrHUpdOf+BXU4wC2b0bUIMbczp8rLHCHS6dVfAU63/4y7O+o1gy1p1bEIOa092
chpP1NPFrA2V4dHu193j2qCCX4tF8KVZQ6xO/2UKOaZb6aPedhMN/L2c22nFi7uWbYMoz/NujIKM
z/YgrHj3ZvRYKcrGkmYrsgZj0tEkzyPhSvdJwZTdKShb8ymtIB20g7SOsrMgxtO+//yjGBKQa+Yd
tZ9LmrnUFY2WUcz7/G6M5HrhXngnomBoVqYJOVMD72vgqScTbDZvyjY5YgFzYSyBQzND+rFlXnvz
xvcYlXkOJwFO5g7e41RDasohZlM8+eiYOITfcNx+JV4vrRjjvOFbS7q26zwTy/5+nOafsdfKRtH1
j4ZGHOsPx3pUihzNpvrdE1l14IIQLtmC+igzLW+GKj3BJogNZpdjW+o0vJWd4S62qG/4TK9Q4oMi
GhaYcLgqWomoP3bZkoCP9VZLJsZKayfP0HtjOmjsyaOQ+8q2Zh+rFJR2e6UVROop3elwEAuI/Usi
vu/Bp9xxfUWc+A/oQ59DF6DR7STeIW+GkhvjQmCSPVfHM00iBKblvvJLqH2BhjoxgwXHXbpeTQMb
nh+gLrfNSv5hEt2/sOTvOQMdU6SBHpWigpkJ94qP5IdJ6U4Gu9g/Kxl3sKEtuZR8R6W017bBGN4P
vUB5M7qLOsv4+5W4mc+g26cooQCWxY1O0wMcgsKO0O+/l5ZBZ59yMY1CmGureQxvNY6Ts71fwTp5
+kCvFWEb7yRahxv39+MMfrPsMjOup9oS+UPQHBcUQF80Zbo7U8nl8+rQIrqXAjZF5wCTozxnRs1H
QIc8pZMCnQcKNzeWbCXEyavDo8GT/1L8NLZVGhiMGrwEiJkiapLS8vRlszbdKDRQGdFF0+aV5abh
v3RgZiNLYA4GJAHxLK8ViVe3dBJFx61kHJT3r4pm3LZsE6WnhaXZmIp27pWq2HmobXoUcvwwL42Y
HcFGxARXX8WUWHeSPSUoQPmEAiroFv4wj/+IWBlB4rHjWFOmO8Ix5gfk8rrErXMct85C4PCwzIAg
UuRLhiMODUgXuu5EL0i4K5VTP4pLKCfIJ28MvH4R2lhJGYX0Cw0Ru8Q5/MMR+A+YuIgOPfBh94zz
yordvUoB3dj2h/YrJzQKzOiDNuUYvnNYwPCGXcf3M5m7JwIRMZDtCjyeGn3H6nmIXJVaqhxQG4kP
8jV4JTWmyD63Q9q/gOzajbYupCCT32oilrFAdfGTr5pLHhB5QZJW0ULOIRXdG4MEmU5ehTQ6vcV7
H7oymN0fNLGd9lDkyoO85yA3gh5Uha3J/x7Kca+cQ0x4StBDtaSQarxrxUgqBL46MLsz5Alx9ggi
GCYieT7ilVhzh58PwaSAvnTK3x1jc9lsWBIE5SQtAf9ItTjfUf+3Aoq6r9eXGSBCd+Dl6fffgTfM
xaJ711O9JDSzGjlx9iTfuerC5o10WKYfJfy+NOK64OtV4mhmdx3Hkif46x1OemlLxSVdwRSfuRVX
mSYai5RVAZ9g4JwKUlSlgTDeuq9wU+iZK7viQiPpiDtw6Id/3JbKSV0dAks71LqhNCWYDXcFAYgu
5LzQCGEmG6dldQNTf0jxsoDmMf9OoMWFr4MQG613341gumRMgQK1ElPj40zFKH+Wg9QCnKAeZHNH
Hu3mRWnmeOSlpS54o9eC3N6tA5LkJl1pfnKzzvwYUglG/SG1QLFzAfKbrsDtAB79JsoC4LA70aBR
5LOd7hJAtkKhJt1Tyn7HIn4Sowr7mNU5ajQSpLbNHReM+pp3pKUktU6GVrZvx0Jc0Ob0P9xtz4rP
TNjhMlGDLO88mlqqqOQQsKj5I2DloA0hR2mmTsylCoKI95kBB7hxqdz0ozNNUu8yHYtW7pOL6j+r
dBHJ24rCc4F+yn4wjUi1FKpshVo+BdmiNCTGFtKvl839s8OijPfUfYPulhuEeD3nfmSX7a/DvcNK
EEDqWQzgoHeQTXq1xlqwcru+wN/ggXXXXeMAQEgOmKziKc0dUMA4+p0q38d8RP6h3mewxzk50ADb
qVVflC79AtIUVtVepUcuBIB3rDzf0IEVrcbyuN4mGDQ/cm+RX24IN6VOotkP8JdO3cSgA7oT6e+8
10NHzfRBrq/gtAiMUFJic9xW5H4mdqjn6VYiCTvseeZpSfjkK+mPJIn8OGJ8Mx73sRVsfBjd80ZI
vYJkYJQzrHRPGfMyZQrXktKRuPMK1JiLoCtdKHK+kNn7W3xroW9rxkRY6p1X7Hj5fE+qEEnTFR/E
nppn0qN9ghgRHuQ8E2XW6bgkx0hrLxS0oIMOMer+lkFbbT8ZYD3eh85EmoX+S63g4xJZMTC4KwbN
2E4rc7z4ImViiyL3rF82xzFrkUmYHUcUfneFwUO0UMBCIsi8stu1RQTfDKF04etEPQ562e2n6KIr
I9ss4pdl8QLcSDGuQRMOHoQs0OEa77tGX1t2HKojrGtbsjdSQKLN6UR0mRBGVB5SU7TtcVjOuyZ7
bmMILhaP0sAi7eLU2GcuNq/Ot3y5mS8DI47R0gt2557ifcG27DJYGhd2PIYg8xgb8t49Ckl0oK8A
dUsazxjhLxCeOtsDP1Pn6aw3SHtMQQg84+N+/qKpIsxuHQFxUk/8a0l+PLhxm0wCy68eZC/+Krcc
OItc0PQv7dXeegBr5jUtCMRyStLD9TS1q8xWgVoKl0+XWf3Bx+O83j2LRriy3+fbh9l92HloUsWo
jkT8AZPCdJFau3+0tRZbp4r0EST9hv3yHEZcfB5voXp5WgPBDYemrDby8HOyu2T9bblPj5knx7yw
imFw1X7vWx8DJlhLGgbzDAhr8U3T5KVdWKHYz51SVgYD4lYkgr1tv63YHOamN+d8xSkp6E3AH8FY
zwxU9LNbGSJyrOou5du6eA48p1jBBj7AwdT7qJTwR+jNMdDQnnh9u9x01nnm/5yPx+eKkz/cvcZF
6xOqX471YKGyK3DsbQuLDS4JNYieGIZMQQJ6Cm0+Mi0SDQX6YhXqFyb1mi2h109R28IApTpbDKTK
g8LOSxjNmohJh6OG0AJDYhF9HCEJ0tP4IZWofNFE3YaX/8NrzLrGQ68WH/knZroVDmXBJhs8ZIdw
eHlUePY+nS+1b8OA1rrtraTc4GPb93eMEL+GenRk31Rji4PWqHiyu28Fq2Bgw4n67XqLm4eF+x5n
4oW4YiLGllXI0VGJPbTPR05VRowF+w3GGIqf5ynmrGazUlFt2pu497JUnkLYQZUVANJ1RPDqUhWE
ear+ph4GHr07M6aUdr0BVm/X5K1IeWVSyIsV/XN5/3VzzTolR6QyM0dnamTMXrJBmiyYtgGXZQHm
pFITBJawtyKBtJ/O3xtgWS+28CZFiCrVHaQqvxELwjfx9Zc9XNkpk+WdpHeNkCVTekzo5515m+KW
22Fu4eyQvnd7PNYgeJPE3aGlNdcULlK8KRAbQoWH49HKCOfV8VRKx/c+iacc890MG6FVJ+3ZtJGm
/I+1iXq/Z+pPIQguh/Luii9JwGTPeRJMmMqxPaMhB3jiqXKWrBjnTjXigygchkKXNC+Pn80nt1jG
jPmEH5dNdwZKT9jo+eRFYMQli8c0THcA37ISP32Dh5F5kY8Lc3kWbJT4GWqcIxRmfi+FYmcc/bCp
NlgcwJVnO5w3FkV0QD0uv/zyt7jYk9BNVfCrlewiLpVpMWzcNf5Il/xqtAFaZuJDDeMLsLGochrA
bcKzLrj14gtaV39Odc/01mlbz7ZTKbt4m+qO3DL5B3Wq3f+/Aww8Zl6GI6aY/+ZqJekR2ZGJMoWa
lvwTbhamu9j+eb/OdgMfXo2uBCTtsbHtF3ydXXhnMjYxzEUUc8qx7YukPqJGrntGigVeS1NMovkh
VKK4f7gkay0BnzNLp3e8uSGzAyy05iSTii/kcjuSwfP5oZnc/HAlRLDS7h3JL+Y87iYWA2R8rrGV
bhBV5VU7pCnZbUc4IDmKf5fTvF5SYXGN5xH/qUKH+8RNNSXsauOVIUV83R37AgzXVNigqd2powDg
kuznLTwgJy0Zxmk93fHd6pC8Zpp4Mcs/8YDbT7MjA/mte6/kjxfMJlR6jqDQbmgckTMme+mh27ml
MfWRWP8bn2mJ58t+ORs1faud21ic2+8py/ASFCB+roojQ3p+0U72svciSRwT6416p029fi2mu6jA
NyQJBMX3aim6Z7nqUmQKdRgc00lw2E6Gllh/trTo/grqSyVAOmwmjJK6AKi2aJTEBdodIp97gBMT
AfOHCrN2x3SMGEg7hlHV9FnNI1FYh/TDTvMrzsQkS1zH95G7xLt2gKzgajwCcukBuelg8JxGQW07
YxPlBI3w96a9PIEXdnVY1uIEskHMisw0awfGZIiGn0YjiZYbQ6/lvOpfGmEIiUvaoC1RzroTza1a
UOf6dlQ+/0s1HNB7A+LeRCJwT6tFzVnKO33pmgfiSD3QbxTS+shs8Rnz9LBGeTaFzWsYW0cP4GOs
45Xcr1F64BPm5TBGszohGusKIH77Si2NWvBqwp2JLYaWTDistjJHuslhM3lTwY2sTYbSTP118+mI
eGUl+3ixO7jr7I25QS71Z2Ycjw0N8bgK4tW0vGpW5Hty2fWi66Mb6wmCFhW3T2kYetPLl25BsMzH
9RIiVOAsL4CU8L7uyzpeAVE5G52MYw9peBOA+SXM4HBDmgBL0UHRRrWDiG1oiwMCNHgITGeGNRVs
Oxop2OYzdeyIvTeIwoxrqodYqDsPXQV840Qzy+GnH4olNlwyQJC0pzlF2ieQPIm5dUhvRLGhbWt9
D3XEMlpwXgFcj9W2EFoaBKNzT03YiNJvUF6wea0mQmi8jW8dyrjL0e8pPTLq096MUJeiwUwb6gQa
wCaZuSqlXHRvLb4RCvNUpr3x9L83agm3nX/88xLaJoj4d1PFa1ANoZAfcpGsOXEJK7bEqe9QNnzF
4LvGKhAuN54DKwGP9lduAP2cG3dfj681tuq8Aipjlm54vFNTtrzYMFuWMVEPsfnlVsK1Z+UbPyia
k5zbsVdR/m+UVLQFDIHniYvybRpH4y7AEzI0a/A2+e0A9tQjpXWAGmhejFqK/+yAHXGMrmu7RbQQ
7SCySFqFiWjbSlgDBvEqsGqUUB1CDAxYvJv6sY5lR68r+TP4ExYd1Oa3EWG1XaAL1wsKjpwUjwfo
NFQbrGLkvXihFxdO4qbvxnGgySL1WXQH/MrgCTqMQPXUTUkQdp029SL4t7UUd/GdhMw8uosk+OK/
zAIMLMyzhN+zOFouGSXJj1RlRfzRezhFLFbhIpqgj0DlbgBf1W2Hj+0NCqlKeaCDezI/e9y5KNQh
jM6y6LQTk0cvkaGcgUy/dn5Hj3fnQKgcy6+j2BLMaSjCYJBZH8f/+Rz9eYQCF4hMlXLhoaDJ1zEn
KxMqbwtbtfZJrWluVGRaDD8P3d+2SJeK9YfNBvF2WBItb9Vg6XOsm9t/Nxcqwcc99I36B2BV6isJ
N72mXhPeS2wCHOYipEkVVBPbIOwVkXjTISeWbaQ/ja4neiaK5eS4AdnlvJG/OSPMiJba4EMbr0XA
SRjxd889C/PYzDtBXxL1jQjZxQ3OAc2sjNpK9OO3lZ78C2n5xMUUzChZqS5mjQXveSZYNxKGVZaV
Bq1FRlA56r9hSfUJzMrcUv9XREbl24SqlXyGlpy5d8ThGAPCOuNEuwqzFxSRJ/BHwMS6m0APkB1f
PD6LsyLNPWP6mlH8pxyOPUF10wDtQYVR4D6PjlQADJjzI7ozGUG6CKz63RmS1badho5h0dANh+sh
jgqMSZ3w+QAQcaNOGTBgBOkk+REGA7XfZ70Dg2EFdoIaa/oBWfOdqnfSpLRT+UtctMCBkByL66E1
QVv5A5wCcpHLRb4MnIzL/uZ4W2SMOWGHLR32owBX6rJmWVCvWr536edeAF8tnfadti9haBbtqvLv
W408DnpRx6880to2taDzDxV9GsO2pasxJJt3X0RwynnXUZX8ZVyNMe7TLXsYueA3tZNwbys58dP8
VpFiRjRve67ILtZEJ38ZY0jcEBmbI8uyNPxHzWe8WdvCOTL0Ym98Yfir3CbYL84An+KPkaBcuDj6
uQ5foC8+gpH4bX02aLH6FcdYh5vqO/Cnan6md2JPeSPa4wxQeXTZgRWsBZMZQPmxsD8Em05GDreT
25OzDFAx6ohgC31SfeOtlCLOvgaQ31rJm3hIKBI7xU1T0cKQ2chjg/95XYAmiYbGHfOH2fxIuCE9
izIb8pdmuHyJCQQh2YXgm+oHSxE8WVpSKPzQkSuzMAZbijWrb0t8/pj+vGL+phRVgm82/ZId4tOb
5cFunH+L8bGv0RmJ5fNlSkGNNnuWmdlhSBZqH6sUJuRH/MTBmcBDJwoWHlQSXkTNA3tC6nDWjRH8
WdXouoWNO+OL2cVRAIpSIfFQpk4OOT9whi9ou2M7bsT+ymDrkz3oIh/CCHJ7MjMM+hvauyWQr84x
aHi02+mOHarSapx6mm/8+IAHawxf9pVaiQIUDQRj7bym/rFEhzftGutKWhbgzn+JJHekoCM7s8m+
27jWtKkGYRh1ftDZKI+8tbu2q2a7I3WqnHh2rtgbA3kLAMoPfcf6FKg7htJbG9HjT+3hQeZtQUys
44TYNhBWC7DNPcOjZ07PMeg0RBwTgM2SClLMeg/OttOg5mQg+ZV3ThDbyXUykGZIsaFFqIIY3qtB
kbtxvsHxAsVrXNpRfQVPjzhD8enLE2eheV++DI0AYIjiHYhS/LEr8flEycr/t3jZ3V+5+YVbnjx3
ItndLyo0I4m5EyVi8SVkLJNtXrBWtmQug3q7yuX4fehoVg8SBhExN/qwl7InSSgREf01jgd8u1by
IEx/yBuPAyXzMxPSb10Z9YQ6gq0W9Nkx9RAeJMGsuIO/sFZ1SpuamrIp5FEHcQ+t6WQ0D1iCCMX9
xmOWX33k/F/xMiwpPnjkGCYFjt5/7vQQU7bGIcS92I/+rkwcnjVeR1KjiUb0V7GKAXn1Cyhifrec
jmiFeyG0uTOwakhhqicqGJ0bLaSljst1HbKDo7HqfSRS7M1jNObnNa7rChJzZLHtgoel1Fy6ttPh
LivzLCBnzky3oCSrmWz/aEDRMlwrPO3N0Cxqb6wMHe2CKtGELJcthj5b4Zy03M1RlDBAzFM/SxiU
h6tpQJhQ3CgTNaoVFw2AhaPs5IL4QrTCRVmcODxz5utgVO8uhBwI0vUa5ER7yXgiBoAQJ/eQoEDk
CMUn0Fn/zNAseP7ziF45138j73VJyDpAKqAAxkt1qr2NLyjFMyD1/xpHNVXM+DIv09RB4w4nioiB
uRIWJwIa+gKJfRC8Z1ixpqKi0lvDjXRlPWlUpKG2KnoO6dowM0ffZ6QhmrOtTtb4a+fqMrssJSiY
vQVrBgVgoKaRwAOrdTy+2ycdvPFpg3Q7ol8xQ4AGBriyDbJ4XlZM4YIaXCM8eOQ/ciF3BQbh3GlH
dyDCp245sLcyqwI+JbpVMukacVdjnVExTr76Rdc4SL1AdTZyyONYdTMoLxUzl3+BW/uDP/hzRUTw
bnFCGy1Ka2IECLQHaoZFA8UHlON+dF6qFdJ11DbIV1ux59emE8Hh438MZke3dAsColhMID8tCnPb
0OB1bWOuCX/VJWmDgJthxPvMOephi/IAyDHZrnOxFarOKJygIZJkVqVW82J4I8oUAml9uNlJIheD
OSdNkmlwy0X0np3HbHlaj83yBzJE86I8FVGrec0sKWJQRKdeSxvCxYBbwOP/x/o+s02f5D2Nbl1V
uLt5LQyywjBnl6MqLmKzFlhbqCoM8ANvajqtPm/uI0WmZnEF/uwbLabnXtF2vhEUfilUCNOcvEId
QlVnUTAOfDeqYiQiqFOBuK5+alPsveHXtRxARdowSVsP8eQ/6pUTv9x6+ZuyEmX8h07m9FVGK3ol
xBwf2a2vczI5TuC5F8KSbXx6OIP1ROSBpFtQ+rygC0EfVvfLpsTA2JumofrEQcnx9MgPrb/yT+oB
OfHXOauNnnffKY4o5fEzXHho+4uDGGq2qSBpdOrhAd3e6RAg6jRQkpYK95YFEwvmxSOELe4QFoD/
Fp/mNhi5YLgZpVWWUARyE38FJRr5DR3MvOAMwho3CgxAUtAhjhAPkKBoH2GV0FJnXW6KV38UHls4
AiFi3/BycnZbT9Ogzk+MDAlzFXs8mcR7dbsETV2ok/KnKbwTnSPM1VbSR8AHMyQ0/Rd/2ApCL8ZJ
3pKqlhraXdZmEpa0jOROHlJbo6kPB9j3E1KxzUKel3k5r6bI8GvvL7KYVZkhWumbgTRz3fnyXPq2
JRjFJrbPx0wl/6ng14pJwmB5BgVzdUTsl500AeugPcVkQt8WQJNlB3VI0W4tQyXZt2iajC9jvbUt
jGn1owkbcz0Xof8md9d+a2GIt8z0epPO67uhqIrosFp7oFhU3BZtqBX9a5v5VC1oWoLSt9cAB7dc
OmPJK7RcjrB+2xYIO+DcD0FdG9ZcGfTpesOd+lj1qArmocdAsmXlRCQ7wiGohPSLxt1yhi/YIVKt
O42L96xw8cNlbzaWZrfrlYrkF4vh/rIRa2ieZhl1Xpytkfq56NsQqNB7Rvauw0ypt1laD6QPNoXH
+T/LXmMCgOWkaHaiKYBs4XwnBP/n4Hly2qILwIqXkG/iP5Vq6w13VUreLlHx2ASBsvD1Ky4J3pMG
W2QArlkVRe2qavoRYMRYluN9Rkxbf+biN9ukfSrfcbCmEITJegfq2S8MIwk/Yolvw5M1fvS1YSzz
RTAN4RcCEVDmWyMUJKxxCAT4XxE234s6LIDi6UF3X2tHlr8e6QNZCShXjJY9hWPoyJoB36o1knMY
9OGOqnMPiD5Z/nUhnFP3Rejj3ux65DsJVLqovebKPZQLJ/k3KAJIO3Chc33xeVTPJcKxtbJSm/7j
phtMN26RQZSCK34yyeAmoFuuEfpObAGPNvEcca/JwfSZrEZ/ndYYNaCx6leSvVzrPpSrY3MIXG3B
uSiMWiEs+BbpUFmxWtgYtTBm5wASxWVJt9vqNbGmQDxAmzuhN2ziH3jbHbn9WbHB4b5HpO7vrWaa
zTns8BzXgEREFPAiKBhaPkWkKrI0BvF0Ch4j0cuorRDGv65jJoAwFk1Lwxci2Z8gLjk3yxyCICBu
Xv6R4v7c85124OOHfPlvHHTyQd9i25QfFXd4V3DDxdhYzWm+BNjdqnYvvWwxns/z1ssmM/Et1lUP
szlxxzV/BRcflrWvRiGxg83W0yEwnq2seOJeHGxgC3kDKnghsapQAgm45yq3Z+iX1m7edCu1j/MI
9m6v80clDHSLi0w/IoyaMEwTPBclPpeR32n8U234wKFK3qx76lxzPOmpkfeWRYI8nvGkF/yCCTV6
Qh6MNlWHP8AwYF8dhU5fXGbOyCpkycxtOynijUTnb0ZqfI8fnnrWOPebE0S4OsnvXVpODhZW1YTD
QZDe3o48fuHsczA9tBYczmL3bhzNldIcjlUoAVla/dNAZGtCcT099o8xgRtMPZQLlZ04IB4t8Mmz
YhHjPJ+a2Adf/NRZbJi6weeauVQtsAYqaNDFZavEX7J6C+rq+qpQnazEqBRFoajVmBW+h3uIFIM/
fG9KHyztvgtFH3RLBywls3YSrMAeeRkBXQbizqI+HxwC2rYKno27VjGCzdgEHVwadqI9VuhdGLnh
JizJMFzi74EJkoXQywTGtZFOWTkEQsXF2fFECC+ID5cJrSNrxpnyA5VlmbogJ9dfHg5Ft9n+SH62
JKe57VV9N2J2t24ZIs6zVjJfp8nD4VCCakdaufHcKYgrF6d0+4QrAH5br0ylAuJaqxmG04R5k/kL
wswI2rOQIRQv4diowH4ZidLuu+wxJqy9lERbVqvhhvaF+isCT4yvnqzwcQ8ywPhgRMtOWWwqmwPe
YF6KyQqAtbEAt4O8ZRRwKctRsDG0VFaKZ9QPVNKGoHCrMQHrl6YpngsC9IiQPPC3sAaE3Mr8tWO8
pV0Z7fq2EmcQnfBqsZyWDN/XsxPM4SCitwzhGwg1UzWrLHHoHg//pFnyE6iGvV3AFyWnlpCFyJNP
BTqD6uk2n0Zqz2EReeqH75ZTrMfgJryPjRgiwxdQ6d9Orr4HfhoPUEgzxVKhnHNj+qrbdV1s9PqF
Vw6hRGysn9TE/MVUiGlZyGcJ7onnagbjrasC5XSExnTRgcG150GNzoVwZsa9umg8YpYZHk7PzpbG
TC+HlaiR6M5IaExOAmTVxciYIzH7+TTS7mFlIb31ixVspG5UHNyY3TLGcwIZttJ3buJCs8NaO/Sv
Vd1vTfVUx/AuuYYStFdUD7FlZ0i28f6ME/Jjar1jJV0aOuhlhjWZ+boR+5gy1d5dyW2i4jGASG43
fzL6gJotyjEDabAjuBhyg/UMk9r1YaS5gW87NnW8h0yRFevia8Xlh0qqTGhPPIhPVgOAg30YFb7V
jTcw4GYV91v2alVbDWyMw7+duBK5cRXyfz/D2zl1+0UM4UNd1hU0Gf6oJL0ov916uADm3NfCPxPF
ORGQKkIAf8g0/7ElYjr1elPaOgq8As5ilvG5EeBC3Qnmt+aj6kjSV7gibJiE0+lJqqKV5Ssb91+w
K5T7nOxvQMD2r3R84Vqy/FElFYJzW5Fh+wM1IaPswJWfd9uQ/w7lKcSLeU9yUukLqFz3EBnF02Vy
r/UH/QmRBDO3uxTjvkIM2rphLNmlVQRSGkPeUTHoxFVK6/WiSSHf+bhaY/8nN4ymZD+NIPLd0iZu
4zry745gkbzFHtvVicK7tUJTPnk+rPVqW8YJEopBiHP2GoIZ0WvdS6OIs8L2iM9WZsI1t/dk7RkA
yO+4JuLnEHRcrTQnyuwhBZ4HcCyUsXTfbVQPPWhI7JqPgimLcJpaiejJQYgAIf8wHVVKs2XNMXe7
MyLh1NNmoymjYVv9Op8U2S2gV6lNK66Jq4M70aKGEOYRE1KC9wVUx6R8TBdM027iAZC0YRX0uw+M
ItUwZ8EDM7qINcnk2M1dOxMwS06XzdPJr9VmyLttMEaUhMYar39WsvHjm8EK02GQ8ptIFPjhO/PV
DxFrKI7wHP067XWnhA2f5EkoyR78Urqj0RWqFO51yNjUEx3VOODh20KBfKHf/OOONE6Jq5NNzamx
WPrBqUXVVu59xq0V4rE5ozJg4aHNKx44Kj5bEtOND+Y45Nx+Z9Ak83muXBeFSxZkUfXC0OOKgYqW
caGMVaFLws/tnBeBGOUf2DgaVwJVOELjj2zOgoIIjcWMKRcA4sExPs9mLEJZecY4yRyEFD1JwY9j
MCWc34PJZqFx76X5NEtlexW+LEflt5R+AjN+CcKKR90FyD16hLTyw7q308j4cgidKSyEEThuE/4I
X4f8zqo/0aKBdi+ZJ/1A1stDCJAPN8Q+ffZVB1OfkEYIID5/Fvkrcrtx3r+OlrCFmmzi1DYYF0hS
aE0HBu3KSmMpOokDTc13xOgsA4j93qifWNo6+OD3s81dr7q4aPUM82K4wyhqkF/zp4+iue50mOkP
DUpqZcBt4LGtyb9IhJUVBP+JuJeBj69/Ja/dpfP9vldocWaQtXr/Zes2FKBI1++qfkNiK87vVz/U
caPg1QZ3v5lc84gDOQdxNFr1AU3dAsXkSpH1+EzgSVz7UpSnfQ5NMQrEtRBqrpXL8uw6trt/LYFm
Z7DiAm70gdZ4vqoKGK5DxSoNjal7QCMDEU1aUv1viOgdle234yhSpSecHN42JO+Ov5gIC0b59Y6S
MH/xLurunDvDIhP4/gDzjPHNIWIki+PZfSSE0ZAoAe1CCyi+Far0BROy87mu13IRdLH1AI9yT2h3
uww1CwzYmbhdJQ6DIStpTYSB7kYWwDj8hEu2p+9fzcy8SJA0U+6j7ZwIpI9Rorhh1gTJTHrmGu+i
6YVKgOhCCS6m3JYCgpst4/D+nr03uULiYaFNJXVqA1nBaeTEzttUreoMlT+HUdG/V1hZ9DssiF8Y
PKet6+HQfp3XHGfSQW94tYhISXtapkPjJOYKS+Yt/geeZghuLCHs3rDMxZRH9/IYNZJz4gIYg3ta
T7b8//DUOa8Lo7gVHA74SdQQ18vvlvaq/cCCXDkmnqTS8ZoG1g10t4FBTKVRta5QEayb0NCGBOv1
ISep4JrLwfZ3Xs1oiGkKn51DSxRoNvrhi0n2Hw0tVxypH33FGYtdp1oDqaGcFXeV7vbQua+CXpjW
aDvT8D6Juw1h/kmMQmqowAIAIQN09SJn21fXryUZ6aYqTwMo1F4LuIiub6ah/werhL2z2ko/QDV/
J473SWmPQ+EOJhJ19t3hNNmAZMi0OOj1lkjd0xVfsU2Hyot5fppD7jJ40uBm7JVPQCzo2IYDgCzC
vz8ys3/jupihH/JSHQRHNc24QlbJ1mp5PvQH7YaYdwUei+bE8Gc9UCk9ltO6DCQYUzrkNYceAcYH
Qi/dU83SZtaVTt3RQ/BNpkOt0r7XkxQGEf0C0GM0uMwO+0NQDwKcv6xkaIG0bleMXQLgC5GP6mGB
Xfwaz3CdMMhmUKfY8W7TEJF/WRFsHDmYnOf6h1TxXl8u/UjBPBYkOmcj2XxeHx6Yv/uaYYFn+D0z
YEUThLH+MwZbip3XmsuJxfSXwIbLU86c7a1o9m5jLTE7XOzFAJNYyyTpglnJ+rjrOGBw7fRi04Ev
IOSrtt5n+V4hvkXOvLelCYimHtWpd9GsEPqg8EG0zxDEyg/ajsD+Pwa6uwMejsgFEXQ9kp8JIcmM
4jMbQYWy7MU6OT32lT5Nt5nZC90cufkHhGkOCg9Uq4ofrxMMS1Uue+zo8YXw6WJSmiYm0R/EKq0b
mnYLwvhz8Uq9HXSZXw1cMc4BcZNoWbvGGmVUgzHa2Ujb3BpvYy5rmUIUhAIF2XcF4pwxU1VJYsve
LjlN/4pJcAI2KliGpV368bMNmlufPzag4p4Bd57Zf2Nh2LXuuXUYS1XzIzpZyU4HPMgpbwTE3Bbo
F7R7V9EGTeTtoKEWvyWZitOb4Iv3RGCTZam8RycSMJSMuyNPomT97ysk2asP3MKbsBuR+0DN8uHs
gTZUZ8qS6mQC8PCUlgC48KoCmYBWYUx5EoP5GEwndOn+jY+mBmXyCd5780O8TJy+2J84V+ZhaijI
QRZ8RCy8z0R/ngvUXeApKehA4eoP0XSkCElzL3v/TVhuTlHvXdeyLHkpQlh4Dm9rtlx3XWVxOfSM
d62Cv+nmHgYUYTLg3+RPtDia8ErszBZikA9vhjrLVwSbW5r6OqGj3rxJIOkcO8gOLB2ORX8/jRCU
Uouq55BQYf82n05AynI4dJKDQPCO42hRdej5vwGka1oBhRpJPRPFPkSWFfyqIY+/c3tn91t8AjxQ
otEj4Sz4dlpbiqFUcc09RlZmatJC0bn0TPPXtixYUsc7mnc5f+Vtux4Uqu/0GWg54X4ERU1zTxVp
74WIneKN2xyq9hFojsuIUaoMYWsjXNdtHMmkvuOiz7Dxfe41D1r43HiUpXFnjbBufJiwweNdWHPL
tcYL4hLsNJ3i7Ew6B1fifopEV/MBy4VRGWex1s7saiygGcdAhGR/JvmlJIrZH6BPRx93Oo6vp6Si
gBQBKnmg5lg3eRgd9QrP2j3yWbHnt34AX9HK4ZPbybwg8WFZxfcuGqllCtKOT1NIW5+r6HCR9gb2
pdtrZyi9EvjfpgNfRyroIrFxoBLSXbERVNbixS3chYMTKmarjO9UHCcvFfVzpzLaiIJsiZw7Jp8w
3+0b8Y9eECuBOB3uqZrcBVFJps4FzsyHnkxvc6WN4FIRxMgGntwrD7abPnBO3VzP9/drYDGV07iY
P/WhCm6zXa5k1xK7oTrz9EX0HjeCbYF/97dMRWBYP7FqetaRcn/j83O7k83cxO8rG/x/sgtSKpZa
KYZIOH5Qcn6ppoAdMBMGvqk03ttC8/KSr7z4/QR11bidOgAwixyX3HzNv2GhNyF1ReWvmKX03Ou4
iwQzlE8C9QQq/CYyH8TA9OZ2tlcFOgT2b1wLUpkB8/4DXfel+n9qO447zEW6rFe1gZXPEpEgWjjj
qknPbyO4ktA/nGepzEm5uTZUJ6RpED9+F+QXJ3CXEa2Uf4ZpXy+0FKKXdRbF9Lo+vvgHYO9kCb+n
f9tE7DVOVw/gWJJmh3X++rz19se1ZPv3B9hnhL4xBHJSGDzwIUTQQtr6r1FLwhFx/SBAj56GAsLG
JKuv6ymeQqACt/XRTVlKnFWdWx0q++LlqWTfWNVcO44hR+QvWBwZIbvNDerP3izKW+J5soI9jjmJ
PFbLdT+z+26mR1MTg4R4U/arKaBI4M2AfEh2XWTKomzdaVULSKT54W6AasfGxe1u6D3lZFdjC/kA
eNOzZLjj/8fgtMiK+WtwtFmcyVfWnyXF+2K80dxKl3jgIvznzKhrdTGl6kahn8BhA+u43figM+3C
djp/TGf7p+MsdSEWTkFdu6zDrE1s3Z1uYq6ZrOVcltNpT7hz7HkiqTbE9vbFllhONoiuGFLVe+Jd
NcuTEt5Z8E1jirxpwUwU8dJ6hyBXntIwLFsxNx4ExuZVDfONZyGKN75FI+m8IqD4JvxseAeLCHAP
fvK+uc68qaizUN7QjbeoCsva9CYOJIiV+EHB69DRE3q7Nj2emmKL82IXajzif5GhSbuqhWCct7P1
dZ1xOJ3HMB+9XY6zgz7Mn96CROUJfnfisqnMFXwc4BfcIL+46+byT75ZROsgwYFzYEJ9bO4B0J8b
iU5BOL+bihPEL321cULjp1O9Ga7QSZyutlRNZUzEgIQFpvqkoPRGgWytiaFoDWy4+7qkEQEE2Cv4
c7+JY9HRY3sVzlsmlEt0iH3Zyet83siGJiqDqoFCMiRtU21KUQfK6Vr+WpXEyGM5DY2a8LJmx3wZ
T+NZ2ac4/GAd/sk/D+NTjUDeS9kIOsbksAFRSPV9gIQUxgW5a45l/9N4jVK5ClpjXqjojwhxQUvG
j84JQ69hhO0hSE/CZNUt94BmtdEm6kPnlbbPG0OuDfCRGrtHZLU9TySxvyyyr4flyk287pWCvlBG
JO17gXRqirUUu2OkAePjJxFUTvadihL8HPh4l9jl45nYduJbXb7RCU38k8H9/itYZo/E7vwDKVxv
UhqXjoYLLzaKzhLtTE28LeonKGXveRKWBUfk4Ja+EDf/B+pwa9Ump4PM8nVglZePNrvPpK2bTt1U
uS2y4H5+YfhYNNlo7oioUY/CnKrJlDv3O2mQ7uX/CGToKgNDTzcb9SItuXUHxCjNv1MyhR+VFTOS
E3D5f6zxw4XrkAe5Fc48RQTLzDiqyUti38pDaEVJiP8AzRSLVuXwAhrT+5CVOSeb8JfSg2azcZl0
AfPcxJ9UAgfvLZ+RfgGEXXM1j6I7P3UG6DbRJdCQIyWbdVIArnGfSBaMm1hXNSv2SdSlD6UTgtST
4Hlf1SkyS7F/m28utmJWUvv2+2WDHZuDyn2U5YmKTcamFB2FtzD0BL0inILQsYMbXE7g4Q74Hj5l
IX8guc4FkSf67alIiZGymU8H6IpBOX7Vxn83xHZ9v9m1kP4DNCywBzNSqPbu8N8lEMcaAwua4Dba
MNwiM0YLpxjbhrXCSU7VfllwkCaVOUMTHNeI6juD3ztwyOA3cXjRoP/rrMuTykP7lKzvG2/zrsrJ
boHlJZFCMZ8doA6ShXAqO5raBNPSjWt+uPZBlivIttE5ByBDAW2C0gd/JoLy9pPOCsfc107TY+0J
bvY7mT7AvM0TaqrBt/RfQ/fomRFDpVytxB0/2Qkk5tT1zzQDdxbOzf6p+K4aBGn7GrqHVsIs8MfI
yJT2raPx3cNsUkKskhtnEPBRF2XNv0UQtb2zBddAoJ6jQKCB8Oz4uYMka/2g4aKonSnrIx9uqD7M
iqzqVqb8QnxxWj0WUqi8WHwZWKjwJSmUIunHW9TrllKEYsSln0e9Mm55NrUKuYn5r27KuohfL33q
bTFePL8YCFBKhTzHfLDJb292C3oylVde7hD7FscisiEedJlOeT9CLiJMUdllUxOE99c6HFs4WQGu
SlgwXXvGkebOOXJF8qQq/DR+NdrIBvpvn2hjPZfZ7uYPfrcEzCaqOuuKsP65wMACuOoIIYWScXaK
iQflK+4FzdegoxptPBKmUXYg2h7yrwjLlBaQqEA9am7GzMk+1sPGtgibn+yEvdxWoEj2YYmvdfJh
1YgfIP3erflRXb7zOMLnUt65GDAAQqB59tgqkJWz0qIq5OtM2g/YWWV1TGt7eUA8GXlQu0W0zsI0
RFnPJXSOVrRhxIhXlXLOhwMR5lQQrd+D7JnfTQYBAckyEWwgQ3IfDNn0bvybfxJU4CfiCwlYUpTV
JdB0V/nS83kBT2XbCFqLnM+zCdJO/T/IcVnKsVMaxqqJuDoinQOVHzA4iqkI+dsctxMv8gyoRtam
2rad20GV3xo1AOcN55e+BlP8jLOBKlexB3Szhm0Zi/FZyqzyFsjnk4oDg6bolfu7CBbh0D599gbD
Jjq6+bEtYfh6eGwW8uaMKZyDHyuSFJMt6JWdrJmCgfbzvL8OnP7Nm+3lOQ9fwrj+wbjVsEdK78eR
EROdgxiQHLcj8KOvqjNxnm/sO8UXUMcEGMCALeohvpv+heegbp/QhB4YyJv3AcbQNxmVCKr9My2e
RAKotMv8sdVxERq5PmtoFAwMxQTmFdMYVi46MVXTmt698s0qISm6nwswMW8VXc/w2mGN+hJzrsld
4PGpkSopKo0WaPAQSFfRzBnrDJdEsNMbIVi5LREbUpHu4q1DNmWrd61vOzgJxwcV+7ipK7oiMCTu
NCdjF4kP0kqHzyM6g+v0/3Wpwa+ebfUXnWcgsVcmnSxKEOL3oc9viMs6OPNXhfmo9LIYQbG/oGUl
W7bj1Q2H5XjlcCXZlDc3LV1Mxa/Z76TjV5THiDbSCL/ug+QpD3bd2c2ZmSAXXOQMy2vHnb65cCF5
rauO3eExLuOn0Wlvfp7/IxwDBJNx2OVPNGbp7x1DtAWrIk4kVNlMG/AVXGfuWrOKkyU4ZScvvcUO
DSXTgQH3CVuwxoHnSFPSCIXy4MlnaSSQjoBZvjsu2Vpw2EbqkySOgRb8EiqiZXtTAWDzpYjIq0T1
N0lOQUhWEM+ZaKvw8voFhesp3dFUATcZ9oqywoSM4zDKBK4WUiST8z/CjUCL3d6mW/LqG/uxKLB3
PkGOYNY5SA9MXvMgo2NJMzE3oWjxmbnr1NwVUX0PfCfU0y1R6E71i4hTrLNBbGdmexqalRU+G9B5
z1RlI8Ty3FrAt7LaNbTnWbh/6Sj1aoo8DWT+KUpyjaXTcPqPfMqPntyrWOJ/GEWz1UrdcgYd4Yy9
6PQIXOJuSM50FJgzpi9iNK+fII/12Y/PZeZaRu32BB7bnbfdzSbLjTcWGTGpzikUd4O060hIGZk0
CVA9H7gRpRGZhdXyoFjKNtsDJmcztS7vjtNtbj4siRnTaWg/WtE2GCMWhIZl8Lr2IwhKq0Hj9GaN
kbagSoXUG88PBjyBpVhTPOFTe6ffs17zKRVrypKT0bgx3I/TZ8nv5hpK9b0+s00H3VCTO5ZGthoo
y4DLP2xTFV2GYJYL2IF85QzqsAU+It7NDR+H9ehmSv7qWyhRWhfxNPaXq6xFKjSAj0Qnk+qf2PGA
5YzZ+oUDuz2UP0RhrHZSW9f1501OWqSfsR+yfyzWLFg/qmdQiryQ49rv/iZ5ZiGQtV2zeKYKl2FT
+FKEhFzOOEbWUkI1ZTHLWuJGgI6i1QmJH24vKZ41FB8V27MVJM7kKvp0hT8P8kyfyoe+b42fRRUb
iIMCv6erUrALew7oEP5g6cYnjeZCv7KF0zmc8HmaNXrH4Q70Ui3yagpN1sJXPUw4QUPeP3VVdQ6k
hpiwAJIFR3SMiUtLN3Siyljo/8cVRbOs8LUXjafj/hK9x/zm0XDNYNsfEnypnZn5kTlhRjFY1OMv
2L4HCn7L+xEAeizPGQx6qr44edUAuv1SZX0WgaX4kozrcRMcWQoYFGrzOiYzimxEEE2vm3F9C8iI
J3lyDNBqFY+9uoFMUnYYQq1/Z5YpBCmEXf7aKsirDD4twTWAM3sKjJ/BO+XnXQz2KdnRx+sLPN0E
WMXLMz9c5BGE7j6gfbCMikMgitZV+DvUr9ejosJ/zGatVkKKsZIlRg+HmZrJE3D/2/Bw/18pM7FA
lvpaZWleaooZAErAIs5vb1jqT/KSsZmMLnVjvBJiAFj9qfV2ODI3uWKp1vXFpadvFFOdsJW9GPIO
uvB8hphaR3XtJhorvNrJPgWijQ7aCBZZQboyMSMDgfRXDl7+Q6Xioljbsjg5wcu1JyXY9NYE6qGX
89q20e+FnjBdWndHZcGCysEAqAH/LCZvo5FURt79D3dnGWNIOu5rXCwoUa21tP44gmBr8L2xm6Rc
ATh3HDNNrIHJRB8IOppFAASiiJbKiGjZtotTqqJHx45rJQVmkrIAEgcCVRqc1cRRVt1AUf+6C3vV
2acu8U+ojDi1a1pZSciREdxtPS9Eaeu8/r+fd/cpz8EpTOCPTGIGmg4azO9N9LxjOnEcCUCWIMJg
leHWUiPSoQooQQgs63ncto+EBfG9/ZntaBBdCThMc9Iz09e8wJTtGeFyaKlWOUECx3JFaf+UyyGr
sMvLrPpCM1u7v0ITBcnY30t/9T0BqmPlrozzIThEUwCjP1g8Vkzg7ejgMq6PIt+xrSn2re+HWaOn
1qGMc7wCBpxKJnqtYhD97JMbqSGPnOrNCIUf7FGkyiL3RLeeO2cVW3anw8ytiwK9gCaUbhpnin/H
tbt2sk9jmMt0DUqKM4vBm507mSsVLRTIMLDm0Lwp+yIhoR8P1KyaWhvou0QIGcvoaHlFjDK89BI1
b5ehFmp2fezyKL6jO1TTLWJ4dLXcoNumCrnrwgN4BxZx/7/sddImZD1U6kji+OBWl6HHa2rf2VP2
3xOqykBpgUAZxvy7z3E33/TtanPutQ73fok1MLi/kLNeh/8CtT3PAgDRAcUt+YULCdrKs5gaO1R4
rV7C5kfDaU4Jj2wmBl+RFXq5YNriG+tTm+PJlrJIo6B7HWHpSzMw8/ydh6esGpU+ZfbesAFMLjl1
GYqxfQZek5w1TpnbsaHQ3/QLINTun21tuu3qAnioKfnFBdiDTkCHv66euDWW/OdYGt2OwSBWiH/x
gUQBIQN1itHO6JWuVOU5cv4FzcNR2I12UVVx+Sj9DQV0RiK+DMPVcFLstqBRzAovzCmLMP6yfDgU
pCnYQ5efkzDjCLY5yulBG44KXI4P0SFMJxXdUM/0Ug6Lyf+exsHidZeev9MIOAOjYuwfTB7MwS/4
c9VPeFioVecbIsqVZK5HBjqN8/QYkwAIkHiV67oAzAdU5mY5bvJfhbOW96lrumWe9Y7DoRqTLUoG
sVqCa21gUvhDBUjipVbcCiPi+DaWvClWKFCfWzciRRfs0zpMSXmYlY4DVqYd65AQr15B6bW9Hx4e
p56viANXoSK6jrQ6plmt6DgpIugpxB2/TDKgxfoIFEgnt28nQqMItLrM2h7bqZyGB4vwDGHp2aTK
u49F2sSNArkbEHP5xDK7chtwgQnHd1K4DJHfheBOEAWjGNuBYDr3I0ExCyfDEbSxYzm+t9faLB/L
UqWDmWQhmy0Xx8VDfqaRAhgcyC15dt+i9h5J8PRCsHb2Tu8BeQusOd9GmDrmOmCEiCnyfKvLaTWA
XPkCVbhwoJKUMM5HhOGGl2D9ANK4pVSTnQYjo0ueqTPgJUuFJC2oj7ZuEag4nvpdtjbnHUq97A91
tjHptjB6peMneJ8zurAxxfvM/tI8OEvDYk/8Cx/fdyEBpvMsgUM5LqdA+VGFf0/b6ylltEed8Hi9
cCx6DagrDl91qNNzZ0YN9j+QEqSzB7MNnaPe0BjxWAQmDY/mby1qDpm8/u/BFlbmGV8BfbHozRJD
+694MR4Oe9iPsUPR9ZL35jrgw9VmD7bEvs3lPH+UJDo0YayJ7BiD5MDOcNDGaGYP+hXV5Zs2vCE1
THuZbZBS9mmnnD+BbHENOgYxUb0/bHnGCv9PpgPYAgnZT2Sygb3mfLyB00AMYfpZaFAHlC2/wgwG
+FWVHYhShKnDB8TPWDQ7oPqUaYn5Xp0fw9gmj/NphRcPz/efk2833h+D5mpDd/l/d7yzeDAejAsK
FMoAoMb0wRAtD4E6zAVLCqWEEX54OdqusMDZJRE/EjtqcBYHFonvLDtFrgTZS+ukQBf5VAXDwnfk
1yLEyXybmrsTiRZzUzF36lXpF2XME3T386KZEePFBc67N0e/U1nyTNeJBBIYjd3M451j8fF1lgIf
ZnOHGS6FhWif4pPvA4OYUA4z41rWKCyf1B0XdY3S+vDME+NhGcEnT+4gLFKk4Cw5S7fmrSBU8AYg
l+DkPhb/9B2wIXwQBp/K0Vs1b0vL6fH8zpfBcDZMMYPgMsBvWzxPE+BmFpWUSzIVezVdI2/W1V8f
4OW1jQG8XjgwT544rytud2b03sQ3wKDAEZ72iad2AkHsU699NR/zxBh/QiIXjopAVlbCb4UCzh2X
JAPAmDdjQehQC6HoZ1W5Y1pUctqCDkIUlR6Z5x1QhHWuxasugi3bbV8voaKnHqOXXzEOziFEkRq3
q/LP/l6+mEOCdbBof7zmb6nrANYt8e/uGB1Ov9qQLtvPeOdHWFbinSaiYsnY0lfyPaPDJ8/8u9dh
fBbvTzZ4Cs1KC4/bk/IWwQDjgKAK1rMyiTdIYZE5z9SuCfJ65Y4RpPtUK1pwQaPzX5f7jNz9lrGh
ez3u/OOR3zLPm342z/04OYc42++3vxcL0au2+ScSUPw9Zj1LpttA/ntP5rTgu5mVw6kVC0XLWdTj
/dq+aig1R/LPHZnUa7v2hGO/PUBUQlb5HfTpMGnhrVmr2pVlMvIxuJGIgR3LPA41TYzbDrsArfaO
jXTM6yTd+hr1WCGiQBnOUH/QkLTn3M+rVQ/eYOAptMokqRV6BCE24C3MYMdFlyXfNc6A9XOu8LCh
EBGifN7HyYngToStAF4iMRtPkHxhlNi76nR72qUpQ1NQ7985WK6irIOUCdiMnSDSawLlvDvF3fVv
cNFxOGl9phnPqW+NfiwGF6f2pbaIOZiPGwmxS5x5yPYgH5RVgdnlUJ8SoXGhdl/6qzrDLx8HGhz2
B9ws2Gp/VdI4PkgwUuYNumhkjZe+e/fTkz1cUrwGJ5NWKBRGZBrZnDfI2rYHCzyvecdzRCBAAt7Q
4vouSsGl5IEdBQCtUfKSlc34AgPtQgKFqj8PNqeRBy/4KyfGqRdf42kbESJ7d/J/Kb/3HV6I4usb
7SooGXRhopg0fdQCsI8837Ubls+nIbKppoCdDy/s3wAkpY6sW0lo28Bi8ig9sK7vYB6qwbiVqEPI
lY4+RixApWnaY4BnXa6UHHdShiLnHfeAhRG/hZzDfJ+YzbASC0x3SoWXQbsGUUUq8Gt9ULJuCij+
RLpVPX239aIuVmdcz7tLvRPqi39ND83C+30V1zg3RvImFu/nXjFAMz5nWjJHiwVEuxD0CKFZ/xEW
2du/7L5un6ithbBrnrT3C5jydBKTKAyDKJuo4EahKnorH7J5EFgR7WUV7BQYeiqtttK5DlNgGIeV
vPtjGh5Oc2JdyXFizFv/67/bDbsftYUIwRkmgvpMu5hO4HT9akOP/ws++3eNGiTcymzt0SW9tQbd
5AXxgUZAYlcwEmXb2vDesJiS5YWAW750QClCgEr/RE+rbL1ybP399NATNl+MTeEz4CWcQTSUNI0B
hKyFWf+RZl14jK8lodMs9RyXrceYoUCSdvtz5+kvLzSuwZyT41divWQPbIwDelMI2pF6Vk/DjUPq
wP8xcnTOLWSM6pzlh2DzRFdLKTYrhmExkdBLxdQy1QhUYcYUUwoGyOZisfCZZ5YHHcTxKaNZHVVB
1HXBFxk4YHdx2uU6koIS5juNOJT1lfTQu02K7yeFwi69YjVhFEsDTdTHIw1VqZzUw2+z62j4qIPv
9yckXiwgB+xCnLUkMuxWO5MjVVHuNULyVQkPma6OKpOaX2VIW7N5cDMcwvLv+NysyzjHT55R0Fvs
Xo30N7roq1dTz2l/4DnOewgIbLp7z04dq1pDO2sHUZgTpiZpMFhOWTte+kaxJ8ZkoIyepwiJuxZi
ZspMn54RVyPE28LAHcSXvRfRIQ/w8cWR2+o+lM+6Gez53tPgrbeNSpFzhO1E6iY+G6vlw1pwXxBI
Hi+gDmhyuxss4WhfqxidJmGlePhsl0dLqs61XfAK7Bp+KLbWTyd09mOAvy2/uMmNHte3JRMYrNUT
26LU238W6BhJXOHemrL42MzVRDq4G2HWglkcM775GTIvbMsWKARjg+tEBv5+tedAf3C34u8uKZlf
71JqRVYFJNJRGWAylVYWfpCu0tqFe1NSU5Zs3zXQpmWpHvfsAXnz5u0B/pD9gsPckYctHt8laacE
XLGbjnrqd4eVdL1cqyPDXej7QE9rknDjOw/hvUUD5s3+x65tyCSW/uFJlNn2lTkV/qwbXZIyQtZ4
0W1veIJJ0WbUWIm9csZ4kV47eiel9KUlWFtlyM1vDD9Z8D8dYfkmjxoRLy9flwdESRr9b296Zw/i
rQtHQP+p4aZ/2Y6FNfQBK40NZi0ckWj/d2rfvAG+y5CcvOL2JImmeccRjvoJmf38r3QwNAmQ7Z1F
FLUq/2pqIdbX4A1AtUMNSN+C9jxB97zWLyhECQWToLo+bk1EgvnI6N7JD11mEtTEGlAkbymnBgBz
bJHfK6lUPdGhosvqHq6t8FmwCp8Iw/t3iOLGXmFaOJd7LG83UyoMBN9qfZ3VSNdE+mRFDLW0E9HR
RMXEAKTXySNFLhtEBnT5GiwSMC9ZLa7aPMA2y7LP7QlX7L16PWlZPRX06/9Lf7L/nTFN3SJtZCKg
zz4iKXAym6PMIHyWoM0C7pPnich1lgJDKqeh0A1s2/cyzUmGsR2UId7XIU6fV27imSRspQ000EA3
oeI8AJs11PedhHZkqOj4WVfVgGv++OOg96iS5d4rVd7U/wRgfuO/24QkX1L8+mW7lu0d9jcwF+2c
BNBrRGcCPuXLUX5Q/0fVQX+Wg97ux/7JWO41Q5sb1rN8U8S6xOuMpdBY8kJZW9sfVyTNTTFhPyZ7
whdyniWz5UvEE+ayr8bl7ugmNfCmGes5RoC5pLDMCBpsO4H/Okfx+iHJ0LxqF0XjWq9xzAtKtGJw
Aj2tlp/FOG7u98i7tyLSXVo+/21dEUI7abE8JvBJMC72vixX3zmTO8WGMfCCUwK+DldFH9DxJH7e
3myT1Jj3fWbiT8Rjc5PGEzbxRmY/AYszuJ51Yckl6Ua5IsOBsbgRHsk+OyaEjI/G43w9U5Ne1we9
lbDJf6D5YFAEtRuiIx/vVEuqgCZPD1Sn6m8TZCop8VcoBECLmPnhWuRHl2JcNi8mlCTh6cP5vjXJ
9Vos7uY+JlnENAsAedeJszxMReA9kfNE/exmLPuqtB9bBTMPbZYDAuQnyqh+0zFsi3CF9QxN1uVS
10xmR1cCVTryzpiLwdAP9sGNEqf2s6sfUyci+1hCKCcyPDVBgf48Fi687HDs1tJ/PhNechvhr7EE
DKaoP9RnNIW6HbbtU/vhrjJldfKbQmVf5Qvsx69vo+QAqLJisE7RL82KWQd08q7TYskGaZ9YjnxV
NVuYPRdAdP8npDW7B1QfiEd7kkHT+JOI3eg/CMUo/K7grCnJsngTeHJmblYx7naWyLHnIKsx6I1y
77tA0O9YTQ1TJ8N7KStgU8b6jl/cqYdjCpub9noEFxyU+VVMiF5i1r38TY/hxlgh+Css+kaN563A
4pYGMgKSJGuJH8HejRaVGwYbXyueaPO76Wo+OhZTfXSI3L8hgIHD6K2A65GBrz8HpIysQQWGnQWd
mvfedei0r8ZoBBKyIMyu4ZumQ9T5VeACqEBjJILIvhJYyCiPIiZR/HkV/VmSFp3Ix7Jw2s0uaGBz
Q4qlxZzijaQkwZi524Ph44iv3nQI6k/ZYT10Ffbg2ZyF9/XEysFcJXJRmWmxaiXg4MXCp5tAJiQt
AY6kt+5SmCe4T/5e5z4mMHj9z+Nra2srrS1ThkObT9q+GMYCXGE7LY0NBu5HWvhwitHAEcbbVWrp
lzN9c7nKg0aCL/I5jBDmzcxfaovRcxn9vYAAIaODN5U3HSVRR5ZFPia6GtgO4w6MR54aAawbavEO
8C0xgYNKDcHer4UdBzK8TMO+SNTDb10RuBWHYwr0MExypQWrnTikNj92yg+m0h6qfNnMySS4XV1f
Mt+g3KzygyyCc93udxdPrqsbcuI5s8CphJKjIRfN+hJ6BvsVGVbGVZR+U5Fcq6YucCcSmelutL6V
YjsaVqh2d7qOsTPoMjeOQ9zCuxxwUQZQ1zNhCnwx4X2bAfCe2Z0tas/iPvUSuU00iNr0lNGiav24
ogAtldls4dqeTq8U5ZqWhB4NoXDwReEk7WxCPBPj87D6gY1jCcyHkFiaCmclKThn07aBSqrnYKHJ
jVXLXmhPKYqEvsnL9HaBot1VDZIEtASxZiNXgApHtwZNxmmUWzjTQslisSRJ3Ybrw2Hte3ijbEth
yYILWKa8nT6+OZ0v9EWaE827Kn6cwPw5X4fw1I5+woVdu8FLByVFEHAMZSuSEqXiHjT0BzTfdARb
GfpQRBU3CZTPYAKU8aQfGc3xXB7LOjaj6ayPmxIWoYbUA7RH/gxs+SWb9HC2WNE/sSGxWXQCn/54
BmDoEhYPoQv8v2zkdlwo6jiapfetVWtkUjYImkBsUmjAq7u46/NsL9vLzK3cfZfEufm7Kl9ClXnW
/HhsofGg9b5ipZ77EGm7zdkazUMd8wITCykwFZgE9wrEfOxFWmK+FqaHkBO2puUPZtC8nT8A5sfh
qGSsVfuFfW8Ob9ycBQ1fnyaQCX4yZXQjvBX5FhrFRGVrtIjS64ZLQfGTuqjlNsdr/s/s8o5S8dUi
NLQoj3M5v/msMpfw5J7gN1mPJf2OMi11kBigN856wtig1WkALStarfRZw/PDqMhQcOFnC+i7pNX5
kDQodFvvHOO9/QnMKAqRDOpI7ZBv4DlZPiNtIXItdKX9PEXD090IGfrnsXj/yqjK+V2Qhqv4wpB6
MPPDHOFtJvDv6x9zmT1P0K99qEL10KyvZnkysQoX4LbLApz/BXCkJaWBRQYujIsCqR3zolEHcsAw
Jyllq4eGCs0iaYcg+VOqGS6VRHXTwiVUCN1r11SIAhkZaeaAsEYBiRAqoMRQZYH7XG2tW2VufyHC
l5TbJ/5jv5O2wa6eFFpmlR1Aqm5/Zoys/lfr+gyBb8UBsjTpwS51vqMb+igmj+g025DcB13BKOxf
lUCvFX7fpGsQecCaM7L54Hphe7u/NUsqKIQMbgyREGZkaCT1HGqpouPI11WhsB4LlFmqS138pjJE
m0dtT02nBk98clzDDob/BOCv44tr3N9xoXGDW+jx8wdv0Cm09rwj4ZoHIZcTg9rCZPG3Yv5XPhTj
lMdEy62zpwlCUxauACxUCIrGU5PP/z0Ku183QsiG3llMJT6f/O85i2QA1j6drxqy9rHuWQZocWon
hSSND8HCq2muuDmyT8iiQLUfVne6V77qnlRN1SWQujhB6gSx9/DhsuMv4jw1B54Up7JPBj5hDEmF
8sDXjLMwTa9beM8i+lxFV+0qCxocUJky6ybaTmDkejHOznqpUMyETHKTAByST0AYupVBLUJ5a3im
mnYeTT7vo5+DnN0EoHPkLGpp7OXxl2jy4eKWug0sOxq9pRKKEw7vZzG7olNy3wOZ3RHK/DThUM0m
/7nVKr7ZT+laqDCo/t3XpobwBz7wF3SOZbtFUHFP3V1JWGF3j46nJjKoA4vInMKItsZYz66cOyle
jRTCS6Cxt0eCe2ynTY14d6WM8eU5AslB4uCKhuqzVh6XBnS1KN1cKIhuj7ITZ27z2eaVBmJ7TPkf
JnV9xPVb1iyQ0TmrLLZqTG6r/cp5Yg9yrFEAxsmYLtOULA9G98zTll12zIhs9tDEeqt/3xiFe3+m
YSQ4xdWiZarxPgnYIN5Bby8TIE3t3tPrTNnH/LdeoHtASGnLCcRXI/rStQ1qmFGvE7T27b090vFz
BcpJ8nyUp3x43rXbdbxMhYDg9+wOgUm5nykxzYz7b+sH+7+q/bi4Ijeor8/7lMJSgeVQeS0ZZ5qZ
M97AZq7bCqo3gfbj6fTGZFTEc6dW8lckKyrm/ZSsdp0/otPJZd0IJ6aewhRoQ6HNWuXPpRiXXdCV
Rzg7kaj9ZZ/ockaw3lbLZlGMOWf+c4MvdgQZER3/16nKlKjhHdiFmaH+VGGOFm9pCk8aJnWuGhIg
g2gRS1jO7FgfqyQ4MW1OIIempxL81URpBMnKQ8uBgjf4OHcuwLOR6kpcIb4j1nPQNEvED5KXYA3b
HaEqrcWAx9GnI2dcgmWKluvOSkr9JLu8g4MVlFdVsuHSkuOMasdHoAFth901X09jE2mdmiLX1Og8
hz9psQiLK8GE43vGvS2HpNDQ2OAtR4tp6S1yEhtnvP9od8AlHVJHzJ/nl6OmXTXbyoZgob0PzF2Q
jX7Hj6it2L1JPMeMrlcrZV8Tn5f/kgIZ53H/46D0vwF+LyLswx27f4yC2Z35pE1F98ywv/4IBtPF
vS7qcwi+VC7DmCgPb7Eb23eVe4pwtxyfCe0DCHwMpn1X+EmW0Iq0PFRPY5lEWPF3eu6Yg74IyFpj
nMB0Q4p+1ULO7NRVKX2f51+gqEhPELRfUBLhqXn0f37YuhER2oe2kaGxxGuBko7Y7cjvep4dIX3u
FM3qy0cPSvpKJy8EnL2HqP/D/Eii+cyI9oe+bbSv1sJsITeUperdC+LxdaMUWgV5gc9476FfiOJ1
wp3HxiZoQ3oHu+wVtyq88TIczYJDJXM833npakLEcE/IeEbUo0+3AHI7fJv/wGm+NWCVzXGrh3X1
ucQE4F/I7FeYUlSvN7i2kEtIkrtM+gJP3KeDf/2LbZGHx9OprnpJaxgpA2aCfDQBdemegBM1SKvF
zPccvJBEsHev3/SkYyLnuYwlzmIAWsa8nrJfmbFAdqxL07eK4P3J5c6addTGxJDpmym8klEC2rX9
zLYFfvLmllpK+M2aZJ0+EYKwwKLcn4Gl06WT/kjk89Y/R6Y8Qb2mWP1+BL2+DNGVdluzy7SzxC3p
oQtqEqyMiVqPuYOLWFolL3X55Vk7MhsuBo404/YBE6yCqwAzJCI0UcsShhUGNt9hFrr8FeVW9ao2
PwZmM9lDQUmfdjJZF/h9Y3eY/q7gnNZywKp7pZUfpQ5L8mfILUh1xTpd5F/JUepM9BtqUORhFswL
m3eLFaxjsohi4Zz25IxvONv5Q9leZA/hVFy7XS0QGITGempfsnAA7uDKFcmXYu49j75b4PIfVvOB
JG8oRwWZB30cdDUkQrb1ZNEq5KxH0m4haiZ0PdoU4jHAjYCTF2HWwtDURg0OKCWBCDdMuaCMQwRc
9KG1BCcRQ5RQPSDHLcIOIV3yMePAfQsTpmm+eeSEOCbsTOo5w5Xq0NDD1cZMPTIF4Xi7a2Ynxv1O
7pnmXq3wh/4AzezxiehsaOLYJV1uyHFFV/ts6PiGaK9poqvzTQvVt480NMICRtzm405xdpUpFTEO
MUkCVC8cNld9OI12ruBmd6K2n6LP+9bU2f5EN23SaN7mOUHYzV9z/0rAx7AbO+jXz/2ZgF9nm3Yo
FORAFOAzu67I534GfM3BHSjXZRw/P9s6+zMj5wRmlgtvkoyIG6gndwGYAa6we5hXYpPEIAu5kgsQ
H+mur9hV5KHoHh9/wpBCz202o2gaNf8U1VGGIGIRCKJgn15Q6WmsYaEMCSq+lTwjztM+FbI7Smwg
6uNx9cWse0PcOVw0O4ryaxgdcc53R1JQ8p48+MtYPLzF0U8ilwm5T+t1hI0YJmjlN1mrdrmiQNOc
4/686Y6PEPWEj/1RMcAtN6A4vomiOYJjIVBNLbPt8m8YCIWSq4Eqh46plDNZ16PlJBODcBM0sIV5
axoJFwkAL5UlUikIAgHUYHn8ZXXVZk/yxX+0OK3WGKApEgvXW3Nw1FRPWG2pYSCCT59EdmWJI8D2
HyzJiCBupMXnVm6YSuB8dULcp7z5EX1AA/Ljg94kZG9kUFHFAtcKwpiqFmRxx9qKVtReXgOhK/eZ
1CWA738j7A0VihZYah8VReUS88GD1VIpdLptCqT2vCI4x6gid1+nAQPfQIVOi48F0RoBCY4q21np
AOu20qsewScS8sRElYzZpyY9pTLIdJKkrbOTweiV7SjlzuWR4Ymh1BGkzEW8fCMg3582PB1bq05r
PoKgCeDXbTvilAZ6Yub6TYecROR7uVuL8/RlbNFTpOJZBS9kZulrlUYmnnlWF/bvkg91AQXquCHA
LtkpqS8s+JtyMsgeHg8m73JBFl4MmOayW9pymO/A6PTd2arxcTntJl7s1ekaTCsA4WtML86DOeMQ
8EXYvq5GuvM31U44A8a+U6N7oz5HNa2aNci9XxPNBcNQiWaWE3l+ZKV3Sf7LKDfh7y0nSzmMOLCg
lrhf7Z4VpN4eRZNXfWbKLpg4cVHUTuppi2YWQRONU6tpR6QXkNkaMlaTMHnFXD38hlVSqiMHhkrW
XEdmSn5yebuB63LK1slG7k7ptDJVu26SYEGViAwSBuEMWGDYzmLra6TyekXysUysFhTggb/5djKO
+jZkrxRSXuSPiBpzcxpCCQxooDlICw2R/Molt4V1xZcTPhTkkcCeFKbUOJLmZS87US/ZW+DcoO3Q
mGdxHzyC/A0cgmVUjN4OiQrjPv+B3K+qfxVCp48Xx/tffKEJyCIs7+hvn2JABnT5oQ5q5nmcso4n
HQME1a5c0UK2Bd3TuqAjb+AUQdzXM6qiRNtIigKX3Ar3kKhIoc3CO4PY0aJdDgTDL6ADM7T35FyU
+239CNntKbWc/KNZPoJ6e2S5XU+cI8KtqD6c/SF8oyf3CDBV7oiAaxR6o3Qm8PkemZVLrgYzFPj+
qRxTbZOohIYVjdQ5cawM9gBzLKNBPCBo9n4uPiPHXJg3NMop2aCqmfuTOjT8mbsRGZqRWAsXwArO
qz8zB7iu5PoGEQbY+IjJlSCkknFHCIxbeIO9sCKlLnfLfckeJEt4p8QqdUafuKOJjXdG+MARYEh5
lVUfrcDRvmgAUa/t6L6Qf0QLoT+ZiAXUmcn7EH3dPGd82rouROIwfVNXK/bd1Mr+rOPjB+iWwGyk
Avq+Ge2BNOwAuaGGAbYbHcup9pt+ETqjyjZBDaCkcgO6BS4eIkjZMUH46lIsiUXSIrwRt/xQhFdk
+qc+ZnC4dFqgCCOE8HRrJLFd5GZNrIKx7MbFMjw23xPcvzHaPQkmIYXc1XFqstaqTFKRJU10YvWG
+E8kvDiw/bGjBcm8wzvuyf7+yJ92oW4PXbiqQXgXeaoIV9aPiyU2FOfvlTwz6zW9YRaxT5SRxLRj
6l5sjlpB8ElnAGgId7+LdWdH4Iz7PUsOc7bpjIbo8vZlAcDGWFkE/+8OLa8zP1uvRZY7abN1ghk7
LTm9b8uk1zCUFKVuf4jmbxGvm3X4aHA1cYQRpCbqG+W1YzVj8ehuNvr+Z0WLiA9Ee2W5bMoMQFWn
YtzdeZeDaodIoj58oyEYph82wMbegdcS8o5nBVpFytvUfDAT+nGMPhMDu8zxCwir7jfs5prGtIB8
661W2EEqujbAKtt2I+2rBtz3J9XHjz4ACHKYLFdgnKQxEHR0Fe4KULvhagR5PGfaNo1Ae6/yFL6D
W+E66BjSWtVYfOfhMcRbtD/X9id3hB6TmuEpSYv1XzUFJTmiYD0fapZIlk0xoJJ55QgeFeFmwwKN
3aITxcYYGrNdPKc+1oyB2x2TsZl3qibleGKCm6VfoFdW7WgIBQnCi3C9FyeOTfiBd31oxYRPKRfk
LPq6fLd67/jTKjxJg9ZO0Fy2vwl7gcfIKclEjCj8hqt6g6b96sTeMMVF6SOPFTQM1HCUhPCsTqR6
BxuIX6aGE4A1L0Qo/7PRwI7umwRBe+XyipcyxBTGzcaMUGuGdyrbgXNF7NPdFzuAYouilq0ulCcv
3UnFUi+gB1FiHnpWrOjcrqbJlMsXI+15NIKKjk+eNBd/Iy3xiwDhh3KrWo6u5pH4zpd6XylKOz3M
LavCNKUBJbxxUz+7xnGyYP3vR5O4naNHBiZ7Jym0WScJ0QGVhI1xYuuNVEGXHnzPRnqA4xM/NPrk
D2Oeul0tIZHK5WgE4vU9MgkQXbqQAQZL0mnYwYskIp0HWYZ9VtrJ627HhWt7p/EWYaIWLnqV+++H
X53VOO6vNBFZt4uM0R0Dhcck1yDpS+CgWi1l1aePUuTjS3b0t4Ej4FWwla9BMbNVF1orcuhw6xwk
5PObB87XHY7TDjOxCDLfWwPRdmODc8L/ncrgHCy7zwFL3TRjJRJf8bOO4fuXBHDm6xiPR7PkXneG
lzwphLFgVFkn2mXlU9WoGRITrDzgKl/Q3EV/LCpcErzmWq/DbaueloXljKnySKUi/JGi8SaNolTE
4RGAWRtZg0dKZk3TamlHmuO0lo0L0QHbj67XK5bTKrV7EA4Z7Ris8JegY05JqdQl6mrDkZDkou9c
0NZG5KnUZIQcDmQ2lUXXMoHd1Hh+yXgfTAGFXrePhSo2jI+TJK+rDSqThPWoA77qENAnvm0M+fbi
cfzIBtaW/QBHJJ51znqFiIqnuLxXSYCJAjJg7vTdkU7LhrAVL2dlUxgJbX1IlgV07IIkYUjuI0SA
d4iWcNunMeVzEzfjXFVM9/6nMlfdLcFvsmX3ixMBSmpmGIa83vjT+qUDc3e24+E1RBqBbed/96yB
xBjs4le7cqJ7RCdm2fWseEDzRa0mKmRQpynZuJx3IpCTVjLvfKRbCyrK1ARboSZ860C5LXRplU1G
Aa+uNtHZbSGsFNyK3rbVXnw+XbnLF/vkn/Q1gQMDYVMs4Kebt2ga0WVsWU2i+JGgcviTtJq98XLh
KyMoxbdb31fcvk8VrmRfWDAxmy6wJ9F4g4OBlrKPc5oCZ3rFzbUkbEBrW1uEgDEgz+KPJJSu6GaL
Y2vjh9JLdMlmjgpt1Ayz1iiUVQi6K8iZcPlYXRU/rYoYLE8yqEHsBQrBHL+qntE3qEaRL2g+JV3Q
JT6Je50pw2G3igTJr8e9rK5OJ2kquZ/ikUj8l3TM2Hl4JQMN8Q0H56SmkTS5V4Vbdz9/jc5GSRvy
f1AGVSiQ+CbJCceRCuWtKR1eamsNBc5rjIj3GWhti0h6C3gNJhWuOJKc5/88uhx0sqdUMyFgu+Wn
MzHBsJIl8iGjIfIqVKyh2nKbpc0jLM9iVWy2wks4mR0gAqTu4AZ0WuWYWXTM9B/kmghYp3IWMi0L
4gGqNKjXBfM9spkf7HYYD3feAo+d50ZFjMn6Frs5m7nmcm3Tc0QI1HuEZ0gpuea5OHm77FzZBpZX
z36JUh0XUPr9DRjpyeuJm/ZnoSRW/Q2H8KyfAp4lIr9ujEP1Fsst42sa0fuppInSQUSXzNZw4E41
h1eW9/8q+AJx5E4iUeYxnF9BAsI7H6CgXADBV8QYHqCOI2/XaGtjNTkvtoQrtTR7Gc5zXGRm0qum
OZxrm2pfsPDI62tECMdWTl29f1gLVnnVU4yXg5boC9CgAT4v4gduZKLJaeJbYpeJjHt3fZ9zo+3r
ge6JUOR9GXKaBdmItZA0cnPbdSKpeqcMQZBjgXWnLYiErWItjVmp28ENA67bhlLImlRtEXw9DnML
U5Qbv6Dok9jRE77LwstXHpb+sMhOcBHw/wsVW33NHzznPNimK2LwQAy+AmyZv4v/vc5SN4h8LJp2
WphyLVIs0qi3O0zH2bw+KbUVXPGnlesyCl4eLRDwTWnXZV1WdsPtZDTb8ytuLVAZeuEc9BJGfeXZ
zKSC5acPDdpOYJACO4pHYN5KLx6snSQ6M+Niv72bE6z3DKRhHmlE+nNmtiRRqXbTFOGmievQjwAB
pD7eF7S4uxHSVMOxS+S14dp3EV2kTzMCfM5z1NC14svEhyHEMb+KOXlQkyxqO28ZTn+caW2fGi2b
M/0rf05MEFsDHE52qd+2NycvFWOokmEXmpg58vpHho7KwfDRTSirFdDXYYlbsJta4fqim3F3PYhY
FOfKk3VsGrafUS4gSIBuR7/MQIuMy0J9lDy2G4Qv3pF1Hx80vMPmMNbS1Gi5WrJePHP3SIsgFVkS
UZ7ATnoGzuBuDxardPYEvuQgS7deoH/N8TotEkkAERSKpRVoy1o5B2n2f8L1lpJSIzNU5ssNTiig
MQb3ZYpzV3BX/j+uDKA8fAUpbH6QTOAPG6kI8SU//4DCHpFfmjJhTE02BF0ga+DYf9g+dGbnoAEc
npNV9QYApGTkQHOLM8aeE3efYd4bP9LHd0zr+4qdzKb4r9K18lGl9C1T9OzxbAByNWL09qrPOuV0
sAFnXGyDF6Rq916+WHp1cV5CYPVeRGKzh5nCyh7aKzU07y+Z/479N7TXUrfzOqE14uRfavjCh+j6
QjrVAVj2GPtMkb66ZaeDMc1NEDIHnEbbBeoI0jio9SyMXxod4n05xoM5e1zlnzM7sx8/rCGnjqyM
EUej/msoNxG9VPOqOxqoz2B8SGjScs5j6GBrSAo14bkMbyb5spRyjqJa7y8O+ACD5RczdYqoQ4/U
dvvuoxaqmTIpMkJo5vE4oVv7aNAOWeMDbMR7Sq+jay7gBADO+kL4JXQRbLWQ47doBLkIhnH5Xkcl
mcft/BGEbrmizoDNgEvI/cgCuXKET/3Rhsh2ZLuDOK6yDzlL8kma/luLs59k+zUlPqqsnCWO0I7r
VCAjME4C1ihiQBd6w7H4BE1nQKgn8EbuTXl+Bqm5PsxxwdV7AhIVJHb+gSLgwNvHq40ExTMouMCh
5Uwphe3jK47z9TgDkY0Y9/HxXEjZlrAshFg4Q4Fx44FdgBqPn7ZkX7GapdyhH4iak7KbWTce4T+7
EqveZEtP1werRy2tUDwFz45bTN4J+rVw+dLUkXp+2UzC/smT/iUv9WL2dPHsX3BgQfOnDSa0kOun
jhKvFAUl7MTYGspifV67kPWYaInOKnHPI1ylUGpa9dXck4Fvd7UbYXj2HGHPgpCAq9SxGQw4qrr4
5HuNiIaJyQ2cIbD0TkoG+o3rdGwBBYJPkqRW+6MOgUmfncorVqdVQz9iBtIRu+ph3Yd6A5vINU/z
dOkCk6dAPgJDIeGLbhOt2n8iOhp1oSzIEhfw9+KTH3ng78jVDXKwzlgSnrD0g4izscRH9fQUvjvl
xeT39x/BqCiPDd4XOsHX2mSTJCLTqkjPeF9CthqCHRW/z9kvbG/kvmPcBP0ikfRRrLYl+yvZOufO
fsZlP3e3fa4/FLRG0TRVyRW88n4zgoOAaWGtDPzDyY0TGq4+2HxYfWosQdyetjH/kSJjsnmbaeLY
T4wLXXQbhWUyjXvAuketIWFf4as1zlaqApV8nLF/c8Teu18J2ENT0D63/sKa8X4teW96uISqxvtB
KvArOMvI/lo4RAVOPWzYZOoVzCSKfzU/wlxWcWBEqYo1TokukrITm0Sb6gI2dERjyymO3y897f6/
y1x3Eo8rmgd/YlFqD698YHQlFYrkJJi4xnWXzo5jUR80IZ2+4ZXGR1bgLNx5zquNT+snRnUjYrX9
enAc8OcsPO0mY1QehcD46+HGN/kZZJXiDKtoWYSd79usw5YgT0rAJrGwceZdcsCYdjV211jX65xV
IEwavT8Sd4ercumvMyUcHesmqc+vcHQlGf9D+df6uBHAoniAz1qECFzOfaBwxAMGB/z8HckSVPRM
nUwos2Q3D+xrH46Geqk2AR3aQhfHl353/a95daj6gvy7h7hkO4vRzN4WbscGPPt4wMzBbyA1a4zL
tQxrNYYkO3ZwcnwEhzJLmwBON/gWxwySpxquq+t2TnRujeOl+rSZlXkiI4bw74L1zgJZyqeKtaJ+
SPo5wQ4uF78pgNpKuKtKmL9ZeAzgj/EGAj0YGazL1ThVwVvHj5etdoPUOioXulCWD/FsaH2nKuAF
RZbZydL2qCCZYPcEmg8Wg3wq/j99jNfYNW3kh0MvUBXEnVEyEzJ2pQ+LFssirsaNsdUL/eSW8CvQ
dV/lWJkdzDQugzVO4tsrOWcexjDsUK7uQgfMTQi6RqylwHRpLCmC2Joska3MN/0hAWIf0vK+AtRB
cg5BeY4Sh3f83BHunvSX7BALRhCQGWfoNSp5J4yB7KC5UJQtcKSVlQAOOglrE/9MuJ9SfPQJwfdK
zESUsN3Tq/YvHRPkWsXMgFoeP4U2vT3TnS/hLRne3eOD2BaSqRZruLXEFujAZuVCbk6SPuEN2Pn+
7/diWwk0IZKEhR9PEGSyPYfqMfPC1Sk+H1Q6eXgex5C5WoOUs7apTKQqGUeqICXOjTmhIUGtZoOa
Cx3aGHhmCWmDPiDnJW9xqx2TubrrTB0uFe0Ti8LumvtVptuN/nX86ewuNSvB5k9PLuYFSu9XPtSM
PI+72oOh8Sr6zWR8XrFnkguCsZ8FYB/fm8KAL88JsP3zQEl1ffXHFAGaFYgIXJwuHPthVlZkt0YN
trzexVpHaJhvV5O4bcsEoOTFEe63bhgvSbYnCobxCC81MqiQV+azI7CVZ1z4hs9U5Z/ZJ8F++Q2P
Ikm6F82vfMvtU7y1JvIOGZY7glWvqkA61L56RSgeRlhx+nNCNv/6qSd9YM08JBl/BjSJdiuOfOai
xGlD4NYPY9lwMj+Kdxh7lGKEHo2Cg1ld23G1l9uS+Vl5qTLLawr/e1H4Y4vi6nTokfgeVgHCrYon
3zNbb1agU0mWMubvwakGjW1GsKsT/ZYqaSGDjvvdp0huFR/rK/xfArmu58BL2/7zXuL+ajw3RvFj
PP0AsZzq5Awc7/NoJ98IHegaqhq8TYX5cE3UYkMplQjRzzZFFnjecXBxL1egNTFuktW2USl+uTKU
6sFSjBpQTtL85S6Gu1GoabHfXMH1RGj9R16acjoBh3zhKGFgST3/h/P63zYDP2zLDQDYa7N1suPF
1yBrSUjwvO0MQNFiHN/5p8gA+/ho+Du/iNpq9ArSdwi3JBoMRqlVq5xFS3YQxO0lRb5vxzHlW1m3
MQAE/wUAAuWZA301UdJ2wUZYOAb2mGZVZL+3/yk2rtPQYsywEkDMfkY9mdqtycX65iAbtdF56IOa
mafK5DDJwnMxXVNH+O43hUjRG7H9NtUiC45xKmawwf3lsCUDlZDeVNEDwMkatVA0ME5wiFuIWF92
8nNzYM+o/tdPriN/A37h2ceW+nokSzarZMjKGtGgg8rHliJBcfvWBzAiPIlfZKwxYur4S5pScxIu
On2VgNF0qN+v+xfRLIVz+aScMJLTQjUFQImb3Pkg5Yq+VZ+Ty9/K93d+KfrSi4ihNuYvPAYjC4qM
xvDxfFCLULRVIs44Zq6KWnCGfzftHI6d0Db5xYoSCgzQw/EAd3eD4AV7RjtrtOgiZzttxm6vy4bD
an1Qj3gwyqFuBgDDjDZpJXP4ROQqwFYjKb7f0LUjlMkLiHALlD5nvcBvggt1ThLGOzFn48917PA3
lNGRzCmnuOSqD/WZCbW2MSxgidQMKo6WZLEuO9QFCHaISz2XvQv1t1f+LElOjC3Fb6yS++JRTqSZ
gWOW70dRZVVfUTfcxoYBZurly8UuYipAkuz/iNzscDjLqomYjAm2/jd9cT4f7pWylz+hT7o9ZOAC
u1Co8lxyA9I26YLQa6fvErZ9KEl897FL4suG4Sy11m3GhvYLiFf7btC+R+kiw3jBCXsS+aD4lzTr
HD5L9qO0BIDiaRgrfE3J+6lxedLpnH4duZ27y+SotFtQO34cVjypH0WwEfijBp4DxbM/wySb0QbT
wgYoDQ9AJx7bB872Nm2le9YXbTHGFeq2/XNJ1Cu3faf9pcliXSEDDome5C4ViZRztD/4Uy77Xjz+
bM6+NkBgSs0k5teNvw+dD2RFsoP2C+DdKZzTMaLw98YY8apvXcdc/hPja2+nkCei5/IF7H9sRQd0
jsulg7yLaBz5SZNqHXocGAZPko58afVHnZJfWU8U6lFpso/yFc6ezMLcF5GdyYC87M4vBYvQBDIr
1i0fwWQAJFHnOQhcXekdYSyOdNqqx8PTLDq5AZKIZgLn+1kN4Mr3ycnNfgpp9Yi1GOELQ3MsfP3u
+ceqKFtcyRAtfQtfHXsOqhUr9qG/b8gBG0ILq11TslvmH1h/Vv6t8FbRSmKQSYR1YAvOp5xFEBle
afZmg1DPkt4FesHCFy++95TJUWt5JAaByiZCrLChCLt/nmdPwWbugTqGqVSvuC0kX8qFanwHz56/
Z/g38fQTxnfz+g9cjgKbsoCGFDojh+PeEHWEzZW7s9xoE67eayKSXXo9/zAKiFR80+D/2u/DJusL
50jlpKV+NDydau/uenb6yUANKjoFqtUeFKQ5uAfSQ9IVL4lLPrfFZWnUOZv3CcCknx3XvKqhl5US
ewCoax7gGI099/ev+zn4TQprJc5hUvBTw0gb9i2/V1H9RMNZkYGWht/ciqTOAFwdZjVtyagKWnTA
EZH66eO8VVJV9Wgj0roPw4vp+NLYrBmdpdg1btdPGJ2OxnGsgycm9IraU0Nl4tI2f7FuCNrqCA7g
KCRgd8r7PFhEUumKNLOWEFGnXxs3S6XpugKW4bbn1gbK/6ZG3oJRs1JxfOVMGdwUStI16Xhocrwd
nMC+5YVYccVgvFYRx6oEAVCxFTavlXBHs6DXFleIfSewB6FtkI+z8yHjl4O/vqs8d+F9wjyqCpF8
nEdS9P1V8tSzbdFozQojbDGFTWwZhjZXPtWVsb7EnHDs2e6c+bSTrnTWSuyeaqKV9tPUJWkQCZLl
O2V5eOJ2EqWCzFrUmM4zuPdf/9GDI2VKJNTB1WYcuMC3uVx2N0s2dJgjBatx1ubJJQkN6stmhEyh
GTrwT8AFowd8TGp4I8mExgJrGknnEDD6MMNQCeyyNTMazpvzUGd8Ge+VBagzoWlV0dAFXBVrRFga
IKXD5eFt3fPpKX8y7o8quxO6KabgaNeHVFkKBgUCe6kYXG8kF/+5pBh+MIeNe1Bnw2ckb8uHnokx
i/vul3fZDpKsd3kXR70cKlIDTyH03EFznkYxyvXwwf3XPo3S+MLt2O3YlSylJW3fY58T11ksAIpH
9J+MiUA2RxV3WPDZ4VXAazt69IkrOSIeH4LkzAg7NLh9FWPG+QaKFasP2w8+Hp3EO025v35188F+
T9zjewGf5U2acYM/w7jXXY7WzRlHjwkMCfownuW1xRcT7EsBgeMdJ1mSQAFVN3nL7fHJ26obIKJP
WDZ3eqOKb/BBsLiVHnvn5l+Pj8kLbNADBiAiNwe6uinDMVRQOkfsDfL2WjkptmjeT1gorYw31+Yq
XfZGj0h3TFftz7Sk2S7tFNCcw+RHU1zVHs5cVYVAT15h8f48fZiFpipMMW8Z4Oadec70kycJPhKx
6kbHgyGYdGEw1PDVpGzYz2HZwDXfGZecu58KezCLn/bEak1A49uODgXROYyTnkm+M/SxZUcVyfZm
sdNsdQEsAf9g3C1AQhwsiOTFHLa4iw6HWr9GLDcrW7N1vhTIWV/jO+sYFAltgXREm79qyH/GBnrC
1SZQGxGHCG1Zi5jughicY4y+z8OLq+U1IPrDgqwScVHPtinaZ8talT/NnQI7wM3O9YdYTQF0zjde
gVD5QIlUcpsBIZRBO8qvdYJgDS/60HTtNSTxdVBdpwPycC262cdOdMuT/BH0VXltGZ99dfscbBj8
HhnRC2vGwPCKmJz5t1SGU/QSnPlFlt7uAkJkOkPeOGmn/sDmGmcJGssp3/nWx4VEWLtKrIGVyy74
kIzwc/LiQ9+ISWeUHptjvJxJqIf/Ir7/r8FocE2MubfMGDRulT0VzpV1UCAKqQbZ460Aqy8x/hXR
OL5GDsNM0AP/lf2rGCBHZXVGcF5So1M9BKoJl6SuJa1m2s5xtezmncwLEUKwbz7atM/vmNIlSihs
SD/8k6rS4WAitc07epuqLyEh0fOqZMNHmT4edtzR1ORHAZH2ejxbDnQ034I5DoyLDJathwkpn0HX
ZJOuCADRv9fv19GOahAfmdkWRf0/I10ctN167nVZu5rpkyhnjHxPYJo1zhPJFLYWTu0DU97b1Rw3
Gci/dn/f8kDbElYGillFZ5lrmG8jxfrVTu3iw2XEIOrLnennTecSCpKGIWTGPqJCRCrb7zfQdzW3
UZYZ/Q+4/1LC6SzUo3AJH98sJCaSSud8sx4XYSBgdStLoVf+Lvra617mmxWJ6ot3fFZxbF1qFHAD
2DUnuD7Tf2QRJqemolBOAjUIMF4aXzuLYteoSEgr9MybiQNHkDlTo8KyBSrvLIu6zYTcQmtOkQYO
DCoCtTTtXGwFEAwXpBgvB3F5CCF0l4v5UNdXxACfM+0g04pgaFwYwvrENFn5K3B2N0/HRpitT/P7
lF7pgxNs5RpMrVI0cAnVweAT11j2vi+CNzCAg4EhkszOaaBKT9SzK0CQhAXwpDoRsACz5RJRupfu
rKOh0Q2+59OZ5ZoMKXQrQBlHOPmTyxzCVmAL1lDXwkPf8vQK5l9TH2yq5cHlwbL65L/w/Iegypl6
MTEa4QDXtK3YITUwHSt/NmUjTxhOCKiHyX+II/SjaZrw2wsQKB1vhyGuz80AZnUlYVqIK/Kl9iDM
Dt3/KWT88Lh5km3wmjJY24pStaI0nh/FXTRMgPffNZB+ZGu7blYKvaUnWsNyI1utmKG8SX92bbtx
NuE4CkLDjI7TppS92419xlbuzdL9rhDruGWFvY6NTs7FdsqwihRsj6nf7clrFWUybIzLYOFd18iB
zlNrd6FslD1Mz1pUAFO8lhRrDpZHoRoxpUhImtGFPuAhZz39WbKALlq97VrLddkrtuBG9vMsphY4
E8ozLlF6d9o0H906hwMky5q1GC+becvJs5OBwEBBloqU4QayiyV4i09yspcBs0YFOSMmYkDdAuOK
qe5jEFcuZyK+F/l+TT+qd83gAoi7M/Lh1HPFqsbsaIH0is6d04fVXqLiJvfS4qU5yo8NrKtyHhDX
XjxQN9RyLUxYCjVZCR3mNaqsYuVYrn9yt/qX7MnrgpAiwHn1aoq6xzvU0Qty374zy01O4XrmiDue
xbJ5fx5E+kukCc7czwyG8HQMNXFNZKgvLmEi0Tv5ND2WWRr7yg2OTPhYPPktQ1rw2E1v0vHX7Sj+
oUgABnWaPfdehzK5KICAfQ/SQPjXr4XCYQsfcCoXXS84TIHr24ChuYxzUcTcnIqk3NFieuFTu4s8
0E/rh7jl9mTyo11MNoLdiViKg6uRvpmcCObhwZ98b5ZscIxgMufy3IeWz1Iii75CXc8XSs/YZPSV
nmGymuL5bXd3VKMmHeGmt1izRxqqO0ZqZoUMnyLQ7oLAWuLPDbl3FRI30CaS1hvL+x01pRFta5Xa
axjNgVMWbRY/a1ZH7X7QcHDWKScbgT8B60+WOC86BbF0neEfd0xupOH3tAvRIsRkF2wiJERMsoIg
5K3GJoJOsYC8h0AEzGdxqv+vjy1c61vPcPIbhO5gA+QQgXY010PkGSbO5Wvf9PWtV99SporllI/Z
k9V+UEfrrBvNrzlbrP9MrRzbzMciBgDldYhethRfH+7B8NXT0508eGMCrNygpLEwBbg6DULPFy/t
OHa7eo3oTNBmOi6HNqT7LngkY9moyjAE4fn7AbW8iLa7wTTPR7dqiGREaMiu9MWXwRsDl7xSx4A9
7DkjcbxfsvuyHGBXHx0e4/fTKAYgGx1TAd3b+Zq6aFfZ8I+kOpPUza13RUanWpotu2Rw/sltGGpq
tfeE6Fo5OEFXY8rR3s1Lp0FkaVU9gTjIfRlEekGSdqdgJOh3ld4pi15qMsuQ94X3/9z82u8Dubq0
kreV7S64GEzQwu4zs5OST+j1ThFxJMTCXLmEZva0/KL2pjkgRfRIXJLrJ8kPu3BnEekC9+B97PEx
tVxfGeZuCZILhOGzM92glOEgrolNl29cufpnH81978HM/FcJ+7AbXdE+zskB14kPU1p1Kmd/jxrE
cQJbzw3CW6f9MdmchFf/C5xbo8Ai3q7GiARODtp7H3vnO2MZ8/oBp0pWgOs8HeiFES8tle7rcQSB
MNnhL+WEISkt62wxNL+L6Xg6IWz+1pPepy+lvCqWJQDeptur+iSUgb3g9c/nFB0R9bXbKH6UVL+d
LJmeb02IbSABg/GENk28fFvFtLh5+iUGVbrkT2p2LSumSy1PSj6lUtwcpx1j5jfy1UJt/N9rbF/k
d7dua4y/PyOiquw63qjsTjE6p3VhQn6zHzbPP29pxZmrZp86ndg7Gt5RyNZgk45izcwjIVbMuau+
6tClaaT2eeSOHcvDnzD8svUgQ+Oiu4pwgvwVAZ+QpgcLL/A0WJ/7phK42f+vi3yA+aWuLTslNMiA
2XwxhosV7wsiLof9vd1k7Rl3QQa4jxFIMrUFFMpNJdPCDr6gFZeDz4y2+xYsboJL7tcC3vwVJBa6
IwAU11CopwX3B9JpwqWaUvIMEJre06lWSDPR7n9kqMimENrTNkVUMbmDu5IZ7rvTCqZd0beVrnad
RCDqsjJ++3Jfkw+brsDhJ4h1ISfXH1OXSgVZIwpVg1oQbanLqNplB660bmAPbCeh52Mlrm2KN5/M
NV9KWM9Qu4k5ez+OSSsIQqTa39W6HpG5sd8eU9Oq9ycpJOM8tKiu4gMe9rG2Wv8qmT0VyG2BtwL0
VHt384FtcWARFlv+gUTQlVo7ybbxaVz1WWtPYgwoC7KgBylcUEHAlRM5JKINduylr4Ho1gsuIHkr
uS2gIoE16+Hd9ndjQXu49bhqm7TKh6YhEnmQNr4KXPJmV2u5ZWs5oFdT8t5Fx2LjXPz8dwMmYhSL
ULzCBocTrdQSmahFV3xaTRDbm+1JT1U0PKrs8C9MP+sKEL9jdVHCxyUUw+w+0xHruGZLZ4rSIwoX
0yYJbysPzmYnNCpvjyw3lzs/YLtJl+sriFpDMSd+eUROEGoZOMeXEZxUgIaBFv8lnXBZqwA1xv+m
G8z2+sYyKtM0PsijgrPh6mk+LAS5XXuavGaRQs87QTB+zTRD+IWYDYaTiArPlD8MZnEXg8muQx5a
PcX8/yWJ5NUd+dZdIILL1NlnLHux9i0lqsMmUGAINUAzRxRnoSYG4vQsF/hVi44r4FULJ5Zbx9Pk
+9hoKw20QG1xRJ+P7Jd1WvAwi4kek3XRt2qvf6NPXjQPPeSbUKwxruDPbNIi3pfvJTF+EjMTFVAb
PDBA4C74JpJhAtN+jCyVjFJ6MkTFAgdryoT548Ink8KtiPKT4M1f2nN4vfIy6FcUzmPuYO+ZcbYm
HFQic/D8B++osF04lA+qefPflPBtDvNuY1Zpb61A+3Xqf6WcPJNSg23piIWSwNflG8GlNq/H4P6x
+d6N+RUoec03YEaDVvoh+LCZmm6IWeJGz2VlGbwj89dQnmCQUYxIffW7VcbP9SSzrHiZ4ANg1oW5
p4N9J8C+h5REB2xLryestYlGiZ5xqS54u4/ov7aCCS5ez8cPUcl6VaHIc9zMeREz9XUWRH0UnoVe
zv+3xSNceWRU66ms4nKGxJNF8VU/Xf7OIF9YLkx/PragVK6XVDHB/H/6tbmIO1UqzfYAJlPfmCcP
yf7Kzp2WPJ8swtD4SRsMVt+S2tTvhoS9LHyq06NP/trQbPtdCw71shCSBoOHHOw1hCCqm0HG43J2
sSXK0aS+yKcQAJloqtLqEvZScDf3bHZM/UDPYVgA5eTLihLSrI0cH/ac+R9MsKG/wLvvD7mHcCQB
LwtwoOP7ukFIK4tFhbwtibduomHOvojKaEJIyivFvPyEgVD2M0HphsVbxoATkayYBtRy/aMSZpLz
wrhXu4tduSzDyj/HSFzqcP5HV9ysYxnRsZXuAcQzSQSFgjA2RmFlLF7gyvGFpo7KO6MoSwY/EWJF
UUhhsAtY2voYSiB5VENZlONaKEmjLL5qLMC2AGRIJvVdFrrW/lXBFBK0BnELvSI8+aGWYkVDaoRO
RqkHIzRFIaisvHQjb3veY5/rBg746SmHUaATidL4NY8B4ysJTwxtsVgc3T7MUFshbkHlQeih9LKd
xVAI3OIrkqa2+hMlj+6gYVUwuqB3w3kCMCOw7Bp9+/UPg8cqbiZgZskemuoQuNqcnVjfZ+exLlZn
WHLiJto6vZ149uk/w2z3msgYNC/tbBYoBeSi6EkX70TYCuLxcyCZM4K3QDTtlWYLCqb6KOxxaCpg
rBZbDmILtJ0XFyTI+Jda4cr2yGbPmWDjMSCs2fdYuU5hIVGkYHsRJWVtX+BzjZSxAPxMbA2k7YYA
OCYHqUk8DtljH5ZJvLWEwUbYqF1oKtAiIxdu4QjN4hFCz0xXw6KVZKlPNo5iHihM2WyyjAiXLOfM
C6DhOe5KD5YTzkhaa09NZ+n6tOc4avK7EM8lTfRhv7kta6LwF2mkqAQtav0UWi74g27tBbHsJIjE
iyIGeiSY11EP7E5bY1sWFtdCxPpe9mzjFjfbKazJd8344cPsqPyTj6ctxWAWLUYZbphjFQcqSoG6
qIbHvfJiEfG5SpOn/YwVp537f2Zi9uKnWGSGXAKinOK+GdB/g/pqprxzX6WP2TTTkuHtk7+33DcY
zvNypG1Gg/ra2CXmQ+u1HJcGptEkX5rDVihAuq0sJmomXhrEiQyckP5m/wvkqjd/3YWKyRFgF6h/
r3p0maokUrvA4nMBZH0f+E0KDjg2j8HsO0+2aWUTxjecIF5DGT9STFdwCMbEcMW4J15gxarJg03j
qK1CtAf5cGgktwVq8JOZDC0PqVGJImY9jjAE/qwQ1RoPtkz34TtEccWHUv1ZGIYnhUCDbVBfTIJ2
QynUdqVbBJycQRBJ8ARMeBxI47CjdCp4CnljaRHYskwpnqGoOUsKUH1Lr+LiqNgY/A5AaPlMkNVO
+lgCvF8dP5j+axZ8a5X1J7bOC35pr4jFgr+8+J4AHmqS8Kx8Ru3CXgXXhKUC4rV1igjqsM4XtJSC
HzLzNwdomj4I11AZrwVL+EYXzJwzwP39EwyKxnvEKTNQJVRxgvTvRLWPERi5RXEWwrcFDGhmJiNk
yvUJqwyQrCLhuQz8s1fUlMBNZWppVtwTm+UVHoA6HiPMEPPOQf5W5jtjkntmoZIfW0icueGtBS+r
gWJYN+m3PgBrJ0Jk7w5Ll5MqkLfObI2yDoK8CX90b0am7q/U85bX1jFriVu5jGc5901Ql2W1hCNa
ISwaN/tLizMxskvlNsgyNqXe/j5+NL4rd47d0o7XieZsyvhJu8m0YMRpcI3whFTDlCUJlviOYLnY
jNLNQIgJElTPIhq+mbI27tUlRj/961WY8hPmsmngV72wPZtKtp0ozykAr4y26hKrFNb/LIO1zBRc
nfPy6f4yU+zP1cFDVB3cAT1eoMrAJx+CdtGgkPLpuQKCD0a7dw09QUv/jgEe0JKpcA4qbGZvESVX
gTbwdx0fmmE+CWld+2JHFOEjOeQHqv2Iy62s8goX7sXZkHvfjfAcxIkb0wz7CIwHxGcdmzqMSlUn
4WSkZnIGgzIlioR+efhoFUMb6E+Zf9s63XB2rnhgKLFwXge/9kwettgivyqc2m/AfSiKCG8MjAPo
DLky0QR3V0sqPfuXom1XyIfBtqTG60bpZReZKxLmup8AJUdRxplgBN8QvxZVLlpf/P8Mzd2E/FH8
q0FqMWu71Ay/idJlbzNflEPCnOhY4CZqTVWglKJnm8DHOQKwWs2BD/58V4bq9yWCZU/qD66MdR7P
VucG9Hn7WZqUg0nzoDlfef2VS86tV6EjS/pHEiAbddLd7fXYXFWLVfEewD+D9yCuVkkIvrKBYse1
gcXSnOpi5wuJCfoc6BaMvSE2DJRPiuDjDiExyr80ULQDXCKVCsUknE24WgxerOzI8n0C88vDTXvr
v/blCi++yCtwFNYCwqFOQGQAfUDc7U7py5UVF0YBf649TyTN35YzrdU/Lco1hmQLdlT+W7LtqTf1
hUyDIKOgiriejv3uY62Yd/8KWFObqnlIFmPOlXiezwjuG/Lnx8ZTt1kpPZShdYRLX8+iRf3ZRrU5
3uN8j5JhGKKx3Wd/dVf0q6yUvYJL8FyHlXjcXq4NGr+tj0nNEn9urq9T2BA668kjMqdB5WJYf4nU
qb7WhNGoYU7BqozBJ0vuBdwsTrNUk/J4DEtnxxivSpTFQsfwuTJnXcOSMuBeCCjk/PtG3QOwkfqX
yKPXU96Z1k9NbFMcHMX90oYsVSlsIqurCrbxXXsgzf+r5VtZQ14mC1TsTH1Slr+WLj9rLHgJvVQ0
9irziEGOIekf8Mbw+ulA/5mI4ztyN5VlAOLIr4jnka0siraUoNMte6X715z4Y39aktTrqBXlcugr
xGkmx36FMe5wrjg2H01+eJm6iIydhZr2RWYGHLZjelx50SLNHrxITiTJVYxh83Kp6DLysYy3wRlm
QJKlVgwVGfgQGCyOA8O9y6At7Geem4TzPjd+krys4uDeFj05YES1zou6JRs3rQEpmQliFx3X/nMm
CHBO5bLCFg/WoquDoo3QoonjeRcDlnov78SX51wv+Ljj+l/hHNNLlepXzL4GoNkH7WGyzm8wSax2
GOBjorLpqMPfHwpreMX9uLu4pT5ZivW4BLXeshPx/r25N6Ib5QflWXnn0JnRRs2AkA3SouxMN6lU
iWYZ/ZX7xFTTq+xDvhpCzQpBW6rABICsfSwxrUhEiWAxHvrvsF7TT9b9nwHO3/eUODMjZi/Yduxt
Oz0akMGonPAam4K1fJlArDXcIgXFVxXhXuSpN1xUXIG3a9/BI1AXBg7ZHIjfZZZr0dP10QdsyfWb
9LQ9SJTJneJYPJPjMv70yuqdq8SLDG0PYSqP6IH/cl6bAJdObTvUPvGfW3LXg6tEJzHbvHNoqli/
n9eYEXm08ilwdc7GIvc81uG5Xu3EvNQh9vmayfNrI0/63t29Y0a36NDNxljGCsJcblTwKHgu9F+2
hkidQV5920XeKnJBjuLxUlELzQxGQ8TuvFlqD0xW0zZ+MfZ728fK+bIhualmxgmqeD1O44lweB5g
r/nk4iQBLKL7d7zFmzrS4MDBsKnX6oP4Xfz05t8elNKnncZxunH5OhbcjwycBPVDVdkHDxlRlgM1
xKioi1uUGMlVB8u7PB7b2Msx5iGDywA/U24ZTRQhLYMvZy1LGjuMj6mDfjAWWof3kj8E+hcd/oC5
Xbctu85t2x8gTXQPnIg8jImPHNHkSH5n1svV5Ue1ntd9uXCKpWoXEp+4GkTPFPAilZbZGhCr4xFK
Y2iE8lRjBSdV1Jhpm+8ebF91tkFw6SqhwDYCF4Y7Ji9MBM8iRsDBjBE2ngFnFSvvS/AZj/GYgmrB
KFGGK4/6Njl+qYvAzNU6UkFLl8S70fPx1FIcrbzU7tibfqeblv29SooeLmnTLu7VYPG2txpcGJqv
u7kihXEzNKio+W6DkD5ZDENSNWzOsPCSIs+cZxoBD3vUr6hH+VxqBOiaUTL392uldCqaDFBZMS+F
kVQQ5dP1kqnDP+YlJ/aE9gWJ6RnL1ngFMhl+pds8QOXjZ0cmJ0WShSwdmEjkn13OLoTfCVPtnTZi
vdKQOvhR6C3F3TTxDkWWMSAFLqGQDOSbi/kpSsEKnEvuiwxN5nJtq9IJMMzJ5Llgs6946ubHfePA
fEuaF6XiphghfllK2qzrTCHG68bSlmvowZDD9BNP2HM7+ImgGFKcpAMDog6Sgy4y58MYlBTR/+z+
SU9aMG1jtOMiyJghr0EGiBU4QjqETf4UcPzCAhNEW7cddnYhk7nAWjGL5I6As8Q0+rogGwM9Z+na
qFn5cRHsu1BFDfh+FhZY5dQPnN0l1mNoKmOsssjF89re/prCsojCdFNS8GEL/pG0p8SxnHHiwNet
X7LcS9Lfhmr6heHWRGfI6fn3tqtldmgF3/nnwoYZmtdo/WrabFqIgqZtH7GhdPVoJkccpI0PgVWf
Ou2uX5GvqgxB41xmaKJkf0qGugQZhfYDE2jv3kWP2wa5dkD+Fo5mSvTNk5LfXUdleE1heyhWcjcW
wcZ9BTDCzy/TYThSQAvwH+rKuWJV/BxEDI94XW+TesuOm9TsFNlk+sgPUVudgDcHauebEvBr87io
ciy1L9IqWfpV6BiDhfSK9zSIfDGy2Dq4O3NRalfJiYqPk7Vk8bCiPg9aYEsCjhXz19QnxlOWoObl
/zJu1xrwx3ugfExypJ3rW44MrTUyU7Y/SAz/KKQGp1r/0gTVzqEX5QJd+b2KoJdOgVNLl8MTeRFK
LzqkUmHDHnyCxR8jnJdI2/TyokwiAUh939zWlcYezNf6BYbpVDd/+OO6coXF/OoxvZlBJsZMA6Rt
gL0pD1jJbszRMNfT6NcjRduOQfKUj6FrPMn5MJ61tJqvQ4Jr6eEWb90CrdMdmyIrCqCs10/k4Dzn
bMbwm6MFHcliuGKSSqudHrmsGl0XzC+xkn1v2L1zHWRjg8cO2E0cHqyY9n7KdUpg+UCoQxoRRxt5
ulerPXkAINi2SHL6imUmH290mzOy7wWsOE/W6VenZ+IdL9hrcJTDrjdxYypuS2h2wvp5YPfSRfGq
AgqhecNAbqYchSVh0SPAjxsgNP3bYPskzNZ8ouGH6oxf4Pz+gxSSAn6KcXA5dmRbHV0QWuNWVe0o
zH8mbKy5aYUuUHxCYu3eAfgDHpds+Io/Lsv2CRu9mXtqQ5hLyeZfvXpAWQ7MfO8v3efwXybM00eG
S1pxEVDaMo+m0Z3V6pC0DK+HxkmmCkfBsEZvXyoPbZU9dG5iOpCrKoAsclWYV7BknCGnHo2AwQ0I
CEF+FHEoJsNPtGXmdUipC4QAIMsASJPjPiVw0hbTgnkFQwoU5T5NLOW0Dg/UNqovfndHkKRnByI+
JN1fq9jo9ealqHDGS1fXSe9v1ihJEcR6DCA+v+C12uiEu9JXXIUb9NnTgq8twv8w48HFNUQ9KjKu
wm1Ot8EY1uzgv4Ny2ecjoRkIEURxoHuh5rIBdE8dnGlBwT7NVWKci7Wup3zKwtjjim4sceKzGTWX
IxC0d73j9n15OV/bGLoB0XRGCGzAN9+Ocb9Xd+s0aDHmRmOBlA/6fcNASykcVWsFAdtwCl2+3BFa
j07MgoGxSxAAm5+G+D9UtRRf+rj2NP1zXbtr8rWEAsHDl16beS26GdJYYdKqEWDGA/80n7GpBNMw
Za9WDMhLuActC3O3V6gsA06mdCOaYtEumq3/Lb+zNSCw1sSRgtaNf4OhD5NhmhKt9ElHb+Fdd5P8
crFScNyrEwXnDhEec9XzH4m3s4shZMZsuGKvZwt6h0bLhMGSHhbACq3o2uhCQ/QSOtxtgpguHDA2
G0gJ9H5/DnV6a9rXKGZFOfMjcv4QnIIARQi28VCs0L8YvGZegaaYKcQ1iLDZkheSWslBT8MlmBX3
bZ8G0J1g1Aa9TKkhl7qEKrTm91+d1YleLjz4laPNpdYV+3dqpvG5NuOms8FKsIBUWZs+qdB8WAkP
e3IFFK0OmC+ltbgrTz8UumYhnlI5jubQ+/N/DbkPsvTXCVx0uVFAAUnEM1T5KiknIF55a0W37jez
Gti/hAgj0PKT633ExHnM1lOYx/4K3JGVoZQXeatz2xmaoHMNopbQD8RafbUYtp3ugfaKnMN97Uuz
N20ltZ7OT9YUzOlBTYFBmsdeqsfSnGnczMtBhf3Gw08J8RLq6dvll8i4/JE9BAtmU2gFFcycT3Eu
e0e/FbD7VKu4e4HafxT4wWh6B+F2f4dRH6VBx72SZuXVOkWQpWgfaQg9IXaP0Kaumj/Z/8XRh8GI
Tpdf+gfoUiHguMW9JRUcme2BFNr+MtvkFSpabMNqmI5/CwFQ1AfnurJ8w/vpDI0hY4GEFsjMv8Yy
aapuA/JuKgMpN4xbOu7/MLy5SIp7BFxPvOa5hGZSre8GhPO9QkxazKtv0SMCziwg0tLsA2YLyINY
FdqflF7ids1gaqXzICD/NSAc/AJxG6wvAaRlZsw69uTke/Ory8CMQ+6DMeuv2joubz1qhHZMQnQa
oE8ls8vsyQWM61urTpI5XABwT2EhbB4PtKuhx2che67eEoaXUf3K8Yt4aWc6inDN0zuYum96Frh/
tihzu6O+ZH/lBtwWGZe93H5odsnURyjo7vFMFX0rvWpOXh9vGBSDBGtOt4sqDwoxbrCA+X37u0Hn
V2T3ORBgCV51guxnzkGUsoVL6cgaZD13K0IbeOBMSzFNE8V+KCXRKZ4XR4+rrggB7OEfKXgt4k1t
Vdcw5ZM9ktnwxJUUkeZwPi5AJYKoQVWDn9ka6tMwNsx5/IVvlt1yYaP3zqrskI/QRIwEUH+pCRld
yii4PUc89hG6FRSzgcvwIN4l9EWoSvx0AVfpasKLUsGlRRGiDwPylJtXgqShHOnmD68l2EZ4DySC
WhIZSun00gmS4SuFgdnYS+jKOm6Oi2h73l73McS9dxK/CJAqqqHOxZNBCFa20kUDi3FFH8zJcrLl
HMY+S9PQcySoW7w/AIzZn6j/l5rew+VnL2FnQJoxAH8Pmh5YwsioAuSdjo6SM30qp6LQIj1BzvyN
IiR8Gclt2ZSU2SqQce5B6NoeJD3Pf38jvhbGeKvgscwzkUH+FGxNlXUVICLawJ+m3kWhYjTHevf1
DW1CvTrSaVao9Rd9aC0ek3Je1WT3cDsW0ioFLahI+7RXPrDh+DCp9OQR4lTVi9oY/5nxx1i7ZyJl
8U2scqDosgG21+4j65S0uxNMPSteDPSppXEDyvjAVQtoIlre25s99RJdI+/QdmeLkGtuVTTpcQKY
Hr6RC6o4FQIPyd9DZpe2DMPn7edJ6B9ozkx6G3DpiQh7s4Q6mGqEomrq241sjdgOoJSwWv5z0SB2
xVMFXPOZe/n168m1Ist+D0BTmHSQ1ruk5OSofcAbBGeMt6XY5hblpKq3XIeexse4ypQl6XcZei9e
srtXJ1sQTfM9Pwgf9lWZwTkJXb48f+HrrktWlFuPikKQ9xUCBDMuoLKJ9ISo++egBZx4ijYql5Qh
5jSItfgw0yFoUVCe2a44bfavT7m3tFpv9Ub4gv+Gx2CRebMGy0aqRRI0R5Wz+oHCqEd/gnnI2UuE
WMplrMdtjiISwWoD10QwmS3LNdvb0TWf9raD7CJbCfY4cipmSUkxfQr+Dc8M+6MIHdi/HSHn07v6
qEG0S01H/w5iX39RHMlJ4Qfyng1L0AOXdR7OGG+sot6Sn83rTU1KLlGQ+jZA0m+HTJBqVc6tplAU
+RpYiwpTtqx0iLf7r56aMqU7wIeQA+zHdkMlDa+v3VRwGOYGZBCj/6gIcjCO0PFaeOlwvdzUYytJ
LAv8ST3iHtCZq2Rmyu3Y4pyujXZYOO7HGOTDjidJjx/Abf450rOEhfEG8mWKgYBnBkFVitUdWV1J
g5u80C1eF9sR4QFlgY/CYvqhxO3PSdSR/nc7fNhdq4CKuH0srTi7FvjK36c/O92t1krtoa4uQpEO
bk+xtrhzPTD7425FwIyRR1WFncA6mRaDeggVYxigPZLpE7Cc4T0Vy371U4DGV2peP9S24rOySKa6
UTmlSeegCuUuVORGMCETQfdiCLbErlvdew9P1CpdaQ1xRCWTwPsoUXGaOeQZVKdGJO9/6/sbVLuq
g8DtdsMN62WqkTVrxP2a/mfzdesZI2u4UeqomFCmzrjbp/4mc8H9LGl0//ug28a4QidIUS8oHJU8
PfGw93fvxDE/xW4/JejLUcGQ/KfuqUMDNy4wIFbvZmQwadmkZdVB4f5YKLgaUsp1qTy/ziQU/fX2
JsvEblHFAe+ZgegVP39Jy+ZABqMeTeLcAFoajVx8taTlKs49E0dWls7X2nJzAg+1yjEYJy8KhWHO
/uXwAxxHc+Q5jTQnYZIT8jkAuEviT/ps89ADGBDwtLcBj+5NAQ0ZU6IzWP8ld3qdLsKUTxqq4bSM
PvKyna4pIkwiWcZrCjpuPO8BJBMEcnN0Z0DiYnje1tChdeUtcohVAV+V7lQt2q763dwIo7W2rcSW
AwegKfHeRld+ibj7KtKopgSzk8mKLw02zZKMCcGdmk8wkzj9gsggPxrYAYMIVz2o4bAbpwJaoe88
svW5s3D1LhdezVfs4wzXScMqLaapg+/ny6CqqAbXtNgcHMwnrVhcicZHezqpPwWHLF6W52imEBq+
/FRJqJv9eAJJ5zy+ZgUYaVTAztm8ZMjnq9WPGjExuHrCWRJLuegJ6UkOqzeOOvQnqSR0jbWJNUt5
QtHsEOkGh55wMs2kX8eR56ZKBWPePrMrM1Hz8WhI8+avo1/EgtoMosp0zNX4Hcd1RPJfrvJnf0jN
hpAhjiYO9pPPfChbIDJ6NHgDV65w4VPsu8mqZF+N3PwylHTRoOSTIbsF4SEi0DlxVjYdemA5HTX6
5yLKQDS2hFumTHqkLjvxVDccv1K9v33vwvUs9rlBWsrpgMdyuehVZAUSgqiQZ4zhvEKOYP1tN/b2
bnK55D82P/TEx0gAR/hSDP11MKpEGf1S/zCLxNff040VZXqJQCbY7rl2QgDWj5uunt55DoIt0lQ1
0EJ41b85fN8TLB+9AMzx4Rsx0wyjhl7SOOZSQoEplNZUB9ftXbhEsAgG+COk4XcGeBZcr4LDnNAM
vG6Bux9VbUvfCGdCeSEj7UJfZVqeI9cgRIbpl0AGuKL/xkYJTzQnAPAVFpc2STZTG6eav+pxW7ec
FS0LEN4P3rsVfz+OZFB+BU8kKLMym3BvZZoot1OAf3HT5yMzljO3nCZb2m/2BV9f55F/NOlQCEl2
FVPU45ZknTA9oLsDEqyBwhqwxXY3P7n5W6asKaFkMec563AodJXTXboPZyQKVtgNSNT+M+2EQwpk
qYt72L2n79syz8sBeX/LW8798taMvjtbx8J09gDHCuQNpLYNcH6XG1qPX6kmZl0cPIlqQtsgG6dz
YeaTTPpQBycB93hwusrJgcPpQzAzvJIHPV4wHCrRNBxftR/fnuu5pikytJSqOm+4s2Xtrg92H4ur
FlhAbcKNnwkGRsWfEnEsNxVL/fxFVUgCHxy5hE1EoPfqFTohyTSSQB+XngmhhGCriTHnjHbYEQOU
nL6/hPsyuseFdLuu+SwYgjJ6J0xRD+CGrg8UVlR1eBTKsBSeRYoTbTWD6SLImbJxjA7dwGH8C8Te
91TmcDlhbT+ZZI9IRvhbZD97L5zzjwiarU1DjTnSIWJu5xfkA2/toGlFsj/cYVFIb67Az68DkI62
pDVm5jo1RenbzbJZk5XkzbP5lLdq9QeJadmERpCs3XMxyE81QCVV4KPPwiPEiPb0KxxPgyIJwW4I
uD2PnoLgK3oI1u6/vVsJazSbGwQ+ofrLMKssLe+6EjDhqT7biOySlkFFOB8kVrFex3l8HfNZkZEA
tFHOKHxPCexY0ju4vE5JnNXb68qLsgzEouoq7VPDX6MBAs1Ueo30PoS5PfHLNkPJZuj7i6Hgmheg
tuRPyxeVqeYvFmLTvjq5u1Ki8usVHcsH8Vv3F+BOdjgBeRdgGvera+R//0W00xPSDFTjko/Bh7Yf
fJ82UZ+KeS7+X3YenuXel5b00yjdUpheiM5p0A2+VwIWPo6Fil3IKQmh4rINYScJs5DsozOsNZNq
VlnMn7cYUg/JkQG/IBjMHlFAoToEzEDLvt8n5ekVfwOy6TJgABUBkc48P6S1WdA7kPY6IXB8+6Nq
FSZTkyh/zCT6q+ZoRY9mBWRhba7EwM3Tu/QGPbJwliORoNFTTGnwHHGtjzn0rRhU08SoBZ0O2QLS
Z2/QC5J1OFhJ9abcB04aNNnNdvINaex8x3bnztUI/ip2ST7sRxSXBQ8Pp36PSIz0NWT2YzWsubB3
R+QMpfc2AE5Sze5LgoasyTF+Rr14PWrHLib/jMdzwDQR/pHzMLpvTlwLRvq4OYqSd5S6Y5uG0wDS
Sl0NhPzzlFfxII2EXbjUG0aFPeiWOIt55IkL3h1MPPy0LCD2GOyoSLFUUBLde/QDUVOeqk8EsOse
1kMjh2X6vC2vnUxJg9dibrIfOYWNNeJ+H5yiOn3r9rJD1AZUs+xxekVaTpo8YAy923dmm+LESy+n
a9eUm2WRp9uyagvcUVaECEgseVO8YcQ7ljz5mUSTLtk7AnOqBaTVarWApz0GZjv5wh6tF4PoH66G
2F5+fSO9E0OM+r63kfT6yMGAmB0zNJ7+0Ztf2nFZ00ZLhl5DU6TWzXWMq+VqOjJ1ZWLasWJknPxB
aK/7jAy+kq/g8PbbyqQski3f+MtLGTVP4og0vt+qmwi9PUQ9cfQM7rVVAXbFyIpLw1C6HIvqKp46
P8CJT3RM9TZEBfq9CLpqhZ+wvBnpwqcy9MZ1CHifiO68bMk+bgY+EhPIrhrngb/YKvIItRyF57B2
SrTV76lFo5tyLpGo7oLOBEpxkCTP99fEvFT5/EX8iYZFxfxI7Onfgiz1mEgK5Wna+ocgulrav4Re
KJTZ85K3+Y5rfNerLgwDEMzM/FMr8czMr0dXci88XaQjf3oX6LuFnS+O8dhQkvt/VGpB4mEwgN4r
K+rG3BgK45J+RvWnfi9B7dn2e5bWmDws5B+9ByWwE73AhFgKIQjhBlDQ5/bJoHtErjHyaf+hQ0Sf
Ol0eRt3t2Zhj/p8R7WwRdK83Sd2JqrjryRpUFA0h38qdQEzefsmm/Ac6ODxAjZosZgo7T5QM2ENo
rtTLsE00/alX6gdPKwNxW6fk6ntVqTRuB8++W3kWCGEY++UgAs0Y3qdQnrGBECBJrcDbEPm5BubL
Y4A7XCIG6leYEikjL/CrYvq6LJsj+2ciuiX2LA/5uVgDOXTTyU+n/SKu40QsetcEmdf8rEq+viKy
+hs2kSN0GrpqiXxVH/H0Yb6U1EgKocg1eSNAlQkf10AHCmuTAuq+dAHEZZMucefgLBfIv1We7UFl
F8qBej0kEXHkaLRxVbADswsnjFUNocpFtr8BOQEEhbosz0RGvyrub57P6uNaMzFKxsCaAqVTpLpN
LSO7EOAu2sVXqHJ1tEzuM7X85kV4RmN+MRNR0Ff2L+/BM0ddpygQPNz9o3cfrd7GF2q9Ct3cxlZu
drVt2Hg/ud9zwv4wLKuKtgbrr6pD6DQfojOqW+f9jTdIHp0zPSvvjFUhKAvh2ITwR3iJYZePG6VB
O6yuh66E4mp6lglrNhajOy0nGpiZv1IFsGH9DpySMRBbh1jtVo6woFrsm3blUMFtHrvcHKFXNydD
MvbM6aWUpjUB6GB3GEM+b35Wzztz2EJ/8Rpv8ycGozwXxrgHfcaMhIMoolrdbXcR3xyKx0DrrMEG
6qsMrRugbIidHDksh94eGWHbt4Y3xlG/QHJMsgnyw0mi+4PNs8zbmT/i7meseXOKMi4eIkgOwQMU
UurwrUxhcuvyHbx7KcXehuWoBM4XwYVTSikg3wzMrQXlTcS+W8ZWBmZRLfS6GXfkQxEygVyFtvPB
tDdETF41YwUgBNSj5auas0/nSYbBG8rWhEIzD7yqcNC2xHC7f0il+eDqLFooUDoe66MVLKF3FJBo
9O2a6ydnyUpsDeft/dI6SMVqaEP34lVRbtT9zslW48djUNbxlNTorhV9oKBZEHSiwfz9TgR22IwJ
5bOIeMu1PStlWC0G8W1WI9LLF2iyiN5yjimpgCevv+mXaLDanrDTk02ox3aJ4kq8Nl5mJHl0MXL9
IylPIfd3Sd32PIE7d7yorGnIHPsV/gdnwGLz4GSYwcDpIIzraW7O6bgTOqMJkwHHXykIOJ23YlQT
aLZf2bwG475I/pCZkigAIkdI0ZYIVnL7pcjsY1V+AE88knmZNmVPTgiiCHXfox9wiNfH0qQ7W6ad
5p980oi8q08JItLmx/rv+HqWR87yeCEepwLDlOB7q5vIYvtzPaq8SlVRkGIcFmU1HzN2GIrIowpL
hoQ+dBAhrzilhSQ35TFaNWjgVx/4aVF3O74ME2lAjpnsjdrArhpyydXEYmedieoVJV/EDU5+/tnS
hSFa594fjVJsmd5mBIv2CeUTVzn4OT2JjI5wyjACGFvQH55MHZp9TuWWPFOjwE5wwRTmK3P4W0IK
6K0ezk2ZL5FNOgzB6nYmZDyWMa+7m847inlTlKMrO5d64g2QdnAxUyPNYL0IeOKTkXIfgbdlU8p/
fLAAKMLAEgB6sNrrrVDtNGuMrAO7UWkJB4acvZtpOe6qLfmI1l+IJfxY85cKG0Yx1nz1N4RCYPPV
IY+xe6nSgcEbb64IQ2AJttP+mLQ1/5SfOWIVMFYV9Sueq56po9LVNovIGeflcRJpEF7PUxOADLbs
QcdXgW2dvB6PPcrWxQolU98zlnT+QCX2VzFbDjNgLDx1ieBRN3PCuI+VpFADCDsVzxQAg65O+lbN
ri+WlukqoQYHeiXdOXJwYSfuOgNjYz5soPV6mxmfjrtmTI0K90NnDWwArvevOEDn+hUlI1jXZqtW
/QOXreroZqUJ7BH/7wGnQiX9T9hUGcBe9OKfNqHVpzMX8h+IL0QHNd6Tri5KmUwB1VMoc6SZjSCu
tOkCtlss2umcyG84pwxexI3qkqRYEqVr62pQr9FHlrcICj2yCK5xqoi31PXhyPFPfk0jxexRGm3r
7URP9oYiGxxjZY98JAy4FZDME7URYO+/K1sPIWhO3dJLiR9EXDkFP1mm2hgntp6IgMTIvzx0FqN9
PVkaMIIAK7Hy7ub1vf4iGBLoUlpzNY6AOGXcIE7A8bupf0bZOgS05U2TDohWL0eXzupgrnon+/Og
HdlYDM4fhEPSFx2+GpcLhTFPS2A2XmBqNc+eLUGCFx8XgRcQ20VH9pGdHMQQ1bmXASloa//0xHgA
QhprrFBXPe7V18qI1bjlz1CWZTOPX4cl0UJMM31/8Fjev1B9EzgQxcu5qC7eEOAPLaQsTnhVb+I7
oob46vA5lWlQfhidXjR2Nw+XyhE3F9RH44LxZz6eMUOiUFqgsye3WqKmECqagebjw3bs3rbXTme4
r0byxtI5jwNy5ZlEKqoUPv7keJTqslhM/VJ2z94kB0S9EvYh5F8NtwdGodA+vONwoj6jhTdGa3u/
qgiYo9UM+1lkA2iZYDe49J9rou1HtT6mM9Udps87X6sYRRerqlrZJIUSWrmJQP2RDxSKS7x7ADfr
r/A4F8tZACzGQSj9t5UdEjB08iVMG9gHZFmaY7D5m8paf001zZEb44VHKAvLf5XzhE86PKIIO2+g
ipJPtz1qMHLD8QadhiKwyJQTj2LH3iDvZvqU3tUXv3Zt4tru0VeKZxb5Eo5UCUXQ4oeRaPuxKb3C
76wEX5k6YiVRKd24y/XKO3cLQulDWevaXz6TUCqNyf/4x4uHBKuO37lVFJhBaFB8LQVh04CVFYMU
B7doqZcLRL2Vts1fP5ZkouSk+gMexDJ1UBiFkEztBxwKtkKRPcne92e/hI8JJt3dJX3/sS19rBce
oHH6XAZMspIw3axaiiR7ghcd/LVQYdW5p0RqPuFwSBXKZ7rUTWet1SI/+J1z5PDiRRdCzelYQn+6
2XziHG3iZ3T1liybzF12ruCwWwje2lIIU3HJAfXAxf6lJyNgDcxh1rIFVFggz2cnvv6db9Av2H5w
aCAd+a8qcfCNQkVSfrx9qqhsuyclaKWAJg3OmUng4YGky5T4vrkTR5RSnO6Ob13sw8LgGhcjKlMe
n/40I4gxzs9pZgDY0vKEAQ2iqsO+I9mWQm7jCnxM1o+w0vcZ1hxlwY82/XJM/7bdzx4PRAj2E6R/
xvUwstqG5RcfXx6Z1UmGlyjj7N9ONS1Qcrl69EyRQRxvuDv4FOXFO7xodkDtpEPjPNq1SOGvnWvS
IeVgU8NHhy/7aBnk+rvU8KqjTINTTwIIAN5v8HDlvIrzoOKMBHif6fVVqRJR2W+UBARhyyuKd6q7
tucc5a9YCnlP6qI8I3rjkoKCbuK6Sxp8/vEyAsjjWc7fTKo+LrBC5MHDSF+0L1CAhky1FK4O7LSl
YUkw2gclXjGXltfKT3n++tYcmKwnxVprsRjCywa+oDrv7uFQA2C8PYr/fZ4twWtzkfT7KZ8u1PL+
UOhc5jsUAtOOc31/KQiSVVqIv/959KWoGYNiKXnduYELcNT1lV6muS+M6OCAS2pPZlRhu9EfZ1mC
JYOoNJ1fIE7zm/p8j7MCX0QrrVMvuEFGF2HVfeHn0+5w0swuYqSy36svqp8A9OMsLc0/jVBYsFX6
hdepr92IraDgu2O4R7g1O1SRZ/sJkfC1Jmw8+/5gSeEZnENGU8kaRr/Xs8mKL4vwzbfar6D+LBtu
vAZHcsW9scCXP1pm1qJ6rb9eWRdJrw2iA+vJ6tJ/ha5MclsILvg1ZQeKFyvenw32AuGHO3r0Cdpn
vch6LCdqsdTKGxPID2hcb3OPChoOVMnBrjLpkqoC/xquM43uUIVS4JiF2zrUWorUAr2LFiWVZE8W
Rf+n77pYaP0GfUKkbgTf2Po4HXQc7geSgHupRB5Xt7sAOR5z8n89Vl/UTgsF8xCgqq4B7LmzC+a/
ABIGtbSYRGj+No6BwZJXjIl/0us7Och9+zDyeL3o/1AKcyvi2O6LZyVp43zWDKZfE02e6+kKLKoy
8/19rynjPiJB0zHqUOXyCWZiTQSOxmbCIdwoljET7v0JglJYWUSsh9OLPNerva7PM6hZwrWhfy36
mS/Mnnyv1ENsz5XKiAsuzEsJaKIUPthLbSiSw7oRRYXkW2xJYPJ6moRAaWI2mYigc+wWyfUsfxCk
zfgjA/CMtJSqg7f+GPCmVJpDSAz7XuFp5JZ7R46POEDKFGBcWbVXhowfpcPoJJkvRrBKt63KHfvm
XGbZMJOnvb50FXc5FYmyYHly3PfMh8kwYddxnetB+PSo8ZCMX1bVqVDQkuwrad7SOx3snzBfmujy
QqsNkYog3XrglS6JcldKWh5s62aXIk4ecRguGl6gOV9q9TL0Y6WounurZ/RhrUGx5EOJypQFTdUZ
q9SdCLGx9yomSJlvCeAtjNsAtFo/OqjM/ZXzCP+hLpU+/J5Xp3Qa+cgL+pXNNHnJSlYJapRrcg9L
W9sxWTA3hywopPVszrWCVxFgqQlLcpRXDOM5XlAqO8S5b9m3mgzSu9IAb3GcqvPuFA4szrbBRFUO
guXhgDiyTp1Mn5ICQm3p/fiCK/8N+pl/9P9PF9GaChVvSL8xoXXlmRrSkBpuc/PkrQCHRt5BCJIZ
qXH5jYNvrqmiMUoPF4WSzvlw/pKu5qevSlWk1esAuW5EHQ7R7Fz+04WYKn0/xx8YODv0iN28ZjQJ
aNHdGZDT+uRdmYi+lO/q7CfhI+gJcjRt9FE38K7ZqntCbTt/4jei0vHts+1ugCW6O9I6qt1dU63U
Dtr888DCQvkqB0KE4Prcap0C0zSXxAeMOM0laitWW0igZ6OUpXMmjgZKR7lm73vQWrwOSx8LqAQk
QYx7F469b7ouWtOeRgUjIuSzBmGeE95t0Hp95H+R7ihjjD0e9dBCuLkpcc4/wnDePqkSU77DPG8a
TUAOWfzxo49VmLcbH4/GjOtxTpoUO0Xh0p/s9KVZU0xZdS5Jh+FbXbLuygEf4CSyhkW86Ydlngac
fjAuhm21q9Hk8e2KvpZ96hRhBjLVXwzy4tJ0ng0BXx7xhm1HDY24sRo9ZQwMSz74xqLZsmkTaZHK
HEoclgWV0N94fHSBwcyUI3ZLJExVE5bCUwn5KdmzWpFACkjtGAH4sZnll7bUboJ6OMvULA1CV77M
mAjjQ5RQ7g93eWpaKlpM2VZb5YtrajP4+Uq/Us8oC+jMcE4JumhmH18Du+V/MIbe8FTe2otLN1Ij
EAi0pNJATYEsZ4sXyOXPpSldopY5wwIOZSq2jm0u4JeqojZ66sAaeBo1LhgJUol5EhPMNO8mSkaT
2IPUb9zScqr2A6N2NU4bFvHnOGOl7+kS1+QufsaWKOe7M3kPV74LbYopH+gPiiRS6xbLE5oGMTpY
xbdsdQCQJ4+F8CSZchlMLJN6fwmSVri3JsiLsb/9Pp+D5UvvRB/MwtodYWkZim9+LIatRP8XUINx
XLcJFSVa2bXCB3q9AMur8YELqlC9zsau2qKMEDBtlQQHLSAOWHYaeBCNozQ93LV4KODVdnrCyQDZ
k4etuMwW8JJF1kir9Z3z9MfP+Wbqn6kZJfBzQPStZ0GtNk/Ws6xs9T1/cZoTXxJadQhCBufscxT/
JWVX76DhuLBc3e1Oz7D+VQixDwjRUVAC6xAcvuis9rO6tteJ5HliDjCLnZ8tm3lCKYolIwRwWf0W
n0JWm+BCCjreFoVdemyXlOgoL7KXcKBF6BwQYksAlAiFyEJyBUmh0SFxDxGY45gCHvaF3t8SrCwp
Yji6AfDhR68waQ7Dgs+q2FYTcp5Z+be8JGGjz1UfoEbhVgGcGJfRMxEEIZbr0OdU7leo2Eh5ZnQl
BNcw2piTjyIRphdu1UdxJoUoZrjLGJ1Y+K2ofKCMsboUGbrp8N4WcQwEAcgpxDUVMKMAQMlCUG2v
aZrTFw2Rd05118gFnaa9VaYf+HLknzDkn2cZRpacs4aQvrDcUhKkgUrhzAHCgvFMPYoZ3mDVhOxV
DCrrPIkNurb8Vt7m3nbLysWWI8LgM40JOwRGNlbBuVSJq29582jnQn0Y3KGn6jP7poEDUNaZ0Z8u
fWGMMBRCdFy0BDLU6cDuLeDouzywPcsK4TwGabCRY2eWaBnbo2468SfkJUCCFParQUP4rHfeDTP3
H5L2b/taxgZJyY9l3OCVk4NUtOxUOpAAU31Fw+Ygm46DhWwrAc1f6EcBrerLFjNPjjHNGiD3s5P3
dV/tzIF+MoBq1Alr+mu4rmg6VYp8SFnyWEXCsBv3d1BZ2jKZE3exMqCnhezS1TRZRFFO8pB57Uen
wDy9TBDIudu0BTf0shoCyjIFJ4uIxj0U2PqvlA3k7m8bVyFCp8bkJEs+5TVi9S62tunhdYyYBF3U
XyPnIYbfG9qCySgbLy9eZK+yYePBs+UyuoYCLZ2ckW8TDfl/BF2q81g33EfY08W427lH0CDVNOvB
V/Djpnn6nzCZJAJCA9vvYkl2/82oyJA0fPDnR/YKCobNa2TzY2u//mW8Xb/k9D+Ah4yzV20xil3v
dJYG+jNeuL951HUG4dWUyI4FaNRh3Vby6mTmCRLS+fgv2HaLUBDigeixbDKoQgq2b+L8/cfVJ66O
4ci8V8ZsLWsjM6LkOYTLP1aRjj6lYHhI8KxzaWVLcrd1K0tL/fd9vcRVBf9otSjUA5tqeP/x0RMF
RnVp5vt34V2gMhuqaoNGISHY8koHhpD+3H324OEKLMunSKJ3YsJQul0G3gY2jlzjpN5KhgTbDgmf
M85VwJjPY493kTtFLFKCVeXTMYQgAV6sIofDZ9r5uvfhh0CTdxFMcLokIOCaOrmeGF+XiUS2G2TK
myOedLIK1pftSPdQyQzBJU2zktDNHmwZG6YJmgeFOlYvlSdvHH/7Uzgmw0qYan+xlKoIbk7UwLMx
gHa3aPqYcK+7ITAmHyPVmkTzDLfKqD2eaW4cqQGM7FZriov/44shreffcS7eS4/o9zXu4y1HLbQq
/Wh0Zt5QYs2o+IFvWmsYB3hzHQn5z/3WqyH+dntvvNJAfIpA975zi3QSOuN6cFq9C7OcMN4H2u5i
Wb28Yn64EJqFtpQaRUXXo4JSwg4N4DVNN740YHqHCvlf7xoqV+EIq3QmF5VQKPo9rr4WWnkJ5Ges
jZUJ0alySbUnLyTR2IOWUO2JZJWae7dkJUUc0/3ad6CNquyl5kV9/Wqq9LwS8B7Ei3ZagaI3zoLh
gv1CqkfWBIOm8QSDSRyBgjAjjFD6tCn+pY872KFnjstOXQhqAneReD4vfLFXdIqJr856SXvhQ17K
LF0mLV4xY8xhkO6ZvrcYZ4quWxVaO/QC2LEiQFoP4a6mmHwYnY6bZu/X1A90EfYIc6+1p0l2Rij9
0ckv1bKXcZI5zW0rj8d9I0KbnL4NNZnOdve//crsXn49LEBji/kghKgwIC78OI7qJEIIlsbzmm2d
UVHqZ1D1DkOY8oJOK62LbPZgTSASiRvs75KdeZGIFvF8J7G3+oZejeMSVpdttkk5Kydumyky1PfL
3xwwbxb+fhEiW/qAiGJ4uVoYpVkcL4pRvva4CjB/rHw3bJjTJHZ0EFGf1xsRIFSIzXmiZumen+9m
XvZlJD/o9svzmRccUE2efT72c0xHQSYtIK3l9GKbnPgmwU7hh9Vwj1PIUXEnBaZj/5kDdnNOfEzZ
/0XuVSoHHOxJT1S8DZWJfyySmMC7+kaBbJg/5yFaASkvqBjdGH5VheVN1hZ67r2yHODq4cyqlClk
kNhpYsILMfaSq7dKHEuLC5Bqeo8wU7j1pJgkHI5o2M4u6qMnYvHpqy0fWkClPFmTcpwg5boNK5kN
0Y4Ebn9nJpCbGU44qk0DbpeNyvTtt/cHJUucAm1CP2OLI0CO9MSFTFw0mXFK5fTu8lFFyWY0fka0
M0d7aZioar6JhH67S5HUccGUm19Ns2RyMZhrBk24Z++oPztLPTdoHoYL1HCPSpj95Ng/RYnYvwDT
EBEm4gzoADGsINdsAVJEGVEP6r7akIa3X0uanSGDxKQezombIdk6QcDiYwgb+657AsEvy6pljR5d
PevVFOqpNEruj8fI/uV0eoFKrTFCH/Dz1yYHK0anQSZqChvHDn6omCfOGbyvOVyV0yo7LL4l0GCt
tUk/R4b+nzO47cT4Kop16f4RgoKr4GYTL3Bs3Y4Peyf0jS0kEEFNFA0sphWHey2UxoiNn3oUDaSi
o5nvco5/qcOikPs2ZBGG3MlWyrTLX8kBYr88QDiQQjxc+kUji749zGtC0BoZBJTwfzEsoDjKOaWM
I4M96r6wKm05hRDO4mClRc3vCyxdGn9GGoFjk0mrMyX/KiRoa9e3e+FqvTiX91kRFsXH3OzaPlO4
huEtM/Wdp5hNeYnvv5yrdz8b5ZGYEWsc/xZhDBF7+JKJORkT8EiUAb1L9Ylz3lu5N5I8FjBNcKFR
0dTb+Zh+0v/g+Jp3O7pYoa0n9q7JLZBbNSUzoS/RrP6SVtS9XV3cO17aa9WTRrwuwTvdCmFvgXIg
3sKemMqVJTf4OdBesPNj7kPPYLn8a0R/8fMVpeKIyVYbzNKasYKbs8idSvS2wEyksS/thNc5aPRE
4caeU/OFzLjvbB7mLQQHLya8rCpM8lZZ8XeSWCGbBlddk2TnfKm5oaUelhBvkNYLi6UDJyd3Xofu
YOjPaYxMTJDU9r1Riglt6T0VxlVOkGeWb2nz/z6KTpaiLgyCQ8lHkvREiMbxeHWGt1ZWYTg+7mDQ
TcvTiXXkM11/pmCqI0eKGrE/2+ke/cM/qbuNuMRHLr//ROlYu/z6ShFxqEU2Urmf0QVORDBHYIDH
Q98ItSAoc74/CuKvnJmA37ldoXCv7bB4N1WtTOjkGQIAkmOqz7h5J4FYwCTCaTMAAPWcONubPO23
NFkE6H8fQ5E2ZTRlHQtgEVREb7ShTZaOlHoU+rM5y/4eJgceBKV9DCQJvwNMVHs7i2U/C6Acd973
1Nb/EfP60TJ1mGQHY6OtsLat//YYnZ5PYJOfaeDC5aC2V26Vd2E2yvIZdiw7GEwKIpWiHMr9vd0C
56du+ZEXAKoRPbmXoqNK+ybuFg6AwJKVbieJq5e81FH7VeCfJT9MlgylNsctvRpVfb38VXbaXx9K
44/9mxNYL64wmUuxeXptg4tWWcXyZgMb/k8rVwpW0IZpg+VR9sLBBHUENqeVaOdldqNYISAIL6et
zqaM2PfiLCIy18HfEXCkW69+qdBWBeclpbkBouus1tkFJGOCEI9+klZgC30XNha1lP+IP+gJe1cD
oMRy4EBi2+8hYqv8gjbGEYXgqgYXLWweZipKb+xYo3ZgkvLJ2Kt9eUt6fUMN//ccr+pgNxEhb9Zi
tL60bfdZduFCBlnqjuVBhHYk4GtlC6WJpDX7T+/aLw4Xv2koqW84ES8Gux5Ig4u6W5eWvKCSxYqm
a+VTUSf0mz1RSMFX1hyD62+LYAno6Bc+vEKuayr6qLUn/YT+bFyX3F4ytM8wYx5kdOOM7m7z1tvT
w7ICZOnC+cbshl3tp6lpmz/akq5lskJH5tmaMEG+fLA8WKmDyeNYWGcLcsrpkaJC4cUyxksOMRyJ
/wzYQ/J0gHDFIlmjehqzTAWUbNPtidIlZMk26rMGDiJNqwoRsPL3CC6A3RklipnE8qz9EOaXGOQE
WT+biZz1GUla5CkJd0xh5CPbDEBRhSBNw92xNvXDXphRqr/AzZG2sAA39GoDd1DD2jQsDbMB0hiE
aI7zKAH4IRqtHMYKJYIhTik+pp+KDETIxNkpkBgKTTCA+MPX7SI3Ukj/+kK6NElY3+jWrN3iLgFX
SkLi1UCfP9vbTO+S5jvdg8gQVgglvK4ODaktvE2quWv6Oxi4gaJXQzasY7Xos16d1N3TWqSydxoB
QpsGdU3/TC83im5bmRPwmd0xFsUxKB1nnM/cC/TM15KTL09DNAY4xGqXBq8GASkiTDnIGlAVTfiw
+cOf/bpvLA9KetJ5f05sBeWlZncNooAm9Co9MCsdhFtK3poHd+CCz+DF5vd9RtiUgBtcWHAhR40H
37VqDd3qSXceu5v5NbjQNMBQ3Q0/txc1KYWV+I4U4OB3fGxPrTsZVSNjgPmmeiyNlSKwRs4oFckv
ZnUXosxBsQVjpGmyNPKYgIV7adD6O68D0L2CUwDspbctldVjgm5Vl5RKz6bj+9XFCURqqPEBfbzI
NyCIstSChP6BtHjLNg541Y1WAMg3SRWXbnN1isNJlrtKz08z//Wssav3/c1nZ9e9iy6JlC/+sX/1
4fyN2/NyZ2p85/BkjJMwuhRSPcwGhFU/sd5G7T/3VuslCsLzZyZNMr1knK1Z7UOfHoKMFHFrF2O2
GfafnUwio8u+KSJ4kpeNK0CfuWdFPP0QMThg5hAEAH2+W5sl72GyWD/xQIqWwPEAFF3Vg1AiQu/a
+zjeXR/5Q+lYgZxCo4BuOs7F83UMlmNsH6cy/OCxwSR66nfx3yZAD6aHqJnYp4JU3qQVr7Pg9R4u
dlU2/En/5WcIyhhMM4UOwCzmATLcGatYVo1VO2kkheSF4bbjzTKp+lRuCBOmHoyqk2mhkEv37YA/
v2MCcH80JeJm981zFeurpT7lkOlK//ZY+Ysu1koJG8Hg2ejhZk5dkTZwNUkWF8uAMJ6ZS48ZsBwm
xh0Ysia2TM9yCZjq8B+TpyqiU9vdOnm24GMqzP51etUcuPRC9NOpYoeTHTyFBJ7402KC0l4OM9SX
W9fC0NHY4nY8aSn4jrSy8MrPyAZh1lLrYRrjb6MtyrKPm8AQOtzODB6tfvgV+5wUKLa9rt1UMRrw
KX3Z6VZRvMl8FqBLDven9QgIUwjYAlXXKJvul4tNZTL9CeKB8Dfc+7ZXo1VQ+83s5pYxQfJe6fRF
wq7QNdPFtOaQwDxVINkx0/n3OHy9fLyXGntypa4xYvYe8Mc1Gu4W9HTNj/8dejxziTYsNJlWCvTu
7LKqALrIOOI0zHmAkWwjM1h8TRCnOOQwIKBkHJeNebfE5Em+oIHiwOipHq438TbQvf1iqiEn8bjz
35t+UOzoRD6vmo6qQQHnsnB4HzKmBeNI7J4/UXj+Q4UkR5c0Pv6lfGIqCpqIqNqr1E/Xqct2NWvG
K9mPAmIWWUlG7lh1BEYs/Z7RP0mFs2ZnyLRJ/bTFx9mMPf4KzP1S0yffhIJpolq3yik7BjJ5qxhO
Z+S7DU6MvUCnzpcktCmiZmpqQzBGXvMSiQws7wnlSRZRW8vHqlr4qgkJBMJ6j4jlseUQVbe0yJp6
gTC2WZqDz2Gm71YUjFmwWkB0ZY7VgCwlGt5Ls17R1xStnMdbd51jhGyFaRK2Motj8GuqKtziKD7F
O5w2lEpzJIF/h6iMq4C1HJlnwk9MWV0PJXYi8PiWqJW0FgNYYVKvjBSg8+BNSo7exh8coqyox4WN
i0G9OrTq64Y43tVJwdZYnho3mm9hEBIDQGObaa/9YUvl5p0xoJ9C2xZ7v5DSEZidpGrs7vzN+LYD
TVxJKREa/3x9uYnGZdLqe/qD83VCZNO6PKKr9l70xnHUoZj8AnslnmSDEUK5fYG8IxxZgwDL2p6J
sa72dIlwVWHep8npGoCYd466w2GiYPu9mKN4jqDNgNI0BQlf/loY64mA6WcFj36ixFZjAxtB/+Jz
3Wq0lLD0OxOohjVShuzLImPeIA2bbYSbZ5k5hnNzx11N6P2ZI9qvv6vTirISCDjBgfzzf2m5Bufr
VF/Dv50DrNeHwiodEXGQsesQJ9E009hGajT694wvpw2e4bPyTrcm80aW/5V/rdL2q5qh+7WPBiJ1
G9d4Hht8yWjT+X5c+RUsJon6zTDOebywhjcQEZJWZpVCktSCBIFtWLJj/RWqp2lvLr1z0G25hxm7
v0h5Loismdam2N0Hr8spNxIjqWk1nBWQvkz2UxhfeI+ItGYuuAr/idKWnVdW1gY6p5Gbr95+pWy+
FhiVc1LVrmHmizyq5kW4+55v+dHr+KI2S3m9+ohq4BsQUR/fsRu/bmzjdm6fFPGYQTRpPxpbWSZB
RN0d3GJ2PBdkl3hVfj/5f63V5Y+IFbgBnnw6Wl/1VyjDwuii5OpKKQX2mOcdJRha9QkXtLsO3AO6
teCx8LrH0eLIm2cCmj750rmkgwwCdZvPmq2Qbl9oXZ0KeJZwvHYa1KXYweJEO6yTpyv6i18+dwcV
NKzR2/Qu04OMGv6jdlSrcmCS5ny8wDTWupte8jsSUZ+o2Ia327PuKeo90k6MhU0Itv84fkB3guyq
Niehav17FB1IQJ3vB3L5ePl1N/QIdQw3hFuavM5RqmV2yYdu/OreKdu0wJflLDJUmpywKiB9nVGW
W5bll/ijPXLf9t2gCukLlxRkciTvEIN8zmphrIt1wTWMjCnkuaG88di+IU+O0dI59FODoyuR4DJf
+vK3uArUcP0oN38QTq94s7X2FW9r7smsGL22ISXQ+Dja/ViHE96wCyHpib+3hBd2t5JJixun5sl9
grvBrx38NlEZd91e/HqWixVgJ5Fxl/PnEjDTcSBEqTK9vvw5HavOecF+2KX5gDM1ZgKBq5IbM7MZ
B43Lp6Q7QKbOsX4ej42voaVxwiUdxwF4UuXVeT3lOtR5rmx+DdmVN087PYIH0zjfi+8xDESJQ4Si
N3g/Y1vPjtMKHWjCf5qzJVBbrMcNTirNlRUsXTicaqPZ/xeIMV/PuigPmYFYAFuFR/AJqBuN/xOo
99qnc0g6N5CVZLwQOomM6Kp13WQh2FAKv/CyiYgyj1a9yo3y26CAOLNbvAZcTRqOTzAUVrUwxCT5
18C89d3HXzHgdG1Xj5CN029PpfqRTSQvm1I+x6zCXddtPVf1vvR6Nag5MDEQ8Dtd+zuI+p5XsS0t
2vg/8ppLTNYWYiAhnGIsr0E+mIfaJwaKPpuvvlC0DRMw7heaeom9BBjh5O1CGBnyZ94lnvtyJTLk
YHDza0Cu1sEm26Q4altmo8gVqYo1JfYuYCk3k2Ts9N312iB/W2Y08XIKFqZ3KIAdZ/R9KI/O6BRs
7IyBaP4Sb//3XokC8B/VASjjvG5h5KwcIXUqK6L2Ix7wKP4oaQCsrUF5kPeOsY0z20/xk1nvApgt
AolwP2RwqlL0VNXF0A+4uOVveQqaoK3ODgzFlSz7nTKhafYJT3pt/y9n0AE+cItVt03BSreOOKdD
vJm0+YzUdyxAtKLsCtTaI5OXe0ZvUr8dIZGhaTudrjMka9kknLdKieKxV7e8vppxVaFNoQqWTFX5
hLqUcaf8iimVd+wMNleLcqii8Lo1QK/cn+AwJi/4tEkBuYoglmm1NanO/WAiyXHqD5VGue9zzb7P
bEH51jIZbAZXhY9n8SRn5ELhVNpwQm0RgYIVwK2rJ5x+ojws6obzxS89AjwJiPfJig4TtdNEooiw
dSiHXyZ3nqPM41my2U0nmMwXD5wAePuvmbRMpkQfQ/0anI95ApdlC+T6kp+JdkOJYvU8zjdtRxWl
9BHLuvoyTW+/WXW4g9TbizGeNe6/vSjH2yeGJWFQ2KRRKiUttr01h/IgMmrjspKeYAAItLupgsLL
+ewHILZtHyB1wLZCWhw+t+EuFgk2mpJUfao3B+RRWXJLSLPQhpzix4kSOSxiztBLKQYsJVTw88W6
0f1PSW/F3jA515qqfFVcc/GWOp3ahRvU9bmk6oPuGH4+tA8/34CJXXr4Vj6Gw5c18608M4lEsXWI
eJzR3H6OCyY5ZzRPQwIvrf3ZdhlisyaZVQT5dwXklVrQb7uFS7GKR6dIEyts29hfy2obAhikEoLP
MOn7aYAaUn2zvm2qLR8EaWpUuCp158yyPMVePRGhGZ2NqVAj3T/HrcMGA/vMiX+Xpjvre2KB8vYt
vPkZpwEBMxXzn9CuytYygfnq82QUbBmXSbSvOm4Yg3F+bGoBRdEEJarYWS+IlD3smmxOVdUZJ5cv
/mPRAsKRGSzu+XkrTEw12rkSR2vlBDqD67A6MNBc0+pzGmXYrFUUevmXIIOzQAZZpM8NsYcSdsY3
W8Q8P/g6FCoptq8yGm/9UdQiwlDSMNmGp03yyUzu8K1qpPJmmqGanhwqRMFX+cBTNE6Swe3vHG51
KBZwXM6Igupt2qUxPT6YY8kcr6K3rqYp0L1s6K9w7eTpm3iNcWw81nvjhw1cEJnSb9VsQRPRmycR
2fUOdcUR+T136t6HEt0gPxxG9oTY6XpUezMfNY6AJ4ZDijzHEHbAF0yGdF9aYh7TY0rTeXV4q4t2
NIzSOqTspKEcHS/GOIYqxjnY2TjagSr/rg42KBQcarMTatNAc2qgL3xIPZuwketDDGVWqO7PCEcO
uAGrrVKCZUxcqIPjauIkDZ1V+VUXMFjPIrp/RWMyCoESl03teZlvYfaU0z2IfyVaUx2HBQSnCf0I
tOqW5CXouExOI3zy992jUcPz++7jcrs2ujNHuj3F9z1/KqNRzi+hdW66dYvbCeSmCJTpiEiG2moO
TZ+7TFYAEYuFinvRmj7GbJ4ILCzI8lXB4wBuFQD+NzCp9/ulqyj2lRYh0VXCUuSXEggHZRkRCMFl
BFcHTnjgGaBHyDJvpQz6yPNaF3h69pHJkbuQUx/ATLBXWW7KJahjvmVHy8zpEfJ89tYpdwh2ptNC
+lTmwPc6MpyF18eO+oxmNeeO/Qyk1oxkAFbAryb0cyPL6U+JJEKvW1bUEuzXnCB6B6TiFOtLoC+K
gWxLygiS9wwYl1yGKmjZKJTZsN2xbZufmNk8uHdNdvfZg8kC6jqiBW/Fg34/J5zS93MkC93xon89
cXlUhbVhH7Q8VpEPDF2OmCv5DSKREtWriyADrWPxRJBdOu64KXUqr6xlGd/I6hTflymZPKcKsa0O
6h9c3FMWrJxW/zZZWpgQzhqz2CCVUmRIDk+Asdy5/owuYKQ+uPjt7mFdkl2JtIlvmRQ4uVOwn36X
GN1on0gcuvOHmBbgZZCmwj4u2aD1KCV/JXvmhevn+ATHUqT3D7QHqtAwTMu9TdvUYZ+I7BM2gh/U
BpS9fcG43P0f9CL9HXOjrjvjXAjYoT3r5dFuPIkf40nb/G1ddW4lf50fgTgutoHRbmbkysIOz82p
woSrV+H1UQ18nVc2ULoWoS5RaxI/Yd4UbGE55izqxbMa5C8K3aa7suTS3p+JrQ2tWM2EYBXLVro4
QC4E0y4IwBx6f5aQaRbUKeOX+bu9PVDF/83SEjEE1b4L4duWQywtLlx9gVg5PjPPRKaV3CYFsaJj
rLvJfDhG92vbiS6Ptm61yVpgwCIfYWVqNerGfDjGsanvMDmaIV/vktj9bwY0oxSSrPnxk9e8ybcl
gvJPIPLS22HK/HfYlWaKEcOntcqTzfnDeZ1o2AmTC+fLrNuNAaRmONFnzLEd052MOiL1ZD7awa2r
mbipT8mpU84WyRer6uK2QFdFlDHqrFcAOqhoiDYb543A9OYPEGH9XlrGVxlC6kueB7vLzSMfDvjV
3g6mFJSLDITwgNEyMKloS7HDUakVmamT6l7hhUBDiFQMQBQIQBGjVtdLs6BC+ayWZ6SMVp5lfYJT
VMZkR3YtYTBSGN7NqdQSp41FiAl92LXjAPWqBWsMQFSWFWe8Tvxw2BVc58TZqDdOwcFE1XeNzi6S
9PxQZF+pPU4pBhnyO/ofNr8sbb/5eov64y0PSMii1RjFz5NZaZGy1kFY7kk7+JVubpQdmCDQ30f6
lVUx+Xc5h2aovauWsJXH5A3uZFaBm+4HWzhxvQZmVOrRlqwIA0DhzNuCDgS1iiZiJBegLFDkDuQp
iE5MnXCr2GzvxzIGZGA9in3J9S9rbAhqGgt1/XGel4tzK03cMuYexdIL5BMrASXoL6NrLD9ThD77
kzHq2S7aNnSNulRzo1jOGET1q6zlitY7G1stDGC3njC2P13oId10sw2/o/Bl6cRLK1u7AuO6Eg0R
L4XmRKFdzplDsYZ8zLR/k5gtSOF2y9KYDGBocRFs9K9+M37NtLoUy3TrGq3IDNo8pPvSwf0BAzlq
xxvDZagDMJzncpnzMAk7mDVH0fbjZImpYFAlXVPBspf2xp/N9Ly4j3LYJesnkzsjcVhMaGaZUeJR
8QagBHbOwgFTW/EDYlqkqZdqoj19acdQzzIbFKKpTXMYS5WbS+qQSpRC+sb/CJ92PXqaxeM9bNGJ
aO2HNgDkNT4pJQ8IbAakLTyCWeF9BYeI9YaGM+ZyePHzlRn+hu+J/wXvrlfBO9cNEJU2q26+iuMd
jqYxUq3Xbxb6g/GETBlCIFpUBh9Y7Z6lvGxkw9syRX2XHYe/guwxsSoDdzgK2ddk+l7J51NvaS7L
uNFGCAYHxc9UMstUn7dKOi9AHnLjyQMl24zCkw/vleV+QX6T4dMPjT/BWY7hGe2cOhyuJJavNCYr
olow2bWdXiGgRtsY2EjLBGfEv2t3oSJOvjTbvU7Y90pkotqYYGbF9CIoSOnTJ5iAIHBUyw27dcCg
8JHhx7zcYwGzSaz5RC/wtZinfdQXHh7Mytj7K2VG6prmSgfJkCSNW0lu1K34GI8jBERuhjCKQvFt
DA+oTQuISUBVzlf8/a8GkMm264OTM7nF5/r58ar8h9qrE9fwqQOrgkFA4T3ZtIsJhfareWxl4a1z
1OkgmHFauEX9ZLkYpog16bU9HAKJP5thNnhzmqWqATeHO9CJJzTnXVfrHr9+oDppAPwID3vOLKuk
aN2ETrOhJg/vcz7cwRfRCAymvU197MVkalXIiOxJDgVh/MlziP9hH30YYl5Oqq8gxZLtK3V2qTCv
28AQHKWxV4vsy8sAvFu2y3rzPM/EesbFaK9ksI4Jpu/qyMaYf8saO7lvXOvV8O4B1AGNpqi0RsKC
L7MFzEXBF62EBa5/TGpaKSyJsFu3ry3Jf6f3WH0aOkzZrn8dqWql3sbfk5HTl/lz/hI50M0mdgfR
hTvyC6fJ4+pzwGiq1p79PHRTcy0JRotpVelqgzxJ/D5soG2nF8mk/dYvaA63fCzZmNUq0Tbj6OaB
h82Gn2r8EH6Mln3MnVy6cHyoktbJ1n0YLUh1zUVQemhaWaP5NVY3kmpZ29veFshdOBY/M5/03VS2
OuKbYudEORTK3gsHCBYazVvIeceD0K37r4YmDbmxQcEpq9ycvUap6uLQN25zE3T18TvbsEqO2tPZ
mUN+TngEbxmI9L266ZScBGUQZvIKnWvaV3ywfRLCQxnlZ5/CqFXDcK6Dz5lQl9NmDrZIsKpv4wht
a0FIO/aMl647sHEPdriDv5UN9Cbvo+ByJt1mc61FNlWDgv8HTd5BwE0JTlBcWCtNX0ZHQVVyQzIe
q11RWUzusnIeYT6Cw5v9IsV9w1PYHXZtgt0QjRn+lWRzpSewZUR2TX9SYaAJa7/PRBemCQ3F3JoF
THOwbt8tI08r1r45/dfG8mpVPx+8DmphE0S4aNr74EcjO1fytTbhL243tAT1P7giSQvabMJowy6m
kvXW6hQ8z7Xuyv0ex1U26K0lJtMLpGykFrnqIlosCJIbRIg5hN043XZjmWwd6Q2htG3keAMHpAp3
wXc5YhZHxcig+DtJyErVRl6gfIRk3aOViFottTKj+mF5qITD0rdEP2hzBuOqfWaGiUtwdtjL4BsN
VBUcxqFxyGyUToqsBIN+HmUYnIBJJb/ooNjnRYGnZmcbyoX86Bfgz/9z5DAq6bawiBqiEqi7ag3G
0Ab65XG2rgsjxBAzZSumJ2sKW3adnJB5QP1TgcmIZKLcZNIfOnZZ/xILCouVgw1HB0SwnnhTs0hT
ZsFCVwyD10Wgf9HfMZpaOm6Il4LTLROfnAvulOBKjSdig+7986nhYGS5JrfY3d5k8iJh/J3EzDVz
XX0xdRld9VxFXIu+RTueKKkP/XOwsQapHEqPhQjJS1bxicbkM9Xe0qioTJ5QZwzqdPBDrmC47Wyx
Exl3gayOew5KFEJsiHVdixgX7SsEqzkt+m1bNyxd7uST8Y9dd1j1vAtUSvqjLfrvRfOJHqz0rPBp
Vnefavt4n6SLdqWGil/g+2LWuPK3fwhu6R6CHfEye53Fdw0fMgr+Dh4o1I+V4HaYyDYlO7qu9DHl
YmN6gZQVYOCMmfVerOL6yX4kC5WKXt3gZJH79ro4xgyInPDKKAObz9YI7QosNrpwj0sbTCHpZAHI
I3VjHJgc1M84sNWFVQbnh43F6mpXbhv01crPA6Heq8SvNMyumCsgnRuncaSQM2BxpLcJgbm7/hxf
SqxNrvN3sD2uPwPi2Mh4O/4YFhB5x3bHRabHIEi1DVf57uKnDDfMMAVoCPG2l1smpV4re6DWGbmD
xi0mkadO2nRpXC2yf0qZZHdep1WMg5q7HW6VtCHikOYPyYYDJ0HhpRwEWVvVxs66rKzrAMIZUyf4
s3LfzCNW0aF27JsxagfFg/XS7x4ohE/gRizQ2loZhz7z78aGUVOWDd76Dboz12A/ShTO3+EgFyqW
PTir2B5yu7Cul++BxAfc915TlrSKAHQGBrY0oRA50yFjb4CF4YzUUhGWwP9+0X6Odt4CRGmYN+1w
ZW4hBMdv7N9Z9hCGFvGLuA64aIav7quwiCqaPumitrHMO6zHSQ9tuL/1jtZu82sAeRm5mwAg6My8
zPKxqFqDmLrCt+VlGAmoA/cscl3Oidw8gJJ/vdfiuEVc1Guc608XKvHS+2DwuV4rdQqkdMcmME7S
ecV7ThTBcEf9vjiOtcGhjVh2WVax1TDSAVqJgoXpnLYx8Qc5x3F3dCEA/uolI6rcDYniJtR99H5j
pVHWlnZnBISGK5f0dApeNu1xV2yVe9ZHE0MD7ZE+l27HdsQLfFT12XvOKvxtGX6DeD0jLDKOPROx
qz5pUgvY9CAnppngBpJVpPUkd7UiLG6bYDHiVkmhP+FfVsruUFpD3Con5YP2wgzNcoN24jGq51UZ
O/Ipt1CspsSc0aGr5X+iFLekB0RqU9scAgyxu4lJHTDE0JHyvyCWvD2cgw/viTwU9s7yuy0Mn4Nr
LxjA7aRiJpcuaDEj9Uq213BwgCG9ZzUSBsBfnxyviXnog9OOvLVNF9Jt37FEem+Htxt/Q7OGWJHz
gv5Pyu2y47T3dUihPDmbgqwP/PHs9FSteZI19LakADfAUJYT2o16MbFq8Z+4pAS20UBtbqm5t1KN
fx9i4g+ktt+AO6ReaXQl9Wx9C9DftnPjNSJudfJcvwQfX5R+jaseL7jh7yO/krW9rTSWYJCEHmJj
K1RkC/MwjBmaUx/JSZM1alXoCGP64eCblaq8n31s/hJwUnTs4VXsowwKGPvUuQ/dc9LgcdQZe4Y8
tDp3+jG+Eom7eal/8/W/b3VoQajC5g0tbQ0JY6znTMXS9EpJOKsQ0QmJ7yHRPiLPvTOXP9Pz8eR9
ToqI1owj6JfLFK6/OrgKF5bev1APmGxV1a6vHWt/E6HD+fr3qIWA3WwS1TGybaA26UDEfAGUxuss
We9XCFiJ9ArUqtCoKUgdWlRl59r26hWNpHto04wXlmrMsI24mBpRxIWoK5hDb0HrMXmKWY2Uzudd
nvHb8flPd2d6DtuLtvc2kBJWnXnlWvlBFt4GM0TKLqPBX/ZYpkv44LBgIstxw1YjWzfdTYq0NymV
2zfFUS7bN5cIAsYz9K96YbatgdppyvLjCBxVzjq++wvXbox0LmSJd2nY7pKcVBm1nH1l4uGiGG+F
Pvxyh/lru7Swku1yE00OyGe+2dcecxq3/QROLPJnv/JWiztsLAtef4kqAswmSMJXPgaO7drcm/0L
Dfb4nK7DrQJ5eHyDrX4cpvCyqb0dlGSzZHJwsQXRKU3CsOS/pd2Ti3N5RqugQfIEkoZRrKIrFTd5
EGUT9grQ9NzHT5WEoCCAN+UitrRIspUFX6CWzWVUwkO92ggTdJtfJkpOAvGnyT7HmRPV31zuyAfa
HVQ07LokPdOrKC2IdsJGoQzr5Gpo6jvhZy8xZnwnwchlfpki+c2D1pulNWQIbpr5M1FqxOcMU0ML
RWzN1d8VRkEzCUiN5Utz1qiNahWRbH28jE4BKwChOfcTewtHt8atEO+18s+bJ0l9v5qks77JJvi4
tUM1Tq1/cIU0Ob/joW+DMME6Rh2GNk40TnkALMBHt4z/0nkkpumwi2goG7xEGmLF2Qm35YVTwkRF
zUpBjIbPPp4cxME/5f83aF6igOTrZU4D9bXSq9Kd5yEyMbsAzv6zf6I9rk2+9cYM7aX80lnaH60E
ApknSjF07wjjO3LzkgrMVZYy/VriojLDAYPjCfBbbMMzXMxnqvou81KKGMk+/xATM+AUizeK3ztS
6huEoa8ouPsyO9GHbu+Lj/zQ04YIApmqF0K5EopVXrvu3I/jmMuFOmixJfFMZefM9J72NO9azxhe
J8ZVbcyzAy8vEUk8hKA31qbcB3Ql5DgQFAF9ib0xRH7pEecSxfU5aMulufeWknNXNXGZg5Pn4Ms3
j/fYpRQNXhsx+bXUOB4Zgj4xVEQPMwyjGBEDJRpIt2wY36BSzZCW60t+B6C3tOcBdjPlqyikLHsA
HLqKh4XDqtEgWM2s5jy51R2+mXL0mbO6mi3FAlSLyt3JKBs2CA9wu4J3tFe15BpVcdeVpGb54wvP
nW8YQmfIbVR8ps5kmfHlFpLBmAa0CoY+g5R9tImzNDJ7uKjgwXOKbQ5Nn8Q8xaLayd58L4KKt0aR
17c9M0aYZ5LTpILgy1w2VL+0S0+eNtOk81T2CQ3jsJqa4RliI4Ft5RPe+BWVkNBWEHKDV6WevmQP
OrmQGZ7MUobuPBcm0YsYK6a7cRwpFhZx/myG1tFV5Fu32G07dWpgGIFfvBXaY1Pk0h6sQuFlSuPk
2Klh37NbS76aG72DKsm3iAUKciP6p3ffFPNOrCnX/1OrCGfvVkgmFwvb3IUzHK3mYe9hfEza2UJd
RBVt+3XZY9iavKICzDEukrOGQn5BezpYhOdli8Of6CDUOafKvQgSWNSPXQFZ4qS2Jxa/DHLE6aMX
BP3E0AhPPN1WgqJlLaaxxTns9vN/MHU8bGicj/2og46EZkhqixlwgmyEEYC99Q8nlN/DKpp262Y/
ee50jDTN7XmbtpbDm9TYbaqDEU1BvjOoDbfiH1a+/XhHVdQF7Zatu/SMstpwatokBGTyXqkiT6tH
Ufo5YjqUdF/K1SMRiLWYeFtpYYWveOlyjvryxcPlgSZ1w0/ak5fsd23fsX+CC1IHMjfuYeIbGkP3
Y3NRxsYZsO7a6bUtAwc9MwSn9OSqB+4vXawbI1ITer50E43hFKOKHMlh77lRfhIWB0fNDpaygYr2
rCDK62qrITe18lBor7g6XmNbdtoQ9B8BW/FKdawMkXDsahF22s4tRTHj/OYKpNbDS1HeK2xd0cUH
566rO87g1g6NJce84Eydf9Bqtp3WXAb76w8UgK4RLeL25AaGxdsRQJcjgjEnJbavWkBopRwlov5E
gN99zkgHSc0n5BsDWxvvQo5RDkx0Ra5pA9ZI7iSPIcmbWBJG40KJ8jsOPo7gaEs0o7+ZEXVbosGv
zHp4xYwzWV/gR743npLkmgmSpJO7tXtYiNPA+F3/fJyzfIQ406EteO6wlT07FTbWG0+5sf4uBwC9
zrD5ZN9FDD3rWLLE5bDaZq85YhchKVJZzDyZpfwi3isnisndOq8jHp6a8xgb8JPBup5EvEJTyFDc
2Me2qXHgKK3w510MRt8jbm1H2efHjBWWtkWNsLKJ94QYN9mqlDeuA7aj1fOXA644OBWfyX589D9j
1KbRuNuM7hnKGPpNUcQ1Xjzpf6s4PikSR8nypuLp8H88hY+tDqpca7rUsXQav5KT8nU4ibTUQqIc
QB3dU4+9kPJv3syklTCEi1HMOHoZB7ZH+9khs1Xj60b+MSBbALplc/z+0U9tIIUplIdIvV4Bp6Wj
EVeQA13E+aMJclPNvVHl8+sUth914fAWGLkB3xGElvv5X9Ggr81Uj4+Uof+Ik1j1/l51jLYTSwyc
mX02F1e630qHpvYTjlc/CTRC+pT0fylmtQzK3NP7JnRveniAySOwx5JMnaC3uBsxXC392XvYI081
A7en4Hyqnd60fdCZpNb1nhDC9sopJh3c0OeSCikFRtYcJsSmCmnIMwmkt7XJJUX++kO4nuRNIyVP
bPhLi4OvweyxLb9d6r3K8n5TBkH0TVysdpsFFsE3FdrlL/CM2wS9U41FJHVqSbep5AFyIZz2XTIP
pk9CSvSQC/AtO2wK3OJMCuHRksQQ4F6OZzGuTk1pdsoydAJD5NZWMiiS36ydSh6yEPmfw27I8IuG
KVNbM5UewEvZO4Smlffi1G+2ggojttdftAM0MWJoQ0ijjI4A2CEDU60tJ81cy/N800BRj/oyszoh
Vchnwqv8RQGh+F2aithk80ce0kvj4q31RbQjrGGbu5qPH6rFHHuHnKUPxFT/eqKDSwEdDCPz8V43
jn39+vu1IA/JvHj1cQM+i4mzy4SU2tuM2Sk+wpKCE/ah/d3tWp9L+4nVU0858JR/zmZ6O3+9UOzl
KZSaIw1Uj0s27K5qRM1RNgGGyoepITsGlEcTzElaGUSDiBLQiWahnDuM8F1/P0C3sM3pHF8a+gBJ
dKy14qlvSiwZAq3/gb7AtmOi50oX63LzN0hPgqH36Rep5PY1yD2lluXtar4UvQH4AVs02zxs31Db
aXfx1p/t0C5ZewaZwyJLlu1MNNGZYFeHHDcGFBhz+Kb1jptUig4dE8eVoVy62Qm2o/w7vlnx/fm5
i+uSyF7qFGQiuL8gQ/+QbSddD0A72cX2ExX5AZrGOOyO5d+EmpgnKbfJ6DnZTIgLlQY9STarvuxz
W5KLupzVUK4Jyn3TYJ9eYwzdxkunV3z6NqmNes0Y4Xs+zeN+jmW71dkPIMlgl0CszOb15Bp71ZMO
WJn0rE6lbhGUhRzx/fVX5FZ9+vfiYyDTYx1inPvb1M76UNx2Thc0/VeVuwJwQ3HZDrgR+npd5dqa
lAzAORWODkYorEtSrECD4wVvfzmfKMR0aDEWeTaRfJIt4XyTJWIUzqM+Ioxd3tS2Zc/2tAq2LhpW
dbl03SQ7uWvLGBwTMvmcYiEAikuEKrH5AbuvoJUH7GzrduaLMeL2/g464h/AM3clDBWS3qfCqwzj
759pb3Kx7jUTNB0qQznWcNfVfhANVsVDNLdYRrTZALMEmTYVmQSWPj3UD1NnwgXabS7PjwxMRdhp
OSl0Fe1Ztk1JGEt6CwbCGGiVS63+TYq1L074vWjlepXgHpmgvoVtIxFKhgrcSi6yeRHRa/kH1CQm
tFeZYM/yvc3ha+U1fhLCVI45gtoida9RwRLyjVou6gumoqz8algP9xoFwQ3gzg35dhbyprE0hpoi
6Tv+AMD/eqKaCbXKb3JXdHQ2wuRnbndSSDxLyC2RQxj6gHwTbwvFiY+L2tc/UvxJJz62Bs6QonMC
x6xwG77c7ueRHV77i569+ffnn5Rk3R6jUdGsNX8A97bXn7c/rFl1luqyvufhpoHkSxu7K5odTC0h
2x8IL5ehTRHqtEfbd9saf16Rwk6PA8aBGrz26wMMa4D1iHKPH83Yy9jViCo9EJf1aLVrAEb+u6lU
2RN02SEm9IS1wEPJLWT4jAqxTLHMM0iMUK7NNQdLTRf1OVkxfJL2LKiD7lvH4mwJ081kMRVoKVTf
Em1WboIpWm/R8MFjnqXnVh8Mi9iUop6z3gt7xZt1dR4ACDPxEVgW04EukSV7HDPLy4d3m2QfaKkN
MFW2PWonssYGVw4dyINlUBCsj3J2QZNqi0TOZnhFf8i3Fe9/OW/TwedbyRQ6UV17smw2N6XGND5R
ucETr28l5bsAuU0wDHAkViROUVmxEwA4/rDHp/tcFOV1cuuq9EuRZX2CGHFqoHO8Owb4g3OVCyDV
QGmLG5c39/7SFuaX6p/CPZlbjt1ioFDEll08XY0lQ3ZvT9dz1ZL2wEfXjCBdDLd0OwzAR67bEcG2
jpc9JYiYEuTtCnu1e51anKxbE7B8Um6iZ7raknGmbnvhmgchkOFCs/J+MG6RUu89YyDgpmLnFcSP
9g6w4t9xr0T5h43wKEGtWh0XvbtncgvfzHINSEQHDPpRmI2WW32qX2i+iDPgq1HD2iav6XOhtbWw
gDYhUhgUIynxtnP8c5MLck7jlVD6bQnsYIRM2XnuZsTzvh0cFjgT9yD5N/PSZ9an3bSmbKSxG7xO
SzPhTRYnRrbQ992mOHzBYEuNgZ0WJ/KluyqzUTfFK38nDTnR9eGh6pB4PRX8bKHXm+0a5mJdccw5
V161maZHZNwlBQfeuPs1SXyA3vkF1tbVPVAKv58cEUSfkLT8cK66oX40rYnaj+w96N+lCPFroPTj
eJ1/tjq7pmGUcbupIu1qVCgkWwk7Bbg2m0roEOet8EhQFoawq4FczcWr8cZRWEZcQxDnkbwu2uCB
AP4RctVqEfeByRo2VBQS5RlOrYooBZu+TMmi7RytZ4HSet2gHanmAabUkYCmnQdVNJppRoeC5fe6
cw80XJtXrEee1MXjW7+f+0H7028GU/im8Mud7/8+xfL6xVYibsv/3ItsUtkzj6KVJbHO16fd3shi
TlnnW9eW+NciGMBvAcEj/c64L4RiD8SjQHFAHnqzCw7rXto1gIBpddh6zxxOoljlalcz7J8RART2
vlJo7S3lkvCiBaSMVJIMNrpoFm4c5DXlS8ziFzl5uEcAlted9UzDwKgCb6y8uelEUUW9I5bigo6D
fx/7b+pOjiIurCG+/ouuKwWKx3Gp9+iyCH0vxFp9BTTsrJBUfpsGd7u7l7zk22vmKlapVOhzCzzQ
jq8/XsUXMGx8+K7Tg6SLG82G/LytgsxIuhYODTwUh8gE7oOhENWQzmGLDVpEVnwAyvYEl7hxRC6b
Q3v4DG9OmeASsbat/toyeMAeB3RoSfj8DH9ZfySmeno9wY8l3FVKv7DZisofhSVkOAuPMfgB04Y/
abqfLeADC6LYCSPnAIRKKgr5yhjau0Y13fP3pQHmAwmdC2jeZPd498KVVkpRD5cWcy4mqBs2KgCa
H2XDMJi3BLCwSmd9YOoRrh+xL3osgAHc+oruWJO7rAn44UVopaJslNV5Cy0ZrUXEx5dek9qUXdK8
b5xBXYLu7g+TWqNg5CtITQpL3vwx0FgwMD9hr9mdpx28t7qVibpIr8ItIbf3bUgAP9AzO/umOCTX
UbEFbehSsT4OwwFgZ3KtQD27tcSgqM1kLYlYuu5x0R4re8W1qGBuvD8qzaNpOVUFk6qFhP1loM8E
ZsPzIDpfUkXHx4tHFMCW6uQlGgmVavypB4UEQ+R5lOBazFlMUcYrJLzraa9Z8S83j6M2lcQ90sKB
TtXm98dc5vdPiAlprTq/itSjoEE8RsfidPoU/1rksC82wfYA3WXc9zikoX0ZX8oGbcr4fFaBOTm6
7zZXKDM6rfeCy0b2T01hPLaYDK9QPG0pjqg8KzWxwKZPPzfHaClGxwDfTmti1rXY2/3dEVGOvA2S
mOHfZpyleSonu6KDIQ9VmenhLipBBM/LmCGPGBL3fzSavYQ+rd9UL5VB71kC8x9a7jAZvPeIWlJU
IH1XiP/CKruwJ8jB1euQx5cWhoDOc8cRUdkMOYSWW3fAEKXLNLx6lHJTxOvWzC15UwS/Q0D4I10H
ijqmNQCHexXb34R5CTkkrcVJ4ijOmd7klkrsVh1GE5h/Mm5Qqb8tlREZuoW2Xg3OOcUZCVQsbmnZ
w7Ch5PAchhhAckFuwQOO0zEZ9PkfxvV+D8h+VDNetQp/yD5C4OK6j54S1UZnnqZyk/rTvNSXn/JI
/TfRTlDWsdVnTUkkiuyQrmnBIOqviJcEpuowUAJCysnM4eyZhroZCNo/or4AahZ6ztjJ3770wHqh
4m04kuKlBSWUICLV4tVBVqD2pUZUcQJA0gdsvz8lpnRXJXamvy98N10H4n2RFdrReh1pANEiVnNV
aTlcZOLphBnO233NwL+eTKZMrE07VYL1MaCY26ZsfhAAm7w9glDTY0lu1ZPS2TPsoubIMWpx6OxK
AU/BPloejGUzSrp9Wv3Xo1m3qqqnP46wdaQaL8mZBx9xePt2+3yBeMapuNI2lFde9N2R7c64K5nz
2bNHZEabqRAEtLhIDaJpSgsDKOTc7tNzis5HFe6g/aiIsW8MO0d2beZD6mCVsOYwEqaNwvEYosHX
uqr/33AcK27b5HH9WI4HtNy9hZHIgekCGxY/15t6JVztpxQejh9u5a1zV8XIBF9kIo9ZLh/s/6/e
NPoMks3bNPr5KZOhrGxyOtKSkLFT/784vvLHD4rLPIIH8Hn+wIouDvshHlO3ruc5LwG/QQLP0gdH
q6M//MzTMbQgfVvnuqqjC92duOxNikJdvGV7+deTrQhrXOQ5wqUShWyh7k4UC8YmV0Tu46iP+nkQ
gIYuHW/QEQnIev/ZLUPeuAGCUnTLXtaeUsSLy7DxnZ7JAvBWtE/UvsTqOWnR4bjLqRxFVT+BZ4Rs
GNJf5Al1foOk8fhUkGEuntJQ/kvuIq26KckS9MPaaMr++tMpDlVmV4WaLwVQ6qtMLblQ21jh3DZg
xbuc3ZfV36Uzv4pLnvmkCqNO5OXnp8dQr319L0K3HuvfJrFI9h8DLEK6OTFqXLY5RQTNvTTBdhGH
TklWLS+LBXfg3o/nSeBH1B+VY8t+o6L8XXHv+xFI7dJ7fsi9HFiAeQQ3wDrYq/P+0uiZgWK9gHdW
tyfA21YgfH+uShU/eWsVth9xylyaaucXZE01OIz9babixoM84fuPeDU3cxZYXcW92fQoChCaJ01x
NoxSD+aLpiSWgvvoQXfrgrHam8UZVyetRvbfp3h5ENmOiGF0j5wj6pSVlZyxOZdTGwcVdBGdaE/8
w2HhbNlWDDtIgotJJfUdphqPIISblPoAahuZPXyr8C75Jed0O0++klctF7ROZLsv7es+owbLdxWA
NVCG3k8HZN/HKtB/sgN5j+VbAsuRSsc2QRryoWoJ1LNKJd+ebof4R9J6PQlhqHQPpDevvRrkD31t
dUvyAx7okEyB1smWRFQY55NS7bcG3/FJ8yEsWtwPxyVVA02T51OMC/7ltAjz5K+SlCinuZbZkkXI
kiV/PXiVb57adfanC/BboxtzA9UumLxwIi7Iq8UogFqK07j0xGiwZqX5pE7iRafK6zFLAtwcRcoS
YLeJ5Cnmq8VaLf9+5c+xI9ujGAFONtA06q8KSdL7Mvami4ficj1035S0OX7Wclk9hlyIrVk0oSWX
wMeWlWRxBZWymaiUSDWTWfI+u+gOPyQKW5lGKdIAruqMlVELsx2RSJ90Pj+mKxN7NY36nm7WgvOx
ahUQTsG6y8Gl0OFJYf4yO73rryJ9kRcBIq8qpMd2SVniX7l0/9warXyi0qEaF1VQBCXZFfj+02pB
FVE0xfRnyOjElMNKeiJ4f2TWAx4pbI++muetHfRBFKFNMf4kzkI1VigWBsBMTNlsVMDqkJ8D2d9n
yQCMZ1BezaRuHmyYlp/awzfKnzldgf5xy5XowHZwyZEhS6/3wxLMN/z0zgCfuWIQXP7PrVZ6aDcG
9mNPk6TClbFoF2wGFwcxkwZdXV5mU13VSvadzj2sLpdnbg6jFUreViojuz02olgDmeE568Gr0sR7
RodiOiU3z2faErSQJke2eJsm2GE+8ZuicTwRkYszcKgRAnrezJb+vDWf7rDy716tkzbtUffRgWC9
DGIr/kMaKBw00CBVjmaUT4EP1ur0OSNQT98TMNNYeHCK5mnZ6aCLvHs1X7ToboQlQbuM3GE73aAZ
IXsFnGPZJM1jmVA/aii+23NxTaq4pXTBg4K8b/Jh1bYPWgMzEAH3gLVmBjITUieYmn3nD+ZMrkvY
wx8Fj1dPY+JapNoz0OmNeIUaAj4EtGIC3GSx9qy4ldkwm+4UipIP589EDu/sjVNo6om0a1UwewO4
bwHKGP14GQue52eVD8J8bo8DRp51vWBt3QnDcTXMwPIc4TfRDdyjs5IeD+sQbgw7cP4fJhhwmwQe
231tjpRb5hX9XAsYphb00T8FwrShUOSGJtdzpdaFNRrJhG3nfVZTD76rFprxeQEtjFje1H371zei
4828ziPtOT0wVsjnX0hXblSgdgXTR761gCU2lRmoUJktk32Y8QsaVAOWGoxtTl2R7HDemChEj3O1
remebgQ0sGU+FyPJ4JOJUcsLPMiy2qBGRu2meFfjLymOyLuLvBrIIn+vj4cCvhwsjMdsbg7TS60a
MPA1Y+q/iarSzcqietJAKH/TWlLWAiyZn3vUfpnpK8/eRcm26Th14aTha6ZoaNhlueo/RuMu74rf
D7wek+ZVS27ErzfG3fEc3uum+dbbM1FN0s2quoMDaCgJ7eoi+gaE27+qwUgCfYAhY3dhxQFQXnfT
Lln2fKjlfZtm58vBJWbts+DMtx3dKF3UR0wxlhQTRfF3IpacTQeFizaQpK9XOD05Gg5U8bR7C2zy
/K+MSYySMvrhQLDeNcvnMHzxwzH8GTnggDI1ZiLBiJH6dWvNnKgLSxMrwbCRPJ+aYVc9sS+Aazw0
0CBMqsVkWM0OzV2N5hb79i9OpF26ij7eY5XbEUg/qtD5riCajpWq6+ZdgZSv7RbJDFYSbO73cU7m
uEszM13BZHsjBH9v3QDW9KPmWZnkaVrv1oXg2QDD6Bfmok8VZqz3HNPuEy+2ytMasPEBdepkXMhQ
wt531jN6GBbIouS6GuQN36ll88tahXYf+SFL+WMVKfZSAiObJxRKvbfGrbf63vIPM/hbnwxZ4nLL
OpLpcvw7/cjxcMnOMVcdV6msihoWKB8zsIaEC8xrqnaXDJDyN6kNYKmAq8hJabgeMMM5qtngvykC
56pSlyxhTb9TgUZ6JAuYje/8r0ikO8OqabDMWZpWzw28oY6jBZsdydVtaWkUtNxnmR51wLSvmMXA
MVjJpyTdxzzDIDoH9CPagcoouSjHx0Zrw9w52ALafIGQrsTHSSWa9wnjrRY2tZQo8QChOwZykgzV
/z5UVaSq2vnDKB6SFlT9d2GrBGPuZvGdqqq9FNTsJB/JvUnAaRHMsL1Ry54l6txO6ins1gQLFcNe
ZTU/wNLWl/VAL8vSexVwC+Ze73qGaVrriAEupmanVaxJ45g8hMwo0LzFL84umH4P7jN9idbshzDh
fxbnrGXJAouePaGygZOTCTkgHgDe40+k1CXO1Hwcr/Z3dX6AsG+2zcAY9iOr9XQf16BaHuNYOMBh
N37j2NKTqD54r7K94E+eeeXQm7Up3DnLF43gHqHvXhC4a86DtxhEc35ArG/OxFFeRkdakIPb4HUP
DW9sipeYc2vrr2XClmwBRxAttKsc56YmOUgvgVXfqOkrd59RB7O3Mj6MjRKxeOkMzvKB0au6WsTQ
y3bTvu5OPWfTQZU1JTwXpyiTF6Ejt0yyU+DqG3QHrbGfuBeSvR2U2z5z0a9YfQJbSGCLvdtoqOAg
5Wf2YDtybjgV5arPsAI7iNtfwvmVZLeXmBLA3mc8EFvcixSAkwj2W8B8Za1MW5H8K+BkUqPCT+wm
x81qBOvMpMnSvpGLzH3+9pfN0NLgbDe8ixUMFk9e833n15Mv7KnpUtuGeYRrOpKkbkHGTjTMsp3J
oRNJzkiIZsl0LdNfmKCwEi9NzIyMMgb9b0/0iqJXG19m1ELtWL8FdF2UFCDzvLNxEKWo07MIh4V7
82f/fmUZoUdHSH98N4FZNfI8WrUlM6vGWHDsMjEOpZhtaqMR2cfBThBwo22vRKTjH31X5tIN/WcH
r3ub12kUpqySRZ07Kal/MjtBZOEcjN5WP7qBLiV1qKnbYd/S+edPU++cMB0paGpICG+ZCHDeAIp8
2mRjEJ3nyIDx7WIZbToX8XPUFQFj5F2Tyql3l/Kt4kcDwPk0TJDQxTGcTLAGQ2/d6GCWU60tRp5l
88WLuiyVzATc3HDgm7vB/XK0sq5d6MBnEN39rDXOx7H8qJQI3lYIf0h8YB+htOFjwAdJ5HHR4Q7j
DSeeA4aHm6fNZW7Rd1EHklGot+1kuYHebpNH5rtHyxPEavxoSXDU2YEBhCjdVn3boi2JgjImaKu1
AtbWsSXvMcZqOmRvifuCIDaqcBcmDVXghxejnX/Nb4a2lcclN9Cz1OmqiQDw3Pp3PMpN9lYaThGs
ypkhpSW79264Zp2TOdh7SdE2KTIzMsB99Tyaywuc+kGzhfokrIwoicU0NyWVt6DeHrIVIsYSW2Ec
URO9c8N1bzMVQuDx56WW4DrzKKQeIovBuLetrVpmfYauq2czi4rkm1/VXMzkI5DrBfi9kYMzZ8Mp
gZG4o6TS5QjBuOM/zqxF9obe9xsOadbrEVWSAVxq3zpxgccN+iqIeI2PVVlJlUC6lanWyiHhcxEI
BnReTirSIJmIbzjlyMYIXNBwVVJ1Ey8+0LyzJmyLvwQYorz3jqf1AZSUmJn31FtET4GtblmQWCCh
wg0RJqX8H5w0H1S0IQKnYzzsvYKCltf8P14AFXCGWie27Wfct4tM8FP3+rqjoPaAhuBK1ucv9FS+
82zaebqDhZDh+tW1pX/LMVF5R8FI8LdB3V7rq9P4MLGJsk/D7UP6gGRKvuwcrpKrXODgVN7fL5Ru
fVVXRn/g/xMPlwETQY9u1m4yha8Or47Ko85j6pXavMweWhRHsEVrg5lYPYQN8/76gXI1tmj0NCcx
KvcW6XrHhjVczCiBA6PFsVGXKiMBlN4ZEdrWW/DYl1WrPUCaIKjbmiCIkI4c3QBdViIx+plYcyJv
DwYhlmh0xdFQJZQeqNARluD7+vNFS9eyVOGEHfexddxmjM69Cm13WXWtc9GhAxl5VqaClG8dxKhA
v87vUs8j1XmKN0n6dBqvI1yzEsb4DkK9viM3LOv3a+IWyGQNtjyKs6e4YdzNKiRjaaexfizW41HC
JUURnetlA2rhelIf62/OuTgvj90CdOX9VFrnYOvFks8j9xEcK5WG2SaMhpnk5EZyddBAbbrxqB5o
ZRQw4wR9GQRyLVcGdBNHuKtO4MV1BIhq8xUVOb7uL/U1qtX7NZZsdxN6NzDATkQxmFg1ViJiyiKB
kQMIHqWIDWZGPubttsH4qV9N2BkMqCvs3OHbvkl7ZZB4EBKyB0qVPGibyE52a6FT9vpz2wtqNjbY
CIoMegD2vdNHTyxtCs/1TQa3RBFrwKgPomlG5T0Hazkb7trypEOXdVIQY6/rddZJoTUoVCsixYoD
gFQHerX5D6hSvmqwf9364Or1eZpBcuJEuB1e3ZLPdWbHKrwLNcZ2mQoq8hKpbJhY0kzYOLMymjO1
WJUQHTnDx0CmG5Jqo/H1It4GpOdNioON8RxZaCLGQxHfaXPCURjhVD2In3ObL/IsVA0wOAD3pjyS
MGEWTsz9S8N3k32GinFY54DRoZFrdtneOPiuFz4ytS6cz56hWC1p2npfyPN/jnGpA2wsLeWYP0Mp
5b7o9rReJgOQ8/bCDucqaRw0Darkw2k7bG1b+Gg+ePgzxkmWiEKkL/aM1WbA3FurIyLNdLfhQ+CM
1cDq+SmzbTca0h6d0ycCpFxaqueF3JJEs5mSCBmjgqJB6XGXtFKnsJ24WWxrPXEh428SX5iPoK3F
dQxVLGTGLg2tyLP1kuVzKP3McxA8LC+Wq0mQrQoMdvZslq13MXxTAKUTsukii8TyUcPQxx1c2oEV
oRLS6AUGHO7ZSnT8y1Wu06FQ/LMRch5M6cix4cux55lcke2Tubg5muBXD4j21oUdDVL58E7z0fke
zKlAqQ5U2K3Oxx1l9aIgFw9RYg4c4CKrSZLd6IolKtoViTkPPhJsydzcnFSoI1LQAm3Gfxl1SoTC
iw3XWjmlTCTwiKoGGSAhkiwrvA3lyzB1FdtJjBmL3oSt5gp9SVpbvHvmiowhAMnLCmDIcJpCFn+u
YGNqWQdCQ8kmTycPxqSlaZJMxqbADba+lHQZ6BdCkgI2NRV2verZLGQ2JqQv5UJudfbXZLiF1Pe/
ls5RVA/g9GjACl+Ibq+YYTMnhb2PbUzwKkwoT9NFUI980nGhnNBIMAB5DRhALv6AEj6qqg8v8BrF
MAhaxl1COgmywJpkVDplVJf49kWzqFiSTRy9eFbHAqD5FcRHslAdk0XI/tS9Fb8BzgIlpLyOd2JF
RcP6RgrQQl6UqseoC+tev2Be7A/X8u31KRC2n6bOJfk6l9e/HkwizWUv/R7Uvu4hBxfzVw8cQd5t
r9hyBVOIKUGg6Da/fAFjfcjC0WUm2Jnry/ZFTtgVXOhuC1GhJPw1rcyfMQmQFUHl+jWycfa5/Jmf
CWt22WWtFG3bXJ1QyfMi0XeouQV/jxwI8w3JwqauIjypUhiSUGeK4SzpjjKi2C8h5r0bJl4otRYn
6+XllEpqGSR/ljis07/o+Ph83t+6S3j226Jjr3KLoV8RIrwEWsA8Y4S5j47DB/n166GbH1qmM+uJ
thy4TWCQcN9Dd0SmXgU2nf4lFN+wbNg+W7oryzAgTYwNMYGsq0w2P8oKONE+Jhs6qttxFoJod6AS
r5rX09PipItcC6V2kQL2gEnXPVlbdb0e6ZZd4+wKGLbTG5y3SxB+5tp9JUld9RXEmzrDyiItV8Fg
WmBBs/rlyEQKPEkagPitnfEQSzk4gTVmUkMuhbpD7l3CgcqxJos0P5LuEaglucsH17NuNi2Aaal2
cn36P8lTLYYON445hT5U6pPWohc7vfbVwlRe1/bKoAfj7ZRST34UOtycfFylzPCAaOEnzquql77C
MXa2gHWdvj4xwpbZiworuiHpnnzkGMpemWghYO2AK29Iqs5z5fvm8LxKKJIbQFkYiHDBiBGnh6hz
/ivm9DiX4nnRQdgq6Ix9h8TPtAf+TKX9q4y56xIe2wT8yrB4wJy9k9g/RACLpRLvGydkdwhPsCvy
i1+SBIENykpkAERTu2hkZaXsT6j1Y3Ij/AqkSaOwuq25Je/iC+C6VdhtHLgJuU+NZpAdzFs7qVZS
AvC6ba49m7uY6XC6VP4887LLSR1pTeomr39U8qd4NQ3AueBg4//YgGAUKT31ljKFaJIhU/K4mQFY
tuIXcaPm+ew4Twby4D4pio6YNRWwPEKUb8ouL+o+eO31Rvawfev94VoDi3s6CKAkC1RpUWjPAHpV
cZXNXV71sMq2Sw4Lzm5iG2Z37mUajdvMf4aemR1A06ThlYqcmeQx1HeoqtK4ldFWYUgaAQ4SQQdk
4bO36g9cZUKVgyM2yOpbWCInsG0aM21SKSgOt7AsIV6D4uHJKt9JtFTpTPxjusEECgpcDos4bhfY
s+0Ymmox2fQ8zVv1tw6SCaX9vVeyTOnN/B2lVDowtmmX/oHq2LOU89uahWhu12BqhVUpXeN9Gdw1
Y76eI96gzEuEl8LXNJ4bU1lJSFi4NAUEMPJre+yl/yoVVDqrQ/us5ubGWyeF+v+BiL3l3ClFkVFx
8tKpKSVJ6fbFaAncw0JZZSeakyF3LL5gTkRFQO6ACvvDHA8orGv9dw/vb+Gwm4NP4f5cTqVDYw8P
XFHixT6IHCIn6KtJsyda4IcCZzAZEWOPT/jpPcPRW8HjrBd6bnCkW4drjvt/TrLJWvJhLoRPkCwb
Oebzz3ennMwYUpK9jHOYyjlE7Wm7tkp8GawJDjZu5fKtll+xrTdvba/VeuqJrx0FGI4ATxADOrOa
k/o2NuqUWBCoSf9bLEkFqmXzAx1plb+pO5L3T5lf5ecu0URWr+V3eTjmtJzeRSeXltpf2TTUQEYd
VCUFfu5XZv37FFdsVKNubE8ls+XNPEz7UyBLlGYW4Jh1ZLwVxfBJAVdTbtYb8AID9zyN2VQAEJzX
p9xJgvE/itUFqvKutXn9yxqPu8UluGwsAQQxj7r3YGyLH0tQNYeFR6kwk5lgYeuvZYNKReA+ZoTe
LlGTToQTi+vJqpFq0xpO8ygeqCXsFJcAeOUfi3fcaNHGOKDxT+zLkYEsrOGzR6hmXL+jBa1l1AC4
JOHxgyJb1kpRjygHmFwL1Us2x2DkBIX3pd6S/ZVIk9sEKbcleIit04ogt2P6hOYM/sU/3gkZBxvi
pnsWbxn1wbHl9kXRj+ZsCR14KxaSGyglLItqNGcMC2kTp3S7k/ZM/gFcI+PP8N1od5EO/InaJcr0
C9KuZYNYASQsNX7Xk1P5HMTeNhuioEQWURqn9mD3g/mreVyK6Zr5u/M9L+VlP3EN2ch0I1G24Xpb
C3tqzx6W2wOPTEnMNRdPu5UYVvZ852Nnkps9bOVktPYnthBLt8kadua3DYAIY/pDFceOZUGXG6nz
KRSRmNZKxo324qmA2CpmTiJuk9g1+2bsXHeRQZLWSi0VB276UM6yKveWCnFJ4LIGdU4R9V3e5Z0P
sD1ReMvogg8x+aIKC7La6zBO1yt+H9uGVhAI/8T7HKxEHXOIThFElIENen97IXujBb/z+pAFpup3
OCDMWmGmrfQSheFnoyUOK9UTtpoIUuR6mUAKb2g/aLZjzG2WrG6nsCMxH5EpSJROelPPbhuVe11Q
GE3hpX7bswy5VLh10INcdnanM6FlpdiEajjNsqkVZ4VHlVTc3AafwoLDWBqZw3o9n/EbsxSImSVE
724iMEq8wWi6Qn9HTTCQyWk20DklCbuoNxHE6Qa/9B9rRMdgiR8vpmMnEMetTRsUs5qY+zjyZm+w
JV6lU8hcfGaMP+3P5o4kVhpgEB0eGN+4ElL13/Eordel0GQ/bac9iqc+qycLJ7oal21IEKmD16Ze
nHp9AkfT2+n7LF7EPqZBTsBt1OwTTTeLuZqDmLqirlYmdtJGryx2zf5y11GrJRAua/rDjIQBQ9n/
6L84z/8bvJx9VpvY3Nau8UjV/KIArqyC+folIQ/EzAhAL5TYfupS8Qxu2SS2j8sS82spEEothbDK
bBQNl6/EAsrQk3stpiWosz88Uvef0gG0PlWB277/BXG113wRIVpO2YsH1KK1X6wpGh2dOGmgjtEf
Potr5r67zQSrwwIXAJRJLpONnN39g/5seX4OLAIIxFMfCTkdsmOCGJ5YXGuUwByg5yYG+/nAoDlj
4swEo2VrHl70c4R3JvKguLmHwFvw0sRYWPu1VY/dLyc6U2PG18sNMd6BXubo9yJInxIViM4ukZ5G
9PkSlPI2O80stJraVJEioQubV3LZY/NNA26Fi2MBnzBLJ1ba6h7l0LdacRTb5r3fiBuvU0YAS4V8
DS5emB8blQUJfu4ivKgtpPCFRF/Cx1lgRHKF9HecnJjxwDoZlISlaRhDfcsPBU5OJiMKwQ/Ai6++
yM/dMYH4jcHLKKTK9o5dlptcEe/yp5C4hVBSl8u0DRq5g0Bpc85OX2H1ko+N9W+TzraPZe8IHKA9
nCHhteQiZZmTYnzyNtzmPEVllFth2Pn43np0eJ/mAn1yobFJh8xwY2mItSjy3Rpfh4JPyXFHrtL6
28tmMm3P6DlTW+yIefL7OW7aCPDrbls4mpo/ycgZcz8g7sTPw9Ys3pttmoLIpzCF7mB/bSSOBlxk
lKqvz7kkbPbdsOh4zvlaztZHpSJwSkjPj/54VNX/DxEvKsrOHdyTgWEkAWbFVv4eZibi1TxaxWec
PsJ12CFw2muPYpB/HiLwmnk2DjCcbLM57SiHgpV60N/3mWXAz43ZBGr1RFr27aYOZgTgCzPPgMyK
itbbUOqYO56vUuULRbNlToUKLNy4JhdNP0j86mu6jwm1jqDq1LtPrlWV4K4DhEPiYZrbklVzwiY0
CjkX3DbvyEEUGY6w+1+qA3llBsJ47K5BlmXBlrvuXY6an/J3Rns5ANThCVJZZnCDhys1awuaHkAZ
dBlmQw878AzYdpcNl1glVFM7zs+q0zv/E77JmBXFj1atJFvmbVlAaCrlFMZUEkZ6/F4Vd3mwX7un
P09tfe/VwHVjNG1EskUyhMbP7DwmnqwcQ7+I5ENnrYED0gKtVdnAFuXJv7XyeayMMpbvFhDM+yUT
NxhHENNaTt8lXFTfCvcg8+YV8GMWd67+1wBjcopFjqxMiOLZl9unaFB3KMgU1RuxDWf4fItFjeyU
ll2S3mtJVJsFrMcf4YhREjTPuUVvqCpwotreyF3xlA4HFg4AhLYoWzWjA4wF+hfLx2Br30deKxVi
CllXe65wqgUOGASlOhFGaeO20M6LRZCHB+IRfVW7GPYGXaka3qi0dI6fGJs5IPSAVOtMyH8Zg5Iu
eKHXCzq48kO71oWFmzonN+tlsKBjFcJfS1WAtpGLwEOybGNeS+sFqBBiy3ZuNq3aioud2ekCh19A
hdSHJkRLULld4hMuotM+5Q8HiEENDGpzLcONkq4Xs86lypvR21VnP2Nay9yv2d8dQ0SFhF/TCGtR
0Y+I2y4oEGXOLvOVMyD6P7vYS9q/iuGrMM5pC6lP3OoRei+amoAFucyzZYLA635owUxrFgnoFfdZ
XmsDk3+7+eKTmmFvtkZ4I8DsAC+I22LyOesw8JnYSHjPjxBM9rwpTAQjIDYG6zC9XlrjFGJNcP6F
V7FLzyLjntghy8lKh7A+bnP3pem2Ea27oIW6i9HvNXxhg4ootr8e2nxxD0FnNdxWVq9vVMoNZX00
SrWh36Dm92WOoVJzPmXLeqoVXAd+N5A1T0yqmW7EMx8O/wHoGigcVQjZJYjF1vDUUPfLjvZgE4we
bjN25dt6LIDnNRzhXl4CGKySyW1VhAP3fQOzJabSDDirV3AFpgJaOw4PbNnVmYEBQ3JyWojawVqc
TlS5MJwwzOWPqnIr2GPBeJJIrJokzOkT05BaIydAygyBWOs9rxsQM3WBOaqsTdGMG+O7XsV64e0k
wcZWncAfVmfd1+6GyemiaaprQOlea2J8Y1pmb8Pf6omAjPsWg6zcOnaNpp2KVlbNhZNKhKQKQLPe
74b2KPYv0Zpx1hfBQt91wF+gOwEf9h5Q2SaEWreGNs16ARWrpapUZmZ/p+jWOyJvvLhAfb9xdTW4
CtwefhF1wmO5j+/kZjHK325AshMFMBU3+kJMyPhw2W3P3lqgKD+7WVxkvVWECllOqwqk9hqek33z
XMnEMmvGnSgjNO72XPovAKU9J449RORgJyfFzEvs9ZT2oWT+mLpvSq/GFlPjDfRt7P/FXqB5bjkZ
bGiYimj3gBGfQNdH6ye5J7exSvRUWra1S9haaaASKq+vOBMi6ubtqTB55GbwT6wfrqGj4yv7HWDC
BgiC3VwIjXv5XjHAnUTRjYXYG++fZw+F1hQjm4CzHjFn/gzQF0rM+ret5Sb8kuNk7iQgGJgzKK/q
q51OlCRrz6jlNu0STRw7GfVuTG0GH8q22bLTg5hyHhK89dzs0Od5/mk9mc91gT48nONvoLIMec0Z
LcYIuHfHgYxLzGGD6sBDan61dq/i8ebWhY3MThhm1fM44iv1O/TsV6MCJ1xWR67hb8KlBVrAtVWg
pHYa9Fd9d+tFt0MMd5gAbDc+I4xbDW/x5fXwaqlV8v43ScrZ+fpMUFRRhzx0TfZsAdprz1nAvC5z
CJuM14VVRcrINSlUsX7FhMlSdaHyMAg3lEeb3UN2Y4RoxYpi14mNKPXMvPUB7wqPxeRMhglMV+o5
MOKAMwn+htCLWp42pjALuG1NS/rCYPD6CJITKpVkTWXcxngfvJkBW76H+slLz7ZW6HXNjcIivR6+
EJEuyUdJUyTiDrK3nORzh/3/0AuVWFKGOjt/9QO2cI+HnElOfKgmVvjxjDw1HqBgHkmj1+fbS4mL
AhtEpL/TeqlHwXl4BWjdoVcpM/OIofQA/Nv5c+WJ3U9oVWcBylvc+fA/y41LtmRa8xgwBeaFP+Wc
zr1C+emk0TRsAj28F6uBuJovlx5yGjTWvd2XhoqYbbYO93T+f2UWn3Rkc6vS01jNW24dRkWnxnVZ
KH2B+9aMfS7OLvYAwdERovqz0iPQjwAjDRAJ1L/OKv83EnNohGxehnKFzHzd3O+wer4MMkMj3mI7
X/7AcUUxrCzuFSuigFG5vZD7v1F6x6cXf+wu/wCC3FtkUrDXuzzvUIPQveK9X4h/p/hjbz+nD+r7
u6zJorKJyPzdL4N31KCA88DdF6nK44nWp2q8uAh3IihbdRV2JHtTIdK6WQ1oFmnQWtg+C7IDYeLl
zhjDBXIipdCPp8qOBuF4vDxQ43mbEg4UFZzoejj5VQGURHWBs/n6jYOnXfrg92im0ORtZzUxQ28V
aphEo4hWp1YfgvryXiYdRyJCSHRWKPsuVAs91X9hH8c26foFSwLPpJ2O7gliwJPVDBUXI6Jqrefn
dBXR4STD4b6UfH3HcZhWQnxnx3qP/QrgSHx7rkkaoA8/HrYAq99HBCrKKP1rloAPK+owoPG+kyO5
Cu5CVopaVbr+oVBh/ETBCSn2tTvCKIjmRc+H+2B1NgAjjWycKaJNOLo0lo+RGfy/0BnpXrcQFk7R
mPnHsQL0erF9gHUAInfQLS5FJZ6rb7tE3gy9pfW9n/N3kSCF9V6qrvUS3O5yKzrxTTvINyMtGasv
Aff4KYuy5vC9VQ+8a7dIRsStBgjymVXchZBC4RtCqjXW5a5Cz9Sm/PN3nTuC64FNMPgVYQy3WkFq
dAzUkQ1uO3qkn4vfx+NIuA49shK4TWHP8+RXZlOdERvrqo1pIjATpxaIuxS6PqhXA/NtMOjSd6Rf
PCcekw0fYeyBWkLot+VW9RZTUFQ/YGgaK33Inf2b7qTa9K0gj/+xPKR1CzUeaC1J+pEWaR3iNgHf
veH+wVfdan4fxIao5X28pp+QZ0qiLqSO9gN5dqIPYCDvZU/9rmnWlqQSog4UmiZ7u3qnZTYfcxNQ
XFBXyjjQzGPeQmp/mHKrGqCtsgjIneCyMeyfM6Rm3+z8rG7NSyX/vR6adegtYTyyKpAUdM44ZCpe
BsivG+GI0CbD7hpTY5WLM7twlNjszma422X2OygWiOVu4iOO4A2r8gkINE+8/QPQ6ZF8vpZQNMLr
bkyStf0z0xJeYZ1RSwqYpJUbsObMrcDcw6ZGQQJt0dAp7rUXocsSE30HkfKBY9H9kRLZWLLiuaQR
H4RHXioxpEZnCMU7gbRUAcVOUTJMyVXz+UaBO8iuZPI+GudT8bf9Q/sdo2RoQmjoIJ1bc9E6K+g7
i21MTizyKtDo8IMyyKoo2y+4RzXRsAJ5MJaaB+yhULylHbrWZNVuEPPRmtEIgAbH+GN4uUYjzr1B
n/q5v+aDJCi0cjAuYpgTyMHxxGhRngfmtSTBJgSueHaOdoiu9lNAjR4XQTOTAQsmgd7ltkBOStKY
FJKrJyXLFaFJQbPWtlQCMekWkBqLjuWNwq85l69+IrsuN+S2RPCKoPGdIp1BmwyadUXWWmczY65A
xrFMRUJe/cOughFbzy4XI0kx2plPFKof64U9yRX6p6Lm8Q/2niVr9n5yIh4vFWxZfErbCo1f/q/s
HnoELG/x3L7BNgjeb1NRUopKV0aH6GcjslFzxPDA2kCW/hwG1ggTzZ2f4ABa/0EcVVCJFy/sZF3v
N3UfYFnM2H1VYggJ6kF7xLnOtI89dr62DSLvxcwGLgfTyHhW4W02US45BEz/bzX+z11g/UD/o1jB
gsn+xkMdzXnAE4S73as+uX4IphY70iArwNSeNOuMGtOGGez+7SwGGbf8B2nTPRS9i3UZrLcLFWvy
zzaRbt8/I+GrlfbpG+PQz5Q4AlM08YHrWRxrArmkiXT5v9UF4loMj1miltXIdDEA4/pStYCUGbl8
RPjTg4l3UxkvixjAgoeBms39PnVwbaJS9T9R+/iPJibhHhcKVrsIfDPa4zZO6Sru7ybEp1kxE9hC
gfNW7PN7i8GVv70MDMGrMOv/S9G5IK8T1eSN75iE48DOhc+B1w8Ov8qsg9rN2CfhrYdiIYBgLlOQ
iSGNjLpPfRAnPjVuVr5pZ18bkVGxlEPTWWQcYgpPqB8Jw1BhzN80PToUgrajkJPs/QUlvw4C7WCc
CBG/sWz/70V3s8+wgi+gShNZh9WfJmp2MxZeOSarXvvku85+4tLNwrm73Zl2++y0LfgvlqI5A5SD
i3tCtN8JVtWNtirwleqaAFuuxKaRJpveLGRI7+jedusnTf24EpgaMcWb651z4GFL7mIh+0ijJonl
TpYrU2etlv2gE7wWWHmwnJGw4Rt+0I6ibKOHweOwtdpSkvtiT+xYrT0KrvbJ5wWPBEoJ918eruxa
ZTYF4YjxjjHNITF2biDE4sRCbolNngLprk9sjcL2sPskL8GcmHMjwMA+OtqgZ+uSzcxM8H061zTG
2ybwqlR58CVieCuQsH0PNfAMZqv5eSCXhjTGkF0FIBm0kFsUxfklFPt+GKF6DURQxnW627oWVmGo
FtX6enc7H8o369OC+T08RhHbOHVJNtfQ678uMO293OfTamZIrxgjPwaS31v7gArEYAECt/YjF6o6
zmmOa+VeV+cuZbQLcSLF3lIRPuHx6YoScqtROt6HiRSY8pFg3GXwDSjhESrVXDlXa/oZ07/vRRT2
JPGZLwvCMWV3PqmFX4B5BYVtRePs21jKMMqTblnl7U3RImnmKFw7rjHk85L0Mv8vbgX894VUWk+1
6cYyEptn6BHz4qHignMG2DZ9zetz5CwfrIJ4b5nKLeqRb1aoIf13HTGm96u0Jut5wLto4JjgP+Ai
/WFDbtFCqfpg2pOBamXdPx8wPgmfX7Gf5f9oazqXOJ0BBQsAzQmUNJHayWIb/3QVNbjWLsxpi4Ux
wfMTZBsEjQ6Fm0jZWEkFZLWDCJ9mnQAKbLwa6mMStyfUz79fS0qMYyAwOYB+YzymWPlKq+DVkpAb
fzjytOcDrOIngxrVL6OkEkmx28KJUr0tQ/HPugLF+DGHtLfrPsCDqEqcQrEeHWCIrP19KAUlL7kx
wYYN6FF1KUq745A+rhoRA4Lm6+F6NVhdZ2iU1oiFNWGLJiZTeolDQfPQvc48ZTiH8o0tQhcwBpdH
s9Thp+SQjxjzYEJV9Pl41j5BbWNDdnUNNSWTpXqqn0lRY/lnpbD9Jev2s80h4GbWp8DVwIvC1kz/
zU17JZvGpV2NcZx3Jvh7BPm/mL8HUiVuAbFnY0z9wmEMsVPOj/td5xX6j35Iut5K7zwaxwkPFFnj
9vJrwgLtoSdOeJ+MCMRUWX5ekJsoxxO0p8XWjZyMfnMxhvyfFfhMzxPtYUHhWybC2sOLFGiQfhBK
37X8m0yju6ElP8UERppTRYKHIaKcQPQ8x75Op+25bFlEwj2KAdqdaDs4GjaUIan4r59M9wLhOqz2
tTtb50IddoTrXGkB/EZnocnTfa9ev3B4pwOgiSDAg2Ak3+x1H8Fd8AlL6+pC1pLsBDU92MeV+D+r
1FKm7sSDlgvbd9Nsw53bAWJIoUpbKEMBTOSxdTCDiduyiUXjSX5Cur1+h5k+st+W6GJ31xDpJYxg
MwW1G5nifOgZZTFcRs6b1rC80hhndGXlUGr170jnDe7Fvw2MJOWLPP3a8pDas1DMheeSCWo9yIv+
R3hRg9XozY0ri7Awb0zK64VyBe6vD0BWI5yuPxCrLjopy4E7p+yHNOV5dMp+ZvIfNORKxprrG3Mt
b71fuybBcj8TFHZOrMIkM+XrATGzD8TgpoJ2QK1D/2cmHutKW3UZB/Za3sLUsZQ2AkGG1HRez1KA
YMxJz9+qEe/3h0DKb7LRGEeVpdfCGBFjjM4CWbq+VLx74qfAPF1GZ1Jqthow1aTJJcdiw+4aaJqR
VVbel63qTsynF3/xa9bd1iHlZNDrFv6OSy1m4u3ll701I4dc+l3aSB7NPq0Zh/jA/tZSMhPjOsm+
8bOU0uKNx3Ckx5lZCqoV1ZuzOtJEXsv+3nNokLwisb0NOOIlnDgwXoDdx8DR2p+VpOuTv2MInKKd
e6PHa0JMAmRlVOIWzzodtNPlvbgedM5pG+5ebfhnzqt6EgDDN7xE7Vtsf9l0rcgaFlX3OHh/A8zT
+0Lk3ucwHVxyloDNSufPCH7eAqsACwf+j7CHOAMnWQLZGJb1vbuyU4ppj9piMDRUdalwOINgvUBz
XdadXqDK5yvWxCbUyapdN/8teZWTfh4PUMQepPsmrLhLWnXR/mVKNTtI1VVPs+FDQKCtNhJj0UUT
J+P7gisYm+ULjEhsC2IbnNn7h47MSDJZgNHMvpXeSJAvmxZLfOPL8wlzGFObW9NU+mHK0ZHUqllG
JQZv4Kai6X8XlqXT9kQ/JrcA0nfbyMM8z99M2tAAPj5a4gdoQw7cjKjqe5+iTPHbH0ReC0gSlkhz
UkGYJuWnY0LA5zAXH4sh9xbwFr8F7V4GmPuMluBMvsWS5MBBMHjxTnw4G1jOX7gNwyjyfu4TF1Sn
WVCDua5TWQWcm1GsQjWhX5falRJe6+yADIhMPuAbr0JzAxkqorl4WAOljxDYSEQu5LHKNiHuDgvf
6IerrXbp5DD8AMUipsDxGSrtNDVfeR+qhiNCZlNO2Q7YYFdXY0zJ5F2rkXkZ4Aq9XY7DsCrszdUT
YHzTl460tfI/xqdS15NTkIM+Jcza0UORk0acZoGYHRdMlsvnz/E+vRMJXU2fgOX1anhOZ03Gv+bE
P/XqxdksqNpMRoBvlaXeoroKaMPQlNfPZRo3JuOakPpKPCRItEjcQ/sXiRFOQOaHjcv6v4PQF2JY
vJQLA51lKSEeajLABCeTfL+2slw3ZlVri+P19btApD4VEcx9xjpKCS1Jt376mWGEKgdggPYEmPhj
ykqkYP9pWxDhRD2WexZnhQ60v3439D8KAmzLlfgzZhTCSNCAaZ03MwOUXtnHeZLZRR/X578E6Yjv
TBs3UJL+2v1axsVQGhyhcNaZRDXtjaJQMqLAUtCJ/AwjboJOWw3cNaErZYNW9BJgZ5hDg9TmQDI7
U3M1KeUPBpw+BaDWDoYKH4cCxR2q/b3wJwaX4oaQntZO4Au5TimZ2on6CMwkc//EGWzv9V+bh3kX
U0I4QBy0AQKxm4166SR31fBVn3elEgDsDMbfiBFLlHgKgSYcUPT9egks+10kCg2np98qVoOKBXpV
mAxcsxksHDC1y10f3nrMc9CebiK59VSv+6cCZoKe0JLtQ5Cms1r79phNzZCg1sTw0rN3Tc9nBPZA
rXUMG3Z/uFiM8giyr1BQCN+3I+6QM4OsJSPIiiEhYKvMM8kQMA1BW7vebPICL0+P6Bau7txdA3xl
80ajVXTxP8tNmcfvxdMQvVHNe3SLjprzEbbr/h+NImyhJXst17nO/0O3EjSSa45gVxdeYVRu4F1v
72AvtRoAZHPgslJKgCgDC7KiAXUFIUiP2m0mwopDXvoXuptGaG1wqV7Zsq7HRSuhNljgq41S1FRV
NKZKFUN1zcHQqZhR+E8zX45vRcZkXsAtc/Z95Q1N2fCYanXHC24HAnOPx7V16QqcKQTxZ0pPk2vS
Fc+AwBbvEyu62t8hqUPEh5fKa+AWGDH0GRbA09ljv7w3/uvic1TBzDMTOYBWeihoRfOBG+cwEWgv
sJx3YJnTvKnmHrvhGmMGXcybPIpPxteRu9rux6vrknu5u+7Adxcfd7hQ/v8DuF/61Kxbt8p1YgcH
GMAPmeEChauDpVDJ7MY04rS73MrYiiBzjewB6u02wSTkiejA6C59qcitE9YoPo22x88g/6YCuraH
JtdQmof2wZYxIjGIyHDHs/RGKUtdNawP8Ed5j19A0Dg7TN1mH1b3ZkPmDXSpkrbG9Nu/bb8JVhM9
oDnNS1gDcxEeWnzQef9M9vmruvOhVaAnALL/Y487Do7jJBeZuojjQJrfPw0hcaCpQjN56IT6mOZa
s30aLTdo/JeQe3whS+kMnHSngJIOXmIDg8+G23Y0WyLbomaAxtcUZu0M86mZZKa7EKtv64XaLRPj
oyK+WRgEfby2Di271mQk/RdyWXkQmGzNxCbF+uB1CR/EKdWC1c5pW+LPFO0rGsGHI+KcjEG4KDDD
7ERoaR6vbImHH+lAP7q/3+uZUn8wKEiyHUP8Hn0KQB6F6GHTd1FeRArMuTY/substfxzWUmekRLC
QJQEPMgm5vBhVP9qDak8iLw2JTiHgIiavagM1YhdDAHQrI3KVWm6ehzCOt6Uuk62RnRoYOYFqgR+
uxdpn08q6F1Vvw/s7PNrB3wSNrrz6bI3/cZ0PBgPS9uDmPs2d3kK81v1Kccaf8GnECFyMqeVPXkH
0jrSr1t50MkUUf76UTDLT49i7hFfY0mXP/r36cJomDiamm1A4rJDzlJ2FrPKT3NlTiEQ83AKA63V
Msi1nRqq/27Rq//NgsJjhxiQry+arwn73Mt80t9wMhyscfOLXyPKvqMY3TUTYXS9F6lsbZIqLamS
PFP5VGQzc/Lp5OaySchoxifZWyumpby4NcwjJXU0JmHBSDwf/WgmVeKGiI1J9hqsy0XNw5SeWcYy
TTQFqg7jzMDAXKdKbLZiNP57VXcu1TbJp8XLVtZl3yWF7XyI2Z6WSq1GISMiSBW4c9bf+SaAXC+f
CJGJgqHVZZCczoYLaKc+eT56oynNM3ZrAJg14Lzqs9BskuYxCpuPm2gzAe/RlqDYzsUvDyx4pyL1
7HAwcBmnL96pZKSOCYdNsLKxlYzXkf3AexVlWlUM2epg+hOvCyiauQ5Vy5lU5x0VFCyBjC9Bj3/z
tthXSKDnWD64sRCo35VUEBWSRwmClERLtNAVUvwcbnhLCCxo9axoZ1FJcxcf/SZGIGzI4C04huXq
jDLhy/YhucbiWPkapByHm9HNE96J36i7gPcoZTQfcT9HjA5onCp38e2eF4nYlaB9hNdCxleMtTzl
hD9gVOFXy4KMVmoGuBpwlj1s5Jdm6paDvuENRDB15i/hULESmvplIU4cMqIBu6mzFXx9/OquFd3l
7pte1jYfh+MuJcjP0PHTMJhSCody6/1YZLVfM3GxiAtjTdMX4oXJ+ZzB1Yc38BTl1SGEKfQoUSf2
e9aDGOk4BXYiLHulCHmVOrEolfHb9bLQpdx7VWjxx+VqXb1Yp1qQfd37FEVGAvaXVY8v+M8MNasP
RGhJz69lP6SgPWAbkWxmXKxQJx4R5zQ4k2OsLoVDeVQVEj/f5ks3OkKHdXe0eh/wiaGbKWk/zyQ7
5Qp6aL7iiXnRrBIwXDu1djmmM4YuD7C3YJkJVgTbqM6DaZz878GEDtupuwHEI1Kb84gl5colwGU4
Av+vRhKT+Sg9NO46d44uD0fWJv5mh27YcTi5jQdGeaVib2WhXfANQEfduiQe3I24oGrIe6ffKRp8
zkfARPQGj9uNFgpC58cuCEYQibDOs1a3ZDp+0ylyyP840eC4aIONe27ulhRmjD645q4w4v5J9K1w
C2sY0jrw0s/ebjvDvFxNzkmbCAbvRZL8xQbMsRlH8A62syOSkGAsyvn0ZKRSWtrh7twmuZ0FI04m
2pEeTNPsaXnSYsEG5YYlY3jnSmmSnaAVK7PUQOu+4PzKGBY1fiS1g1irPtMsn93ksbrAVcZ37fR+
Rjya8BK6p7a65L4xCOYrFqwwOoBlPA/Mo2yMZGcobl5pYeslCTulHcCCE+Q2+SU+TJu7tWO2EsVD
Bc65WflgrZl+RCLSK6nx8+avTXmsX3MafNtgsGK6FZYM6iqh0QGCz8xm7n22p9zWK2eAFsvRI79C
gm5ZxlbArOwS0cYgqfp6AGV6J2GsDWlmENdjK9fJRrEk2x2F8DtF3Hb7Mhq6ZzNnZ6TFO35sJZ9/
P7LB50/T2VwW6nlgp1Y5LGwd6YaCGaP3/+llk1ykqiE/TxUvxxvf2qM1l2yMQO1Ri/usuv3unApB
ddXxyHWVhrDlotLHMIPwEI4CPJ9wsnzb+2HYH5keImhHm7cZTa8IJm2diWhkMbbZI7sNl3O3/TNX
Lo00zYLK9Loxc5XJSmtLXhiE6GvjvFjBNaAh1dc8WKGm37edP5mHA7FqgAj03PAu84DnAZjBnl2W
wQ7RAutaVsVXbnXYOoNNy2W9oNLx9nZxEQzgVteIKcHbrCVFfz5fCN8n14CRJozRYwr0AHpgZ1sj
UN9xLGwo5RW9F9RfkEnSP+XbKPhAX7K0p/Nn9CTgIRCYU2/2l26hN3fs5oFDU9oiNjnzWWRqH73X
UNDq5z71cEJpRe0Jxv4oc0UcRqCuz/5p8+XJ196wlrFHXpSrPzBk7GK+4A5qml6PCmGZ1SdBcpb0
xE8VHLF9wk5AfSA9BqSO5D+A/hiizba2sSANd5dBPpZwLZkCNQI6CBD2/m1/eKaSa4zsHm7DBTUe
EZOxrxKa7OwFRX9CvXGbzyZ3jjMay2ltnaB0zyvOBBXehNVB4JzRL02sOT1pKOc8lbmWb3DBa96h
PpUJgrzVKWoJ5iFt9L1pODs0o8QE/Pg86bCtlTlWizQWXyif87yMWw52L1q0mZCTHTJxLMwDsZw0
4MpX9DJ1iKYc8MhggNQh5xtgP3YRRi/cSv+M/FnZzt8KRoyagedsnrStqHMXAouC/o9tGxQY+gD9
JE2BqcYNpxi6zefBQH60cZjDtRS66u2NoswtACBepgc/Zj6K/bIheDBcaZGyLKeUwjqCzjjc4k9R
7RC/6loPm80eXISJPPvYVFVfHuhDBEDuGlWd0Ff2mSzyH4jQUedc4i4MpbA6Uv74rpUCR+JVbK4F
8GGZiwxZe+Fhm5/8fcuVTfWiZX+w+Hwh9VLzqGSA/PGsObHD6Li/tlNMf7NF3dQ8AdY3OqbYEjPx
MhC5i9F86uLm6WQLhq9j+/3x9Cg0LeiHfCkmnsJFbpcqOSgTbztTJoHXg6KOar2fjCO8ngO9xhDL
f8lo6cYF2MOZK2evvXd+BGIDQVpesD/wdUt5Is9bR6lbgUVe+y+CO0cF1bR1FpKO4Fmvt6hcNjbX
AI7EgIiJujS+uAiNgQRgY4hkgHMp5PDKKk1shHuoHk5oFQNA1RCf7Mhi2nsAJA3jnWzse2fssq0L
sXYnjgPMXe+bXw2jmbwBYB829PoVotkRSsDeUCKPl8GohFCPPm7POct75nukf8W5cWHqq324+1nv
9jbyjAWQFm6RKSV3AvQLfQerU0X7jy/BO2tJ5rlRSOT/LVXx2opJswETW8lPoitN9PUuE3zccBuh
lY9DW+iA0J5huGgJnlBK3dyLkAh12n+Gsr+3cyY82NT1E5n9a2YdoajkBWAp3UnOY5C8rc7+2d4I
iUIO4JZ897+xe5/80FKW2xU1zNAWyUQjEXiESeLp5IFaa0g7TbgH4rdkTgQqQlA6DMItlLrDCk4B
Ir7H2p6sBNJOR5O3+qmAPt84YxRAQ8wbmC3zIbvufMwAXRg8DZO2ADVy101pZZ5hDe/RGJqjswxe
3p3UQYe/EvGRIgeyQBcVlx94tLD66XhoNL7374DCPPdtvIVvq32TxTbElUabppPQIswRijucRjf6
BQTlIkrB5J8wbHvpBxnkMGJsgAZjxjKpcwuhg6Gm2TGbEFAphEjkz0qPaq8TocoQ8B0X2DCD8OEr
o+lMyF1ljGTfUScRIonOr80H45dgFvE1XQe14/+UcXg6Cs8iJqs0RfMoHA1UWzEEmlqNoNNPuryi
PkQW/1cb8IbifwEzP/KM2OPvOTWNmnVwdHLsv989dZQHQ3OvyyPQwpiGrbbzoTX1V5cThCM9MjL+
jn8u36MmazAAilPZklHfa1bqisgWLNLF7KvFLNKiLrcl/hQGlid6cP8TcEPjlQGgfkbAbKFqUQsv
wwedfjSFc7QJr/Iystg0cJgQGwGhTy8D0dlBHjIHfHn4ziXQGtYxG9ffn0q8ixtQRqSUlWq5S9LV
GjLEivcIuer6PqAz29dZEd2U2wZRZiHT+Dnx7i5UDNvOth/LRBL927jocIyOoSflJAX9I2FoC+Z0
fIcDA5eVyMssC3KVm+oNA6dwN/BJRfjrCi4j3Mx1vzZpDIQ9RUTSv7nHUxw0Dm3UjA/aWttTxr/H
yXEmafao+rjvtrJnibcR2LNL607FGhyJnOQCvkec+mMcTwsHCEc8S7rATNbvw/XKlaUarX9QIs2t
BHDWdvCfheAliXAXHIAhLB1kWKZihDP3tPM3b91+ff8h1/6E6Hlpaut1Gj/mpwWyg0p+yTB452FD
UWlUSvHi9iWw7qxC1u+zKIkqHTbKhB2DN+SRRV19VUtohmSWM/lzxZ9irl/IyJAIU83ReiFq4RqL
ZgCcso6RHtcmogcNbLzQrcZtqPGlRfxPuvwUivN3axC47jN2KT27ny149EPmo3atJPdd37aJVoyQ
it7izv2/Afx+VJVgEqcuuqGdnIySPr2UPnyBDk1TfzshdeVEICFJvrfHgv5rqXj3fYJFBznzovvC
XU3qGaUJupC8OeOGqf6Z0THwoaBsjhZTXcD7udXGxBVZnjNdcyIGm8U3NmhC46C9vshxx8dhhtwb
GHOtQ1aIaVVKhdeRpYDTX6kC9rzR8tWU0uzNKjCdqb2UbcRDVlB50Fyswj7TY56dSBsXGo/PuM7D
zWqFdQm0IARU373K9iQfkoTWqHW98QkDw7WQ0QPukb+ffzjgm0ggxfFyhk0a3S6v55qAiiVHz15x
YY9zYeLeCqEBnZcDqNHSirpHL5DzC0TGMOfTothlCmCQGGqzCmoro+G6BOsi6EfhBJpIrMaQBUAn
JhTB5o8mdEfnFWq65kMAbT8vBhYgvbJDFOKislsxXBG5nb/FhT4Ok1q5/Hji9JcT6okOBXu+Xlxc
ygfQbnp3bzE6l/huXDegyvyf72eu9cvHdqyCOykituXTGQGWJGIbauGnoqZO9mC50w0Cy5MOByTQ
I0q7t0uhZ7xNKCuTzn44T1rQAQHbKGrxFNjyN9vGLSS8lSIByh0XdqIl+ZqkyhYVOEIBkYIvnAwY
FgQbBk8uBaZaeT5sSNFTxd/CKZQmhciBEBa05gTs9VZ78s8AfB7mVr5F+peKPeW3M+kcxxsb0vTJ
0xaRVsQ26o6aExDmCo8ANB7noSa0e1UYU+K6PVk2/dqsTs/ZzJWPkIMW4a0ghLO/LK9Ez1D8mVT0
V5EBTGOrJkBkhDSf+2Htd0xjlDPPDuM5Dlk+JWiL0HXAs5+ksgNOw03XKcfgwqb3WY2oLLW6EJr1
BRin7RqJ2pwafVwVeqw8vB/W0XkBnEWsRmKaN5AhQ0/IatoCzraQ5E2JJLD1MkSPItnIk/S7CBSg
KuuQQAatVgLOWyCQ2Vxjgid+nL2Ip3f+CKgU1u9sPSHjfhwrd+s6DhQQpmo+S72jVjNyH9aRw3ln
sjv3rFcR/NyIdx2UGInCbz71Q/o1cDbL5X3WNfxG2TjwY9SiBh3FcMkZHL3YhdQXylR36KFFh7cV
8dPAtP4bY+5PM8WCKiGlMqohikbIA7eiM5H40F4Boyu+iHyjFOisZiF2mFhTbiIR12Oty4DLMTGi
0g7WdtgRWUffs7NqpAcZgX7WgYu7RnRHumldGutZePNE5R8D1s4qw0BFn84YrtP19TkFj6Odue/Q
v/2wK+pwwXWW8l9mg2VyKGiMaJ0h/TbpVIGXYFPTV63/Zd3b3jP2G+sFh7txQlgSkyHyL2hFWdiW
h6ZuZWuFciMurQGY+iQyuN7KO988igsGrDlcLr4ZHqsy/IAdppPX2CP88eI/phT1BaebK/l8UPxQ
vQ+kB1+A6B+iLNUxi0Ur30zN9TL8txsThsuKVjwYB/841KvcVmBKh8xJMSHnDrOyA5z9uqhOmm8o
OFVywYrryX8RydggbHa7qWETut78tzg0zATjoibTkZjE/rq61YSlZCmRSv/0IKGRx6ZPw9UyDyIk
qAhHJaowEgDaBT/fTUa3JHxXY3FqN5buXdPSq/G5GUYGC5/D/YVIVlMzJ27VzElKrpxABBV1UUmY
fpq9tM8xN9bI5q9uqS/2tgXDHBa2PPh23dsoYnNdWTeoHxZKXtgEZSHvgE9Nx6iJEGt/I1tpy9Hp
VIedVm4/VpWKjyCRW6cx3A1YzL9nw7gOujcZwvjp0uwz/hFY4j66dkzkaYrXqvRzsT5fP6nKA663
vgdy6oMyUX+8TzAhmjz4wz617sm6GTjg0Ov+vKtaHEmKo0wWtF4ojANNKgB6BFuLkvTk15FaaDwH
vkvYtmG9F8hEJEyE5vUj74jUONHSM+n3GZsM1PiwnwyGdzAMU6X7Uaei/ZhinxFwJB9enXF9JZ2z
57YdefWqLWyazAqJ3UC9LciLgZv5tc7QhYhY+UcfBGlZ8RNTVDc56KnP8EzegFwM3hqqydXvTcyg
ZRzBIX/GRXyDMWo0QB3pPAUmW7n9FBqBQWbhF1WBtTEN0ehntxj7MdTA+2M7UyhHFlLaLzNtXfG/
Ysc+Bxj/QOF2tJ31SVdNVV5NPHxDuRTzfXpJAlwnua/Nho30T9J9swzqw0e2DpbnVgLOmVRAOut1
VnJYAvja8X6rDk518Np/IA2mSUIyNQGERIL9TxePtgXro7lnvy/6am12WuJluY3apUXlDuiE1J4a
00yy69JZXE8Z6sixGu4QXqh9jBlBgAiymCnnPDbJWVrCYSroJhlsD/zZBmCM6kEIPcMVEu4NsJzy
iakRPuc7ttBBP3MzfYnON013YZEiYCe46zhOWKDTW8v+VzOyRkjRjMm+KgDowUX5qei6IBxsfXna
8p6EHMmdtdesj2eOQJO9FRfDoVo8mT+C7khCoqua+qeNEEzO7Aj5+AM3/ckQx5ejg/hsDRDiHZHm
44NOb3wEWZN37D9tR+f1eg6eiOKoM/udzvYPQe/Vk0qpJgiLXs4FN06QC6Yc7fVFlolg2+wDvlsG
kFSp9+Uo3C0UaU9sg2eEGEDMAlCvPJlC5V5Wp7DXg7bG0n+2qWKT2xpUhs5Fyof3Q1oeZNbhM4CO
NBZVQsYur/F+X28vO0bTN+89E3qgkTz9+a7mS9jozA383wwcTOALWujTvwNq5DwjjzIeaHwY877u
1FxXSITnqem+hu+oo1IytKybzb9PxwxwMxax056OcMrjo91OKvGWK+hU3OzmeD7Nm1yR/PD4sRjd
ByQHyZfmokGkT73NTYU4Z49miZcXuTyfLLSHlSN/8qKoG4o+cOdOEZIZgV2ftcNF/XIx7r8CaGfR
BNETTGCQfvM8J1E7B3/kA6OTdFhBhZUx2BZ4YFIUMP/IOkbSmKDF9nabS49f2k7P5BplPV/xoVVN
CaSx61FOcRVsAc5OP0EneceFS3Xt2WjZaIMVfpL/9mLy0LkSfBu6RDNGlvSxFLglwi1DgZPk5OM9
1FVAbHTc2DV0rl1Bacy83Pv8a+4O+qOW6DONiYlVZHn53JbD/ceNpVVAEYvVvxZDbTAVcaaD4MbH
thc3DLRCFO/g3dyjOtaqHriZPYHSBBFoThlP3DH0kFnD4weh11Ew5jyZK94OebI34aIuRU8PiQXn
qtkJLFRIZ9FyFp/J7bffp6vpH7BHW+d07FpSo4HFKkl4e+0FXJLEa1odgVizWhcak7BMcHjy1dcx
Au+JH6FyQVXzp/BrHbYwDZ/W7L62EdPpLm0iIhpg8BoJN/rKJ0kGoE0UAsbOSG0/c/6/sUZatUeJ
xeA+Aq/S9UYLzKzy+ZAr+oRDV4BuemzpU3Z92upfWuvyfxAz8wMoyfCd4hVFtn4LJLmsfKwPdSw6
C1xqtJ6UnhP2KdWZQa3p7uZClxFhY0BlWYzt7FM8ZCt8w2Ovs4tx7293lY77Ox0+WhPyGGbttbRU
mfx8t4PJA488s8Q/o2jbjBWLW2+ykws8CdJMz/bVO/3z5XlEcQJH6xf7pttS+4jG3kBIT2dN9uiN
42Bb4IgZZsvbMupWFkgVaT1HZ9qAm1LeZko+A6ddpZg7m69vQbm0gyfZNt0I1qKsZh39zUnBukFI
+kDxsl0x2jjUfUiWwKokLvnrnpm7kP+y+2sYg0LcfS8g6o/7PHYQMUdJ7BvYDKltHcZ9GCWd5VuN
bVEr0WlJ9vvj7oUPZ8Uw+wj0LBcc1IZJ0+ggb0nroyUmmUKCBjuhQFADQuwM63ozfP3RmCCKZCEs
Px0J0EwxYsihQXfgyiK+kWjlt2sjmgskn8Z/BUu5wQnysGd4bXRxqPOGgxs98+VRfzstnwYtWv1b
gCB6+3MXbtKoOmotdXninY2DC2pc0Hc3j6V9dOJ29JKHgTjThlq2DNKg+7Zxw4LL0rZXz8Tj49DN
6lC6eYTP8oRTAQhLXto9cwKNQeC2ImmscNans1nBS+7mLT+X0/iONoVhiURmlXhckk6OrxTKSOhK
1NoTayqIUZm85MNf3dpQL3JEEGK5gOW+UVQ8c/E19YH/TUYI4fWjCIOdoQoh6i54yYXSorpbf88C
EVjS0ZMzR1TcstnrpOxelEfWAviwmrc7KKK1kLSApn8bPMXYYxQjY/GUZW0qd3d0WQuuXssVOxGo
RCIZi0KQAzbezNc7XfyjXK0XG+eas3rGavFm1J/kGUD7L8hNyHuIINEHzXrgLUdHFyklREKC3XON
y2w3Np/77FqR++1iIB7ms4j5kTSpqxKBiYyDCLPWO+qp1OHYNT5A/I+HskzKj0EcT7bDbMOLUOe4
j3fTgun9TqgPWsRx7vXl/8HEKnN872LQBNkwTjiQmT0SRN/ib+T8lR/6qos4CsV3y6miB3X2Jbld
gccLxUB0hCksZ+HsMYBoXogc7RG+nAW8/WI0L3pvB0NbgdleiOiTIT9W+m/37+PCiQ113AMo40J6
1YpFXdesUboGPfQd+57u1d4EUf9yeSffLESk9He92m87vWD8CFGNAVJG1njmhUF7ECXu2DmD8mP4
yTwU2at9wQHi5mojZjBp5whLXMnT+IgMo9JDphF21LNy9k37rrNBdTiMotuhRC8Wv7cBMx17F7lv
x4pj7IMcdrdXvqNPfjmUvjSTBdO3CKqaiuPnS0FmQJT3btcfCGKW86OS1yv1P247DC+wmktaEi/D
sGokRwi1arktuJjJSuvMn82mW0si/KS6g/VHi06hc/qgeelGy4EzWUjBDYvOcR14x1SzZmyvOUmp
50VuBwk3xobd0DzpNhL7a2h54qGwma6ZFvxHNj+i9a8fiBOtBt4uMP0gRrqlwEUj/Zt1GhgL/209
+mOoPNO7iJMfcEnh28aHLPz24krxuRpgLaEGabzuTKs2mtnFaAtHzzFPzfuDDNZC+ZJVtWzgd4u/
I+YSVTRBe7d2PU5TXur8p65MPRuK26vrhbQoV/uEao8Q5dA1rYpAAIlvsW5X6q+7zl5Wkso2yT08
F5St4M7HVy9fBXdzDyBVFNN8HsWvKj6/tjza79Uk1HcTz5dBfP+QAfY7b78H0Ci2qJ1cHCWEqgP+
AIJ5/0p2IrsAN7/hbaxHx+BUd4hkGM8eTqCCRK5KWJ/nkGbfyos59kxMkFI9rNu2EDQIY0CrC4ff
CzxmFLNT9dq2jE+2gucq/m3VQH1cG19g/dWzCZRa9Ng8OUcNi8YFNhblIkSaheVVyoCnR9Ts2ujB
SgoG+WONCq2NBPP6RonknWwEsPbBMbhlSysp87c/wxeP0PvBEiSOSIH9u//XF40EmjQpY2z6bOYg
wzYgNu1Q83LpO12KiGtxn8i0Gz7a6YvwzURwCmY8jmVghogkYu5t8hOHNU5DCkQ84vV7ak+Ob6Zw
+T6Xem5OH1NR8XbG/8BmsqC0FXAwuVQXsmeBpIPoYPzLWbIvSNu/2DnXlahS+1m3XjS8X7FBK6jo
oOTnBi+qU37MMhD91WYhya2welWwrBDkIL7qKJGFtbnH0g8dYChSrQ183JUSf7aUSBLMXWk0jqrJ
fu7mGa3elT2hr+SaYrGuMjzhMJD/Zi8xgqlyRclY8xP4LMxVl2j/KfoUN69QOPB7U6Gu8i1vsasG
L9hqViXAaSenxCv5uoyL/qwB52HExIzCdFe7SaV8dp9eazTTFUqWUlhSkPvfT1C3SosjmX7+pxUP
pEWIuqjtcX9YWdC/ZqmS7EAcA0PVQVQr/rIi4oz7Gad5u5h3zNlhSURFhvYO/XeSP2M61PemU/DL
SCCsDg0jbClJPQz/eOyDfH/gscj37AyWhrw/8KDmAg8L9sr0xCdkYy1wEt+/j+NCkpQWAVhpjIlh
yNzYT3ucSRfoRAuqxv0Oqg1A93hAwHicUOAbOWhcIByL0/WSSN5fXSVZAnv4RP0ZzQuYO/PBLX5J
4yOnX1hOVyDu+r8nbgqtbtksnLIiqsLA9bGLKtsCUjqMt4ZXSzjO83sTOKsHCi/1zTB2OGS2PA5a
jnHGTnFkuagIRF03Z52EOEtrSDeQLRR9TRClydfLac66fMT/xiiFGJs6g7sICEBUWmW8ZA3AVacD
7SQFZpwCGmYTDPl5aREFvlxUx37ElIChS0GPFFiNh13klK30GijAtfvSy2GZ0Fd+Uf9nOB9kEe+d
QLiJRQd8Wf3h1XD2Svnrha7oHJo3xUhm2lWsFvNul5qeD1U5LwWM+KB+8+CW4YQAlKEF43FG/T2u
X2eUigbZ4kQ1NxLCF6ZtW62Gfz6Ucw0B/t7V+cymRYaMpievMk00ce5b0gfFi3oIdJf19/IGQA1G
hmdZ/TAsqWrDHRYWEE+z8BZ3Ei+dG3VsxQGSUJhVdf6GmeBNKFuGM5hJGYLLtwPo2me1wYz27bpD
dGr+AlWPz8eNRqpWeK3tBAlwoujijI7KhY7ClKub1dkurDPl3Eotuzd0DH7msBVZ8RV/QIh3aFUy
1fyXxmzUeMHvqZvIe3PNTsUCUANPavA01Pc6sSpfQb3v2tCc4axx6+WIpJYAOWXt5XI6KsDcpDFy
LdcTEt4Gct3bGdd3m5mqrtJLU4fdjT9DsBPVxJTkZKCkMKzF22fA7AJKH5q1ecdVEWXT26MvpXp9
xg+plA2wfru05av3CPiSPcRjaBPomjX/+z+yNb8Nf2lUK4ionYE76EEQ+M37DdHokDJC1hm2GKNX
Zt6PcxCKEpDuKCsPhzRFCwstihGnGfCkfQh4SJL+EMFOPpUDeMvUvV1o309TE//RC/Bjh4yxKhcl
84FqXvO+i04GdidLKm7Hl1PLQD9lcX5eUzgTnPrPaLIjgrhdnGjxLvH+HpS5azljos/BojBRl5RO
JxgGPHpHZxRf1krNY2/eehiPLiJRHPMiVZ/qVl1YhGzHyWh+vS5s3P2c4sCDH3AdzC8c2zpID9Pr
qFBwe1TGnbOIePaafUUjFxrHbz4Nd6RJYT37uvBc1wFOUzJ6Dzqst+8bgVvScmk6nz4hIoda5dvk
NXt3mk9He22ImRPzAjbSSKRAp3dTNxuoy/r5J10vcsMPadD7LU9FIKaV8k3sDUC+peIs0J+3Np2i
N352xUxlA+jflAjKO9/pSLUryIPte0sutLwbEtvVMfaclUHnhqf4Oxr6wyrv0QjNYBmyZ2Pypg2D
nLJ+/mLkofxywuzbbcvimSt+l0AHvZYzSu6w0w8/ZjzB5kiOXaCUYUMGFF7AASShAvAPw16Y0Dux
stPXYvQ43ygfnqqmqgxXdF0cf2hPjtoLEN4cKQMYWmtIOyiAMXpxOWzBFuhN2TIn5Ec+0uQSxiEx
f6X9Rgida3znMKDzgKEFCQR3l8BjuW0je6WpKzO3bN8ohI1rv4slxDYMonpDD3cOfmscaH27442f
p/xt7CwNFe9T8aBZL+qE5vWXBVq9njCNAxvrEMVCj65daj1tOAj7QUU8CW0+wR41VYeuvgSSpIT4
Cix004n4N6gGTjRVavx7fax7/M8piy6EcedbHmqF1UITHx74bvYh3JAy13LBON9Hzjt1Oeu/L2b/
SDEfinMuvoEjoy+RQMFPLovJ3OhVfWPEZm+FRuoucUp1ZHu3vxTlNVzLRc2XLatOSjo9mjWSfPTk
07SOqCbpybejcFKIUY1/8kpFqdKG1YZtN0XlBWZ7E170CCMMjaLFOunNWiCnFYwNHch+vA+e0nFO
OJEAyFFaipGZpjhI8a0l7ey5CgcX2ReruaeX7nkdijvQJmrl2ZSLh0T8yCgixzfwTv5mQmJY7N0U
dy4PAZo4Q61MQ+n3wH1kDrqVAuI0FDVNIIWi0m/YIu7ykPfmWsf4rKGAtiVvu2eCBEI+xkMFm3Uw
7pgxaCW1RCkPSLYh32zq07k+ZU4ID6bi5wDPR15J1d17pRESRgGEMvVBf+UbB5fC9ybWwt7Edse3
vrxn1UHpgLPdvxR1EHOJVKeYJ3fzA1WIkteinUsfATeqhCpSZJ0Pbjq4ABhG4hGEQMdpuNpbCDNi
++/3AaqeDUt3uVurjxrUO0eiG5Z/83kMmxrDWeoYqMymwEFt/Wt+dstt+teGsboLQ24PKgSagM8g
dHIq8/RrLRFtFWE0L/Q62fZpyFeXJ8gYrvcak4euDc+jXvuCm3TFPKArhGtmmUZKEBkGPYH5V4SC
LtGH0bt+M8tek7aZLN1u4wh1/WniiGu1PMTaxyWlRIYPfz/DPHDuO8PzGRfLDmseO8G1rTlb3ymA
FLxyvS2t/4Tdo1KM1HDlTw5GUZRkVES5VacoWt8BEGXT36hVcagdWjC9VxRh3ONKtrPZ0gkJfwHj
va5/qa10h+2UguF1xNzWSMC/CPoH9qDPGogxcf3jVWKfwP3poDzOkHxo9H4WiKZG7gk10XCmYd19
LYD2vUrez5ik0QwMtFv09HNdBPjCMUJ22KZSWMbExOfKd4/Cwj/I+NgXLyGAMYoxwVXt8PNRHcjZ
vlBerWdBovam/nleAG7EZDbv2ie68SBfNgpuIbOteyqA482IQHpjYHJv3bgVHudWoA5miGkApOWO
aB7NhTXr1XqoRqytUbwF930LHWr4E7ENnbE0aRkI8RP4YDTi4RTKX4EOQCh7WOzK1+/xs+DccetU
gasvv5qAt1LrYl0rr/8vBNGpTd7kX9lsgwXT4rdIHQyWzsxHV3z+jc+GtNLk/pdIjJTSslBG/rsM
/5veJnnnN7V7tCIah5G/dRO2WgsgXKbIvyz2xXxjQcNcgjLays7Fj2irXsLtaJcgaQgJO2ue/Iwv
2tZ9xFxu+xN6/SmO7JivQM6PweGvQFv5NxSdZ0inaIuqrOvgIZmpQ+8waBPpYKSo3OIx1V74CjDG
MQA4N3qUj4/Z0E51epaCmzeSPoV68EDK/euLSS6klbRKra5o4CT3knPZwJhxGQLL9udR8lSPs9/0
/nycUzaxabn1h0OJPFYBtqk1+Mnl4Eom6ksdsqpRA9Bz4XBb85g4aP4rwQPJBoby4vDzF1tWf9Hc
eOSRMaG5AL9cwrVulXKNxF8sRIqrC8021EwiKydZqGWay4SB0BD1E8pqqz052A+mRm1R9Dwg/PIr
bc2jbAWbM0kHvcyB5oybToxxs/a7Vh2lsQh9oOV/42tBSrZY6fdcEz+PwNojoY3EK0BDAgPmDRFQ
/ViSeD2XnJsQpqbMlsY36lWDEDhab6CvTC+sDATyKejgdHPPPIURWYxx0z+NNmqKYX0zLCQ4Ez3S
cKbmy9SUix5jL+2U1xouqk/M7u3NjR6eKfGISVDq940nS43hekwal4r/jFRxNJNxw7t+TuOVV5i/
8cMfhVR/GSH5yOZugwEdXGTKxCkUFzWGAFTyQa4KC044mU15oUwQQW8Wm1R75M2gEAabJ8NGP+Pq
zbMEFU/14+q21MqXHO0+EyItszPsK/DqQSvP7x+0dsqGOyrNieNRRk1FA/bXAs/jTxGRU57FZLk1
ZK4db/hn54rD7ZAq613zgnNV1T/JBG6G+PdSSbzQpd/dZaarq3ywMpJe7KuFgoh/fa+bYoqJvd2Y
t05jStxhKTpThRHWPzPn8LITiOUAsjfLbsfvTaUln/f/5ALC+SCGQAr80/lVEtTJco62/bbLpeDt
5ZcYZ6u6s6xd9wbDzoTfLoK1fi3tzlocuRvlPeAGVQmZ51RIQC9DVz6nShH6wvSrOmkYBAEYay+g
MaU/PiPxIbL1KkTosVz3O2M+L5dI03hPNvrydmyDPHjCFCSHLj09Hf8f4huSTlZUgizwBdFPKpfa
Q7UAovV+o2RcQAR7EJJoM1NFU6bJHJZIq2MAw7HX/jvQ6CeevtokvkpimLJWPUg8vZyF/UYD58jZ
q+F5/dEamL54TOr8+e4zOMo7CVw6GpEyr4Zs7VK9XlwtogHjpLlASxwd6jxGgVKtZwujmeOGyhAP
tC8/IRSHzVcGdSm6GVwQJ5SDdMb/F4OsXohjdUzWcOEzZ+KkVFnjCfHupO+gkiyCyr449H6nXj4m
FmP9cGSMZCb7R/foCck1akEbwiVD05Du8Z69elJR1c7qtvU8Nxy1Y0N7XYrg0ou5AIAK9pzug3bL
ZgzjBxPahg3D+ALJkvLTzA2C30B2zNfuAwNEZCtUpwkl/47JODlVX0aoR57NCaoxvVfPqUwaeCiS
6Z/DTFKhs5CImS3W1ruXhemtTtcd4TnNHAiPmtkFkCkTj8dwScAvGDSfNVFX9ecdItA/dG/ZXxxm
EhRcSrg/H6ZlbeaT65O6Rmj5ooZtKMaO0c7lnJ/mHL7fPASPx1ozVpLBoztdb0etLVsLNeJBDriV
3x8VnvD7PBCrvW8HQJjh9kSsLCeRwBfadKC4ytLSGJ30v5O4K88nZoIF+9lfG+pkwkIc0vUq71WY
t4sa+yOHL/1lcYMzHMSPDOFVVQOtzCPw/uQ7UPCeAKaJOzzCiljQ9xBOQxO1u6BX75JyTcKdAK2B
CYXPRsRi6BywQpFxA1vzfwpENJtH43ChoCcyyhBjWg+hw0AMQGBFpNmtPIgOyIwF5nOV8TT6277T
e+b8ZKsFUxP9++4cvftt3DNyoAwee2qBQsJzz4vNukgAVLu+/qSCziOjx9rx6JJ587M5UFWJdYLL
ZV68+EazhUjw6WhvJLe59uFw4TAjaxPUZ3t6CONEFFLGR7qb4xab1g8IQJ7rnHTT7s+3sr5ySMsg
OarjuwI6A3Eu3jo0mKEL1wpmmPweMtH+eXdOVv+ZAYnZYtHIe6JTQi58t1r+XDjsNeLFB2TNaxig
6wIm7ARWJNDvBcKR4zEdSv/1nifbmo1C6D5qGl69Wu3fpfALvL/1oApPDRsFvbW17jMeeSY2U8m7
8zhq2wRcwk1fs3cdQJI2+zUuRBWsr+KbrUKH2r/9fD1UTcIeapZj0lGESScUP7wPiV4//es92QRC
ws0f6cdsqA6dM2dnPYQI5R6Vfly5mZCu8POTUCMcv4jTG+o/qEN0Uzcvo1DC4kmGCvFC/pJB76G0
CDojSm1Wha8fk+a2varVlWBt4LnLjNkIrYE0Pw344RLmHUOCOYchxHWocEpnsqyIM2Zp+TAB+fs4
6h/yv7CgcwRndCUcUFXs73ztPq4IvhynGNkkpwhjvAFX9DQJq7Co4xSvILJF124H1q5K2CV2L1Kj
xEVUWI3GH3Sej5PzDVouIAWJZJ5heXED0EUhE7xRXjXdS7wVHHV5ITFzb4mknNF4ZulvIaesNG10
1vOr9uBWPECbULXB7RgqSXRmkhFmhFZXBBXyionGr+2FoLyCudIAlFm73/bxNUYZA6vP6VODLFWx
Mr/QXNJeprApsdos7UExhtEi6Korqeba/TvvakGYCtor0Vtln+oWWP1vJszqB+PbGmadCn5Mn23g
iUksdvXmF75uXvryPDCfqStbvHbyVA63g5/OBYercPaipeqwPeqcXjEWmlh9i29MUEZop4DTAD7Q
zClGzN0GFTZYFJzSrbE2zfx/Vexm+3xUYkvE5iHBa7fVHGvFrYxZxj7YkoZbZC/+heQXGY9IZDc0
X21nVfkzZxNrhfh0yToULnDUMXhKq2DWxvLZcjpMqSz71m/4wBJy6MRmgeZY+m9x3hiUUFJsynzj
TsPU0SaBKPEvbHRx/CjtvzAxXoj+crONGC0KMvnl3xMUQQPNQZEdln93mwzcAlzupk51dRT8+PAS
S3RS+dkVPGEAaGikjKBlVUGZ9ikI8Z0pAXU6P9I4oEE6GJFrlj2aDN1kXKA7AVW6YCOJjOhDJI+k
d0YoK+hhy9dPRpMZAkHejK84cOrAdcGilqNRzhodPJQWm0JqziCadjoauhwJpnd4W6C5Hov8Gxbj
nQxoh2tNUg/ZjY7YQIC4OicNLC07bza783CnXo3nuYqcedY0ahJGw1yFJvmf29s86SW7tQiitMZ/
tS3YCYKD2fOjo4CwKW3x78l6TWKz4tXieOB3JWB5cCoxmh0vcypAL003lsBiPVsqQ9s2MSBLt10v
gvZ4V09ht0gimM8S4GILz1q7M0Pf/uEBhqRN9E2xRkoln617pjmlNHg73yZhNkcEWa/4Y9LRDU+0
A5bsAqIZeTGTvo4Jt4IqSPK2i/3h9O9v3u3etCT6jD6m7uA3X1tos3/2SI6vknLIErJk1urTUBYi
rJRabV91oVFk8JjiAzV/CSEbnKG9GlS+gTiLZNcPXz9e+aCllqw8oXKOr+NO1m36EcnBmdPIzH05
qsLK0b1SgYhG4A7ho4MBCxQdMa+Ozlht3SbiHnZHJl3M70lR2jqKyfi6wdtirlRdVucPinQytYua
W8b3aBUlmE4XyQtmuP3EYrL8B7QoHh2u9hRbPjrq/hfLUKYHEWEF1bFV0uk0r9GwAVzVRiCmwlXs
rXKt0j8HPhwYhyOAc85PmZR/T5K5ClPrlj06pmMvirBz0F6g/6axa9N/jJ6whC5BypQ3QKFeArZu
ZZMjYWxKxG0kLDu2p9ofjbfxte/mizSVFRU2V6HABZQOshB09xOG3xKgM5Cd99vWvW3b5MPDXxWa
pkjkKkIFC09iWT1HMlE6LC0iu6nlnOtHw+GYposiUO69S9G6kJdkp+p4yEoQ9zdmSCbn+MrfzG35
t2N/Zv7MnDFtG716Qgp+Ws0t8dCgccYqamgfcS0KpL7gJEHFZw9we/dzNuuIIWZr6b/ydZMWm6u/
stgSM8BCpHpRPKi+9waBDR5Vne95lEDLgYqMozr6Rywttav95SLM/7Je/Kgd5ZgDgdV6WkCiqPim
CFoEohSIuXUwTqmaJnKm5KP2khXrUWTajtUeqQUiaIP8fvp/+7cNvfFZf0biNUmoxn6nmIQmUWIV
WeY/VYkrDXSRjLYHPpxjRGsPStmKO5UdkRXJEor7ExaR+vbLK+EMdsXj3d9dwiFVvq01W7t2UN9f
Rgl9F6P9jwGTy9kXS4HCHhNG0dQga08uCDEyuNPBzVcm0RGJtSvIm8zrleC+DtwFA8olywpLrWuY
ziUZ35CBE8jYoQLOyO6jcDthBres/AFP+GyoAD+cK4lqoztO99N56Qz1FsxwqoxabWE7KTI9t6QQ
3AUpTyCyDHDd9IgZpdtxyIGzpYba3CQk9Ixtd7fSe6b7CCRssobcXRK9VV3mxX7lpo8XUopD5/Hs
+Ue4v3Exk+gXlSUqlc0jsV/6RN4mXQMviWZsl5WJVAVszcC94+mYLx7dmyq3NCYlKvgKQmZ2bln0
VhYsiOz4T4KFGw20SaHMBsXX0GJDxtj6eqs5m0ZRa3AhmVV5wbMXAgLkDrjA8i+CbJ0fCQC7reQ4
TMGXBIXs2PayeRpALx5djpLaIO8dcZmpDQ8O/6uFWmGeu4ea/vB/oYuGnmXHxlv6oBJdSzQwXNOx
aHAv5dDVgQ7F6v6igUI0HgASnQGHCDJTPe/isG/PEGT/U3gdgFYovRxbqMHO71Zh0TCMphO0tSe8
VhwjUjswwAsrJsTbYy/523R6lSESuSldtodOsOq/v6xx9q0LifCeggUpKbGMN3ahhMdBXevvOae/
qE3sHcAi78HQat5Lvo2U9c0iB0/xzObBZhgolZWneiIlWqkNqlYFyD+cdXkb8v3cE9wIen9MS9gh
pAg6mep8mXLZ4nt4GTptR0sxbMH/eNxRtKUm5x8/a1nb+E5SbrN69Hj7Np4ieM6O6bYlyM233MD7
kSh+/Rh1SuiP41vY1Zqot2zHlC7Nf6D98NQI7IIm9BBVU1GgKWvDnz/ycpj5+lJktGeD+P/+Xniw
dz6Rt+rg9V09EHrqfUVA634GNREAwpGhdxiawUsgi/Og4kaOaGVtL2QcEMCdaEcHU/Wp/8wKlqz1
74lIOyFhUPGEukwJCNrZ/0XgRWuN7g1MeEqSFwti0Fp2XeaEigeizmoL8QbTQU0vteimW6DSvynP
oQUbzzAfoCPDY1cdVvKR20eLO/SQ7twKu1nIRartmPi6HMw2pyauUTLJxoXz8CQCv7hAs+tfBO4M
2inoX9cnrUSBC8qxQn6sUqeFjxZp7emcB98fG0/W07TWEMCyyc7zJiBsskkh6g40R2l2p1+4EFrc
5wWZKbSoUASIDjWuhgZpKtbcF+Zj9/vwWY6jPjSEIiGjHEka5lN4L6oAscrr5NPqNX8uKlpv/pvG
E0n3vBX5oKb7c608P4XCpk7IPBT86jrgQIPMzf8W1X0MTvs+lg/SvF5qr8aMKJFtYav1/6lAwGaz
VOkllArhgkitF3wBdqkE1AvNd8/GjUsznrxFOY5K+UeCdplY/c6bO4y4gRUrJA3nWeu467bnTO7P
RSuqzeqxvnhR7DgrCTEfoxehSsztwrUC3lhsq8HcF0gIp+OEm7gv8liq8HHHBT8xZwhR9h5qdVxg
dQ8JnwYfXuE095Lv1w2qgGqSlRcAtQay0/LvfwxfmPo1P6NVJhmwi/4IVXa2aweKF30ngWm5Q3vM
luzvoRVRNTTL8aDsFVhu7b1EHCQ4Hj0EXUI4DVyz4+dha8VnvDmENkDZo+3xzNQQ5Lrt8pT06qdA
pGdJWGcIjMootqPI0vFsyiHt6liCtDO8cSXf0o1RW1nlMwnvJnP/X8X68SRz0dmChTfkdM/HSwBO
IHBJjg25+IMannwT/fIGIqFIps1gApTJZznL4sbUYb70l+KYM4zd4Zc+mAvFAb3YXrefY6JwE3Wk
Sj+yqxvM0mYBjED1fvV5WtFR5NiFOmzKK1tZ8Dfu66tl4/Ap7RSC+pGGFaEunQ6ynd5/SnTo99dh
IiMKFEVy8jkFZv/CnZMdNDctUxpQ5Vx01vbPyPhf4QRdVn+TFN5iiaBeOH5ADMmzxWvBElLdNHcY
WoRAIBTAfbscJLfYUnxCd8cFXLMAgGi8Z7ne+6H6lH/U+vSGbKKHE6NcmRR6/rdV2uDzEO8aXbuV
o8fGTEnHcZ9QP+OMZTlrUHyi2X8jvef9zOx04ByPKcgfdQPDZU7uMWGXLqeWroJh2qSnIAKT9WBK
LgLDchqqgCPE6/V+qdsXrE16UH0EN1Er8MJr2zY5ZhqnfoPA1GM+YoAUQ/QsDT9aXq+0qnx2u10e
iL8BO8P/Dl92ktZ5VKaqABzwlt6FhLAvqCFTn1QhPvpgP8Ikbqt2pqtT+E9YcEcbiupoMmteXOKE
NgQ2FscKzMBmB3xhdmOtVqfI2hXJNlT4QDtbVWkS9YV6uWXI4WDLyl/drQqbO7h2Efmm78W2ljIH
FGxhqcmztk9B8ZQ6Q3TabvMojNSvs1tguDqSiyHXCPdc3aDlM5oho5ID4TRgvmGqQ0NUXJC7Pr+l
6T3bPjfnd5reIErikQk+G3uUwH2WuOHTcBgGSIYauWV73Up5AWhJ/KmQKxIjbWIGMedsDcvZUxSH
qobEQ5hNNKib5uRaUCyWzVvcrSwNWr2D2lEuxXS7NXOo7/iSWqY8ao+bRd8XfOaxlv5rKzynsvHj
TFbnD+kLUUqgG6b+FiD1Acl4px8jmkw7YeiBMri14SNs1CQxneOCZnL8JuRVdwaLIuWEV+KMgEgO
uVubj1L2qLuc5flHouPnnpO10O7phHMswX4Xip8txi5OXyT8aZ4h5T8r9t82kXSdchaRmv0OGvob
JJqeu6DNXGzeetVKSPZPReUlcICXBTo4Zs+m8WsAxvBowUHHS3fNTIMtB6yTnftWdeGQAy/9GFSB
fqFLP4zrDM94FbecY/rcKhxcTDpUkC+EtMtf+UVJTYzhdMIjUPq2j18+wscpPK2EOg5jBfIrn9hX
Q9cAPh2OS1E9dDsuFxKq8Nq4KaNF/84NMJoPYg3ONYs33kUTTGDB1tC3+NmVzCy5r6Qbjt7EwE1C
Bic+UQ1vuYPt7ZDAQh0FiTo3Wir7DvUZY+9QQMWAdVPW8nMCs1DZw+4xGLRpZspF2SBMIMUG/0x0
0wf/6y1uh1vi7eslnsiYMBdDiWR371zQ9rAeIUdCyxu7lhAP7ZO1+XWInoOCL6NcAsuguUOsQBqP
uchSpXaQUyOGkf20VK5TuDsH+VtxTLZJYt7AFVzJwEQQdfL/E0RAN2ajyCTAdKUyLF9eKvwrb5OP
qel9UfWOaEb8Ow7XxvHz1Z6ONZE0y7EZpiBJnIs0c4jjIcUKpEkUoA0IwEJvTl4Dn/QXkDQRJgSS
uBUYO/BPh63CTMT4063SnLw59vx+fwHcL7wlrZUoQX6FSMg3kfIq0u6ZD4ExY3n6yYEZ5AVSL0oR
Y1tO+cTriSBT/Wg0i/4tvKpiPZ3zKP/GmykuWFgYYM8msXJb5BZu+cMWW1g2hgdPG2hES5lhTM+e
2D8m0+GRzCaR9EnM26N22sOHDEOat14VONrD6qBxMEIgahtXKxJna4qV5Bwx2Hj/TMmKMtBGt46B
9ycV4m6rcOn26wLQ9DlOZAwaoN+H7ToJVjXm63OVs/zegnQGH9TF+a6fQv9dKyiNVngMm9ton181
DefnUL34GfKK8BI+AfiBCr45sBJRn4h8vtXc1gG6QXylIxwoxJQkp9Lm8ADJZGbiDw/i+aDTGmFp
g3ThW7PKMA2itcZwZAq+GuvpaxW4PEg5fZKO4BIB+JwVMVi4JGjMUYxjggHnp6otPxQytLvKmZgQ
EDIiuP5Z/m/bMRjwW+KPewRKz6Ongs+W07YDaacU0HGNm4kPazA5PXnaFIwyhzdNUdsiCQyaAMqe
n2TrN7crH7TmCjo+nNTdGalWGCN7Ih7lW4JadYHttRyffr+yIHERMbZyTkxk3GN/E9BQb771B0yY
fnRBMN/9YScK159UkQee1FYVNDvJS6paz9lmX8tHeSjTg+J0/bJpQTa+EsHN6L2DY22EiB51p3Ws
dL+jPcPGc8/R3G0vSQHoclqpBaov+uJvla/AXtLGL5ZtRuqEe84xW5fQqWUYG09vvA3dBfy7St6Q
q7eI6zhnBK/jdKpzdQr57Kh7lcLSLpNTcOIYMflP/Qut3tp7+TLVNRrCS2c8ekgSYbSzBw3oe1yg
tFD7vjQkJZSjVFayyayiXdkUwvDnWi4IpsX8D2NLzbuZApg5k9ciMf7gLnxLzUBgzEMsvHP4b3K8
//2XbSLv7gBgi0O4od3NwI8U0IY1mg1JQR9BC0+jSrNcwuowRo1IHRrfid4ay69YYXFX2cQdcTeD
ImYI9yCeIkj1EVvvFwekOM6hs2OQJNu4NUfoNfHgeQ3lztGRYPe8P+/nOKFMM482vlcKpE1vH1uk
xpdHKBKJ86I/UGguUn7IXbHpSaU9jba21qnVkdrUjcJtDP6WN6sxrSNKpjX/MDbJEZJGSax6oJNG
sQXrYsHCa8KM4VGdZKez+CfBQ0kPBbfwD3huXWNJMQdHm7qZ17Yqikj8Cie4pzoEqMtJSLpdDos3
rhzkwohdpBo+0wEKITvZHKlH8VDZEbjNiG6cifOHPQavI1df4Ydxh6kbFUvmbI7c28SfvNjCpaB5
hqMZg2XJEh89FYiSw3YeaY1Qg7HZOVaOVJx4dgsOvUWpefV6DaIlccSu9ST31h+gff4oojT7pn7a
ucvrwkmXlnteSrbdJasxGqktuXjl2FqdVHo6PZjvvK4h3mtIhDOQxPPYjNWxW4+xD0ijq0VQmu7D
Lufv2dSBtqwWistL/7H4ZjYBfRku+wnyeO1uc0FUSmqPaB4CRy55b4oIwL+JFPwthkluS/BpIH+6
UUdZvxJHS+HTavsRuivuDVdyoS0eG4Osek+CiT40t3KToWZQB43HfeTCH3hufuBkqJZYUnCjROox
KCSJv6VAtWbmGFkyKwkuUs6EsZjlxNY+l7hwIYN+nMDvRxu+93xYHW391nFmjzF7r3J+ZH+YAsY6
bLtto7sPv3T0EY5Pv5ER7cNF+EdMyIv6QkuzAfSZoqzOfYip+UOyD40v8kH2fA/7S7rYoXhhy3rA
t3bS1iauqT0sc8Ur6lsfuw5IlDdHXJqMq0o3ftZWG8cbj3XFJuhC9akh+ZY/SV7lxq02Nebr8BSX
GhR7pK5ntC0oLdRaD7AXDZMkmpw/nct+iEzPdJ1kkVBXrEDNjVFbsU9Hjbn3pDd1O8cKrAQI6kAJ
Gtoih5Dade9SWPP+fat1ZhAvQVSkTbx5Lum5isjsUKEW4h/am8xP2m1cqLVOUVPROssUPgIRkfPV
78wrYESVz0T6oRKKCO2FOMVmCYRzBSA/lcojhRfBnRDqQb/wDmpSavhbD55L0z+UF0eJEr+x1bG7
oS+y0LlcIbWp7HauYoVO/N7bDpAwTFb/xuHA0OqfMJQb1y6W7u2NX3CKgbYXizVyqSFvvFJmBEbk
whiTehg24H+Mb37xEv4bFTO74mU7676EM0tJxqYxKhsenSm+RXQx9fdV3xbfGL3zkgOkyqFLb7j2
Wfa4btFr4XirIOn5daeDcMdloUBvHBZdPXYWbmIiuW6nzvym/Gzn/hmTX5oPcr+a3W+HdwdnZOdZ
DN3b3ilH96PQfhBMhtHEfIo2/gTHIFD9leG6T5RHD9vX2MnTzHCJFXYYV04Fkliz7LNuh+a1QkTa
kr1F/rnDX0JDN5FAI+j6F4siyJ8V811+FYdM0QAAkolERJGlAl8h5pc5MoORegNNT8f9/Mc3iFn8
C00P8sOl2iCTVFfz1ivkp+Q2ff9xv008uEnvRJkaVnic4yrJgNl1PBUTty849/wuEP1YGaHvO3mg
1HZOmydcWRw27Wcg9U2khlbn/DRKsdxZJSx4d9NN3Yj1cwASXR1xUUeGBBw55LHRe9o56KCKmCBb
H1pkPOB6U5Or5KggalMNDr5dSW98xQmrXA4oFQoKULdVluf1ReVBxSTpz03sBGwMA4wQN5pjmcY2
Aqb1g0GRN0pgiVIT7N2muUstZ9usNPVHWRx/C7Vu9PcxY31lWtOstVK/3U91ePon7kqd6+GlRbCC
4SvpcfLyLOoEsCjgL2EOTby8hcJYZAosjIsYf/WRMJZ3aJ5QSmDT3WkwxOfXIT6h8PA/W8KePi2g
fIoCZV5sviZOd3d1Bee8tBn0mcxp0a/WvYLM2pfO2WJE2gtEoRz1m6l33Qgns5mcYaq8B6SuYalt
kWRrsdwBeihI+2CcYu/Y7xLZVADl4c1ZDHsUMY6svskE6P+zLsF6s55JLQ3Dmcf1bI5lgSJ5P9yj
Sgq17ltjHbAvjJ+EMX55CKOE7jQY1DWy2SNVXi8+pyPtN8FxmzODzpRvMU29q9W8RbnAjTU/Qcdr
zclbx+zw2FLZT4udk+hDgUEhsgm0kCutazU0IcLizkJ/ScRKzVGhnG348CX2dYSjxn2xe/V3bOFD
xccr/4qFk0BFUmD1Jdaixy+ksO98xMt9ak/b36rnQiikzLIEzH+hQmvaE6Fh0GOUb8fx0qKols/w
WSVYseP0AXKtgZCXlyvr8puImWs3OcBCYoR1jtPGO0U8+rjeBictyniz6d036GAXQlckQNwkjeNA
5FlXtusiCP9o20CuDtpjkeYoyRoEV+H6yE97CIE9NzShc0ApM3eOUFWKngHDlNGw90q1ILcW01zn
WaYy6saie7CaIJVdBcTZXawzvY+6EIdAo1/6AiqfHcSaOow4IO76jk4QMp9iUo9B72Y7BOEJzVov
ZIypm0jrEgkrpyrQtwdo3q/qMJ/Ka6L9YWgQ7/NTItFhYHqI6BsVeFYvG4ZKS8d2MyjF1UH/p4T3
h9JyN/GWzPX/vwPUpEMf1s3C0G7i/HM9uOjXX0XBFX9CiLKpoyGejaxwKROoa9D4FIAbyimzoTv1
PXSXY5wJ1ypNzP98nKU7RK99W3wADBllIruq9XeVUm7s2WP8vOkfFnVU9ILoMrzNXMFkJ9SqX95y
t+ZQiQDEuwFcokYMi+htNosDsh1xpnWbvJJ1IfE2Sg2BYZ9yZIaqzM8Rqy1i8SU9ZuCXtKRSakZ+
ylX2q3lQ2ppxOO0OKr2A4sesBSgP++jaYmGGOtbd91Eu5+4Ldt+SAVrW+Q+h4Z7fJB4bGk81/rdL
P0LqXZxctUpJTyMFgzbXcZNR6Nup4dCd7ueHCBa+5QNfwY3T/92k9iNqLnc/3fAMVyFH5VOPTbUH
QY+XBRnanhGyK9IEvzS+pXbmLFdJ4afBMCzkADj12CeszJ5Crur94Pw7ZURSgRprZeb5NEeXq2mD
ofSvwjbDEcwhIkmacpNJp5giQr0fuwxSb5EHIdZ/6AYopVuudFTkQAN0UZ+nepX0ZL8SCumAeURf
NmR2mzYzN+YytwlIsNltALPeV3Eh7XrFJk4M38hZtQqSUxWdaRoNsM0/PpZs2dQdW8rVnEibsxIO
rLIogOdRXB0R1jmmujpaEGPh2HbfDWNZT4OTmdJM3kz1JZGlQBZz4Gqx6pW08EtMDVE3NHU89nbc
mj/YDhUekdM8GC3KOoAbK/xMmEj+aGQe1ZbZ34fql9FiB/aN30ceqDlGXVB8gTv2lFG1uYO+oV85
4Abo/ZtupTwN2ariooQCAvweOrchX69UOfrLlBrHsoxIBSe0Zxw8ovOgpzAZ/wbHgzzsrF8JhTgx
kP95nJiTzF6OJTDlEqg1da5DsOz5qKWHuxrAjm0Wq87nGzoki8ynujRmqQg5EYleA/rfVHhD4fOK
CXjCT1EHg1Ys4sjIeK8Z/kFxZ00VqkZvucUviEPKHXP3PZOyON6W8iYke60RyIC6yjDafAWHJ+qa
vNfUfjuJWwUE6ujGOivL/Sa8CxXPNrUKEuYK+C1PHt0UU9bK7o+5YT8U/n0thbls109w6fc8Fp0T
PO6PfScm3x+HWvqfa+JsZ29eNrMEf1kNhe0/k6+VMykfzyCm3ANxwKlz6viC5Av8rbQy5UK9dlMN
/EiSCzV4t5jUY8TE6qabQx8/2s/6eHzBbwrtQQ37WJZBvG18OyiMjI2XA+w+H1/FLVNoUKTi0vvU
HKoa7QUW6iyLbhuGn3bg4zOoM0GXaTd274omGr1GUmF3qV3s76liiiR2ck+LgsIEjzpOPxWiCouw
qO5XWbyrBWtlN6g1JkJeUMUsQyoxZBFmJyspgNWelZYVxyfJtPFHf/kP15MdQ5eH0pyfzSYKMEUN
4Vf2/2nTWEV1DSWxIbXv8R1J/+YZisg6HYyDCPA3cEysfVbU8KkBKyI3rBlohScWCZ6weyIV/wqi
OBjIYJItZrJuruBO+RNDAz+2B17QJ1unIHDYQrhVtVJYy57YnSwwTnzOJmUL80rElNqwnCW5PrWg
c9q1sq7w7qNjt9jfCncM+CUjI4f6xgKcdj2MShHZYfq3voN1L4q/5zYX3XjOd2e3Wfe7uYBoXDh0
TL84x1ov2S0D5W0/lz8fKsgrcr8VWIqjPfBID3RZuqdt/ZFDLjAlfDuxL7lS7uq9ach7af2qWLl+
lw+S1has5p8vN9QhSQxj5Gz65z+4OvnNqbJg6jH791ZcaAsdxLHsmiLkSLLSRzjyOec3oYS8NUla
GvpNWFHOS91nxEQeKptMXAEpkU+kJr4dqjLaUxugpnlhXN4Ia8lJ2WfLDGVBVhBEadJF1Jds46ue
wlnDX9U5WgTYHq8nA0JPW+ik04ZtnVtHtz7FUvGoSQeIh+z0zGlwgu1xfzXJoThB4XWMVJSRmmoh
G2dBI3d+D0VW5djV26Lg09rMDBUvfHllBwg3X0lkGK07Py0V4P/DdPx1QdQgNz2NquZDZVQTLYHJ
5QJaFX5fuDk1cWsBy+/yKJLhT/oTb2i38wkJUuYgwCBxkIctYq7bLTsPvefsL2Qawa2m/snIMmZ0
TC1o3ijUfDEWYSqu+ozEPGfGN/Gbh4bw0AIHc4c5wfbWnG22MZ0eB4CRjsGVhBqVM6w+vrjmVosR
VU+aU56jR1g5hCSDYG6mZwLiHSonWEiMFJz1ftc/RrBYK/Bdin0uj71fECimS6sICBc56+e19TXb
ibNT0wsD1auAXZL0b0MQWLVSUW73FqTnSTYlBFAkYAPd7ftjv7aV6/OR+sGQO4bYf4O4tHojAkD2
+49B9uwidpGTtsSAioklL7YGrzl2viUlEztKXenXYbztCe9lbYvgrHbKOl/xycB5lC6Bj59mDb0K
cacn/dL7oohiYBTUWi1dRtaFwo4NjW4weGQJX6V3Txw8oN6pzavA0uy+Ko0fHu4KciQqk6dcng0e
/ahutlvaqT/MJnMZ3trx8isUahMsjMYxeeYo4/Yz16g3SRTBprc6Fr+IXdM6WVyimSn6pYZFXjXI
MIg2AlJTcsIy5kIh3F+J6b5SNEhE/r1ZScKDvgHx3lAKHIT+8wROmuDidVrOh0GbznZLH6Dj3AM1
Nk7cZc4EHvawjb4s0zKajnM3ZI/Txs+hnIMP5qgmHstUc3wk+jsQ4Htv37n5Z4d9a1mnHh/P0LXW
0M4Pk/onKnfoVTIA5UwPkwgQKgGTAP1CgIHmewo8JAzx9LloWVczWlJOADXR2ogYGiXpJMIhJahc
Ui2kLYQ0NsyOOOdCP490I4TAuwKlkJoKtEKuaDZckKCz3/9sAYBodECv97XocSSh55YChp1oRvnp
0hFmYzEmwrxHwM07pwlAJCrsfUfth9HsF0UwPUrP5Pr9cpMEmZXuouLZScv6AywgbMQr9OFC33TE
LFb87zy9nxsgGNWg8j433t5pNNhgkLjHMABA9/VTemIwA8Vds4b5m3uBWvKmgfsTmfX0qtck4d3Q
bdMg5tzew2jgVO2fyAoNflk43ikHnGFjf9SU55aF5hp/A2LPEOLUffJuDz+WiXAMOx38IFeWl5wU
VXcN/y5RXPMosEm7quv421KvThCz0jkIm4UyAqbywlD5K7j44PcBGNtb/nw1w81U7Zievb8JeYir
7gj3OdDTmNsq/VcCCM2Ge2yeroyYqyCH27Jyrv0bHtthi4Z5KWBfe7DUoCi56Xm8fCl2BIHPl5Oe
QoHGQuC7GVNoeo51390/qhV7BpAb2dE1jlLjZ+69BmlRMg0qYihkP/MApLbFqi8ja1Rq1S8RHdtG
ZHX26WFyql0SVTF6T2/b4FaLHnw1/aZp0M6XJaMhlrsIlXqJExs40HOWgNMMtzNWarkM9PXhtq21
Tttsf2r1ajgTTFvC0kkRqI65M2p9Lx7GyCPwkf4bAGILufz7iXZ0aVj2LhKkyMlGjMMTSrEteUqf
dfgfLzZy81qvw6eo/zi6gcGshZa4vD5XKYEzNJ3L0h/DqSex4DyXYmEF9CF3c2MkyKHMBr8q4tzu
h5gR/ZGK9RFukUJ8zSljf7T9enZJKcct+cZ6KsOvjWsxnmY15YaINmIxPW7FYn01N7FLwLAEDD0y
ECZwpwL0W6yLHB26uniOHchMSdy3bo3jrVSPMvW8yxnniNaYcafdRiLq6J/0mIpruMc6ykPTM1UE
HiShbOEH8GkboxVaLJ8BacGyU6Dg7vxn/BxlQuLHlO8tQk4hmeMI+Ay4QiIhH8FksnGVLt31Y9bV
yA1+aB+IYk++l2XJ9SZHPWq8h9lmYX2QqTbwNp+Zu6pJ3chVTykm928wJjzFDPSWc8NrHv84U4NK
ZaefD7q7rtoJ2oE6XCLpmdmySu5KALFaLUVNkPk2NgS3sjU3sGCzbFKQts3K0gqemxrkbh1JoPYZ
B++k7v7IQ8urifnsFgcL+MTd/v+KoY4XypyeehISJdYyp5qDNOaJLp9ZtZ7kFTYGvtoKe+yDUx3f
TDExisptBp3K7HXO0HXOax5dawCK8nByPuqpG8jm6JZawRTUVmsGY2ga4kl6xyyhrONBheu/g/Sp
cARCFzJFqS+xXGI/izZeRV2euwxvzJp6PqFXqgutU5fY7EV2YJObo9slse1b0uZ8ew+7Mi1IHKl0
gk9pP5sPAXPRnCAe3uLcwg+EURykQz7+U1JIHmFezV6bszte8MLgGyWXgzv+RDWgK7McKpwHz/Zp
4pQYwp0FwtESC2zCr82PXca2lx2uLU1qCNfKpEZmA/xGwQrhbJHivKNJTuiSd9c5AU9z55ybaOn5
HoXZTPtSaeQC8aNzW72ZXpK1CYdpgokRrXBGNwXE9fj0SwArzqc2apnxmD4q+hqFnLJflUHxbZTv
4i+/dQrM+KWFlpovgTA4G5BOMlJmkA5touz8F2KujqwEH3knpbwTzOR0HVdSWLPk4ngd84t05IiD
TIa0LR0rC3m2R37wHlnhRUHoBjTGHRN/L6Ai9qLLj30TtSLUn2J5uKyy7TrRBRO32dp+23Frv2j6
RlZ2FYPgrJ1aX8bbIguHhqiDoR0A7WuhcrY0YSt35DXWxnLpoCHjekF6hlcbGYiQTNg5YoLvTA0L
i9asKoFHQrLvp4DneezDrO9RZmXl2M7DZJObPpd+cHjjZPjZmSKJlhBwIkyUCiuYEI54onvbAwl/
F9AauYZfTYyZFPjla6surjUAOBridnWzqDK0VBdgjv5fajjuu1hvEciJYNdMdA5EwfLizQC2BY/x
P9kpIRmrLeQdRqE7jR7dmtHyuic+6rBbXKYihYv0WmtFbK9/iwCI1IA0peGKRktUjv52g2h4txVO
w1HRbcRpFhIqUlkXvTaVAmAnMWm4xscjCB07g/vNk4N6F5Bwn2SKM3dkpavXw7SyI/RUfj8900v+
dxtmvJyOASfbosuRIZ8/OATZQiyKg+LxOlb13gOUcqKsZG1HZM+JwJvbJpNusL1aHl48Mtws/AhR
i31T/xI3P3EQU95LOpgYgR8Zkj/9fd+8bXnyjGIMRb7DhRllcPXHgQztZR35gXPXWy7yQPwja+Ed
f4NNbDQEmzm2yGUWmRoFf9mPfIJmlPKr3M2gQ71Ivc3bbeQ9eizO6XBDf2p0gs7Y0FsThYO2F56A
IZavqWclb335qL8ezJQWqb99UEOVEvidynxJHaCppZueETXugzJY67L97dGxQCqcepasu0pxWLv7
i/tlBzNYhJbPcHRhKbXHWgvdGtpKqtB4OcqVmOnPZjb44SQo5ZnZi34NFkpn7Xf7vNFg7I45ewhj
gU1jzu5Q9k2xS4+xjmqdxw/CKOV7j+LIWAXcudKQqNLTSiHBIFvuIxNz2UBFQMCrCPw9zABxUWyA
i3jaLXJDrXZRvToo5vibw+poAWNnaUm+NrzmzIk0T0OJDU+KZD/81GmXYqEN5wSJ9Vqm8Arv3TfX
D4zibhO3xJV7FNNkP5X4QwVsR9YwOpsiOIuLOi5PCy0lkC4ix5pDRaz6T6vJW5Q8ybWbtnCR70sk
Pp+jNhy3QTaQkzPcYbqH6Jkr+4PHCaIHMyGuBoN2UlU6OaJVSvfEAOQqj/gVpkHILvI5+OvG1Htp
UY17SZvT+N9cNgbkS6aDS6mnvVR0fdMqnFh7XAHx7GKzs13pG07NBj5lM27O6BtiH1QdBhLHbxdS
cSJvUxDtwPzHX50qxQ/q1Xkozi7NXADmAlxt1IV/FD0JhJwDL2nuDeg3uvAsQI2ex02C2iv+Qli1
dNAcJq0hYLm6fbarbhDEFVdccE5QsDTkr09YG6IaQTniBd71dRcOh8tU/3r66j/9tc8BAQ9nRJwy
fzQAFGYiedylF2DfHUsB9YKDLZIFbi1SbuDGCm1m0GLlNgDO2DM1vKl5LJbFQyojPADDM8uOzLY1
Bx0o2H00kfQhmuy6v7Iknh0eKgLO5Yfhw+MFr6LGKhQGNwpV8E0k9pz1qcRMQyh/oOB4b+X9XMjM
HSfm4zF8aCKkG5h5bhFIrNSlkfX0GlQhcnFR+Yo9o1GQYQ/zoVT/wZNOwxxbM5xWlzC52jY7NeP5
I52kAIlQ32GowFWKlZWK9mFYOeKytP4VDfPt6CEUia/th/JvTaw+MG3aw6E621lOLCXJOyiKiePP
9twdob4sECqLvgvCREHP9BDtm3bvjQHypsgr/GAo/iJm18IUyLMPeTtC9mNBEZFZPpKhHWxwXcNh
mKrKFUefxvixRTdOsMcD0HdI0VWdoujKi3P+a3pZf1ubcI0bHJqaUc4D2wRhU0yGx8i6RIxreDzb
KIJkiwY23e/tL9Q6SB0Fy4ekg7YG8bFGUWPXWLpRecFay5z9mRQwYd0TrUsohZPC1xn6zuHpgEfy
oOxT6NYa42Lfsa/pw8p776PAjUT3KQiqeuxKDYfcbB1N2WtiNeLEPqx0B9oTFsi/2q634jKIAKlm
2esvidRhoJ9PBJ64sXRndsj1z30oLt6XvULdfhojQKoVme8IB8auxOjH1KPjIOp8BQranhgMzKm+
H13Z3n9J9ICrGItqSur2kVbP2bJGQ1qSlRmAxbK1znobcRxp1E/mDGadRwVAoPrVeZUsdL4MWlaC
QlT74yIiHmsxouFDwK0hxYaQys/Pu78Syk2URPevsTyhSAIzz57BjnIzgBGdZTkP8+tifud3UjEZ
l+mzqZfk/p/IozlUB6HC4r93WETU/uhDVECw3yu/FdU5Xxd5JsRfVlBl6pTcGkhKhM9Gomzfg8+k
sGvl1xfEHqA/5reBV9PoP2NalrTXKF5ypjOxG/VRsAxbm4z0u3i8Zis/Zx4lCF6+9KJS6y2T92cj
Y5vJRXncc3hIrCxCj1BEKhpXml+UpQfL1lMsQip4GB3S5DyC/IXj9B5jPCo9sGNuYSN6Rl6IBLEz
F7cl7oNMQtM9v3t05u4oN1UHdpfDq0FSzp+m+Pn1PsFH1cyUMKlE75+hbQT8B0JBerC1ndHfrG8W
ql8WzaKJ3njf4ICw3N2x+JWAntpOad+3e6FmW10uck0YbJh+SWt7yXU5pXGkDje/3FNAYn/a5rEQ
d0do9+5hSxr2G/JMKnoY6DHbdMQehMulKtJ9BpTLNhCjbriVYAleLpLa1NZhI9lKIflWSl3TB08E
EiuYGKMBsGhpt1W2uKflncDVTAOBxzRdbRP4PIkLN67kGze1FmpcIevnB1CLnEEVt/IY8Q0dj2cY
p+l3Gs0wMnmrYNesmbrCYt8SFteKdMiw+8Y+BJVtGBGtCWVhkLqs2Ey7xnV9mJusfCJbbKSgx4hW
Eaz+G88DFpTdyKHfHjyLnW9+xUWlRIwDo4FBTcv6DB75VmyPTZbSQ2mjQoK82KKyY09wjh5SPxC7
ccXR377Q2EtZkBidOq3VI2J3r5+UgHZ/r5SPD30QYtQfp0vYKRNz5QIwdYf+9hVnMi6VUa44jZpq
A+KNWPzakDvADo6F1mdJrBx9kbOUS6IGgo6NUI+yWy8hLYkJfFSbHL2Ou4mvhBa48k4MitHDv4Hp
eDPh7CoP5qF4MKo0/8Kdpr/L+gDu/VsTcZ0zvMY3EN79mKXrspx3vVFbzoQtqt4BQrLrxBljL/PI
WXP5ucqb+1MDt4Fn6lEjwwXDOi0MjuqkUCKDQxG4bzJodZeNlVxiVTFzmSs6kfBsaq00cUin70CS
aI8gAh4nFGJCoKYrxJngAkKnvah0paeLvH/vs4lzXHN2S54bEoEHvdzQaNuU2VF1oNLbjv92zPWg
SYuSrcOQnU+oyvqGcIRejBffEfMg2K0C15gUQS6oJN6yGeEVpkuovjeu5IWMwARJwkYpasi95sRf
zBecqEqk1PGvxSyggNZ8Rk1ebcCfa/N2TlDj3rcypRIlLcpBFqC6BRK4VPLiwjHC7qFVdeCDkErr
iR+hAbP94IoojR9Lnh/7gYxmvZLkav0SBbYTmNbJyhiuRtzPO1GJ2u/tiKk/wNPU391YvK4nbutn
MsQBzftOdhGl9HVOA/2ZwHJU6vupj8LpsBe06uBhGlwwoc3ujBh03uBswM/mQGzD2PPqOditicQy
0cEFd/M10ZKrpdTvLRXHdFyNl7YPgB6wgfBmbONxf2UvnM904rb1f9k5cEpd4q4dRPca3kr0btdi
GhfNnAF8qYBtmS+ETAsISbyK9shoG5cmNtIYS1slT5fG/al1bZbQ4AoU55sN0d57Qa9ljYjn6kjN
xtW3EqhBGUNUSaIg4Ave7WxvWdLqrqp7HquctZe/geJIYQg/R4BvQ+zhCduwcQysdDrtjkGWmq2o
QrSD+OirefWKwKNinYkMkH69q0gwl3OPXauPoOpN2NBLoD21+HXpdtzwlil+tRNiIo507WgAWIxN
pLX93ZSlY4h9Hj1M31ii4AtLR+cCfanNbA7G1+ixcb8e9JLkhcht01Z31ziOLmDPHodqK3QwpgT7
O4h71gN8jjdJ9IuI4vX9i/j15nYbszeWbcXBhGijfAysqm7sw8gnP9mL/8ou23zHBe0dXQiFEjNE
mBnBsNt2cEovqHmm+YCn0s7neyLAk5ksAG71oo1JKxQGnR8HnzsvguzKGEBSejZYGXeZztvmV1Tf
iXcxFJ7F10S6DJuw8GWEJfEniHMBVJ1LlqN9bvw+9AfWKWky04N0RbWdDyvAJ8zEhMeSkYC3IC0G
Cw/cjfnG/sjnY7uEiQwdvP2hz72ux0glS4IRTEk9eIUXiIeuMthstF+POTsDoMzt0k1a7S8dTmQR
8WRnB7voE53FqqLSmk7dsltp3MH+PoV8+8zuOWPBO33CQqec/7IrcVHqzdaf3tCGAVzBuls/PrPC
TNUqtIaKVzZnJ8BPxJ6rrNeFGZ3+uZLeUGKgGCmFZg58W84AlE5sX3U27MF970ky95hBiJpAnP4y
5YNWZYzY5Pyn7ndwTyq4XnfwwNsX9pxpQy/7bmHgS8E79B8fW3+EeCoesLbJ5tT4F2n+dj8ttN2p
0yKmJWrR/UaO3ROMfcfUvF604uCW2ngc1pV1cw9XrJN8DHvkXIacWiG04vWLbuPld8Mc+R4XAzTJ
V6ZlpDnrrIYyOPqvT908kZ+njN1aKytZmti30m6kgUUdRUigCUd0MpnFiWW3hHxbKK1PP7GUXIoz
Ttp/+oT1laOuMFrltIwLLme3YWYTddH7Mt+uxAg5JxUr9w+kBWdUOzTja4JGumiIpjAabJgVB2Hs
lFHMgmZ8s9rT7BTfHGvLJ+sp1M3lcb6V1Wcm9t4ZHytWljmknzu6OYyKMec9MwsK2uS1Zl9Gitzd
tTgMoS8gvJ58I7RQEzDf2J+MB4M/ep8H7QuAWuF3M625UdO69OunodcjsjI/jnu5DD+XRMxrPc+j
qeh0EGPrqt/4fn4jtCSXOj6QCdluPob8VKxUa88TG+TrtPO0KbBznEeRITNVM0+Wdq+Wqlo7PwzQ
jyXB2eNWKAeN9Ap5GrhDeQwSz6bIQTPFz4FEKXcyrngy8+arfNZp5ICzj175NtzKp0GwyzvdMLn5
OJxgKY8YmRFKngBhPYuDVCv6DPQF4nyumgzQxbv2y65ZBPZUQJbkFJmBhTK3f+qqprH1J0ImKEiQ
KdO21//IobTD6WIJazTwf29bOqQPcAUt63+AdtqYINiFLPhJCFVi92+nB86ltSqTJbDa7zX+OScj
xPDNx70s7tPk6uMPeC+/4Lw8ew9d/4+n1BGMy+k/fLSfdPv4raVW2EgCMKzn1XJXDIaJkc9RzH2P
0c01e2citMc680a6kwhRjmEuvq6281YWFGgcbfU4U2K4BPZG/CMWzJr5afFlpD25vkKY+aSFbMJ+
7upEgEA9zijkOYM6Sq/TdaIjH8qEDnYtBUWRaWtuHPHx5GviPy4KWE34Fd+OsnjA0VoD3RsHdIhf
X2R0yTPX3wQ4IL7ZytsOQgjsZ2mbWcM5Uh2ABc3orVgRNXjIgg6F9lElCSxDk9cTxO4oFafAIpS6
2Lx4itZ3v8kTqTlmlOpSJVhP5vavTDKUYoyn44Fd7M89NfWAwCW40J2GYrsQwbyWoq2Gf3WvQhAE
WjXrfzr9BZOlkbnSS22KrurRHAkfguDI1V5zTCLB0NPDCa8NXqqL4w2ykUK1Q1uuSqHOwiOwGJWx
03MhawQdUCgH683QCdNEH8Y1jdR/Kccvuc3xznLNVoN1YmmahatgPCIlcOvF+0m51KLqT4W8YHrM
kbs4MYIuVKEJbvjD3mcQkk3hpNeQ8sKX8rEdkgK6X3n92sFvnxD1+7r763BSESSJQZE5vo18mkvr
fSeH7QqrlLuC9uPX5p3WUpkgJHP5L8LaMu0W0vSUkRnh9EmbMXATEGAEQqbEFCHztl9d5q41q36Y
tXwiRC/5gR5wmJQ50+mKX7vO381i4+alGKwUjrGK2RJ67XoWqgMpM87A8azu8ZBssYafA0qGH5bi
8hBwagRIR314VBNpWXE6Up9E/gL5YEyF4/3eA7iI0tOBjNuQa79wXTwA9V2Vos0Jh9XSo83pi19i
fUPCBDShLmSfwiedPuTnt4CRdw5y9X3Kceu1rPCjWd8h1g8nC+++uUOZrXLUvGJCi6BZW5QaGi+P
l86euEtl3NWI7N6wkx9smB5lidHTGDsAC3FXZ0E90x/vzimPtJGrVoyTi8imxj99jBFqIa7JEYYd
8sgFetc+hnEvG+kOYtlQO35cRm7+eSshLbiIjnht+xntNAub63w4HEL6JA3OoEnql2CZzc0CaabN
HVwO/+qeXvS632uZPmprur88U66qJj6sd5Z1gjZfBjb1Mh+MlGAhOjwch8v+p8CVSUPoIi9apGKP
Tam0z0nDI0ssRuZ3v3OPH4SoPlz1NCn4C2+Q6QT/hYlwCgoD4aTnV4blzM/nRKQTIl/fDO4ePNYy
7tmDCATFOxdCVZ+ubGKxVehyqvVWSwMsfchg4MPn4K7kzfZAgp0en55/nk42Ie4uiuaNxMULzfYn
OyJXytVqG2BoHUTjEkaT9sr6bIfcrfs/q+2Vm/oWzI3VRwUxxoFYsSN59hcZwwdQF37kTwLRkwjV
Js00iMZfablGNXu/5ChuKCiuKQ7gqREOrwuIFNpKqt3HCS8jm/Bib6b3zczZZD3tYHS9ZHJ8pLVt
SU7C4yYi89hgW9s06Y87c+i82wIOQTZAllbJsyZaot5pqe6CKdKRknFl9szWPrvqM0JPH9iVjBcg
+lPtpJsGjvnXPxbh0vTZ8KBCrJBGBB86rwC4c7o2nw6CsO8B67sWSC/5y1i+XAKhgB+y4Ih5GG8U
9tSFEAOZSKEPklRj0+Wz4HF+s7IaK3TdFiyQNe9hSEZHByIXr8fGQ0PkVU4iv7PvsfEfhlHy7kCB
VCNvXL5DADBPeOwIUBeb162C+CRHDUqKfqbQrJ6Qs95HN97X/eWbkpRIGycTYqGjiXwjkrJwqAYT
ut9lkmEDQCZ7XTSkEIpoUJ8wJJrptuAPNZFLksJoPUvCgvHq3kROcVMT3Fs2+j3Bfxbi0gIOf6N/
tfHM5de2r+HtjmDPtAqkISrKztQuHIa26g/eFqH/6aOpADJHYVTQtRBu9v/bQ0f9IOP0V492EA0I
4CQ8r8FECBNI39sA8PibLi8UuNg8QeYvPesGAjyY2jA3QMKa7Lhc1wSP/s36uGRXFRQI8qe3nBa5
KBYZMlALjnEpEE6s/zGJoB4xBsoBX0dqDvnxjfriQFbrmxymA+4A5+Dqc3IYQXc7CsyXqu9N/cCi
uxjbt7ginqPBtSp5mSoTtse/EFenhb1xHSqwWXMsoU+tCe5b8yk0dn2DS1TvVcIkpgTF7je3cKz3
uzg/V4AV/ZtOkRAcpRA2QPBUCqCT3WZJIDe6yUKmPNjhQmGIUQBwV5rZKpAuoEZnRuQCnkedwUmJ
bfRiNjf3VctQCi0OlQr+RPwidQYhOk1rP6anM/CtElJpxJKgdAgc08BlNbbOpJ4mbrWGlwUOJ6IG
zoveyWp4/gpT6zJVPRVOUfqCSkRnui/hT238ZHSYqyNWZH3ldY1TJZWHgkdJgdHgc3xFE6oD/o78
98y9lmOIQsIM4Os8wjq4ida3ef95CnYuUpTFGtjqmmLcqnFutCxvlL4bY/RXSROQodA1EJU4gFs9
Lb+P5gubod7U5Fs20Amj7UfRyEB+XYkm60ZrsYMGg3N/3dhugrQ2CtUz91x+tbc4LIF2EATVd2Pu
9Np9S3KBz5KGv76fuCuSxap3n8Sos62bsejAO9v1wAKra7v3R0R+8zFUimP9kGzXotV9OXXsXiqR
rVPIAt4MGLxjdzvJa/B3U3aRun0aOB+DajDSoL3M+h9KB0qeolpNhksV4h9e65ssS9DUDpv3HrsR
o7snO1NyrKQ740urqiGluMsfos/13ujxhmkVbJqDnnfnVhvmZLIq1z6QTk59f2G3riLXbYaO9SA8
dszQlSKlRzxYGn1ytH0wEcdypfn/2wSDiaPHcBiC/8B95IWjs5iNWkIb9uVzJuyIVo6GWHoKXomr
ovYvIVcD5jTkIdVsWKFI0pMNCoXXrh8jQWqBq/wwunZ7a6JKP8Xoc2w1sPGGRzb1/osOF2mZW3XL
HztgaVmCbTramRJ84gP2X3Sx84mj/gsDMaTLWcuuyN7beuHAnxlkerrBYKhYMIk6vo9Zkectm29k
UJRHetsZ2+AHcAWRw9O/nTshBdwG8GNfIhqfk0ExZ33FLMkMNPUpCpnvJkUuao8aOHCOlV0P++Q5
NK/wuN9qbS77Fbc5QCOWf93LnJLmi/98YlzAYsnvvVEOor3JFAsm/c+hSenFXyr1T3NA7J25x/3Z
wwg6AX5sFkBQG+S0/iPAkcmcb73CpA1C2AQuory15qDNcd7Y/mXEAMwPJQIhJrWqD3NLo8WoftCy
JDAQoOyhCjIL/FnOZs98ZcuY8yS+19eLAH3tHUoMZXKFuIGrWXVtMC8bXBWyqilmT7ZTjkAivaHw
PEaBq2zbW30AzbzNlDJglpk5b+f/pTeMFpxWpWpwWM+sGVlNNfgUUGRSgtNu0nRFDxU5hHnKmwFA
Is8/fg6YEk0tk5p6UE24JQZOqTF6DJt8FdZ86TUtjyr2Qwi6Eyx2hzG2q2wu8hGjG89qPxOqggr6
nBwk1m5LWMhzPpzeprrCzuweYC6nrxqehZZCuvnYN2JOLaVg2fUdDUBgbd4WVwJRaaLr4jGYxkdH
0Ou1Wg4rD/I8qjqMTyVqxzYSspNYP7gszAw2TWGKFrifZbTTsFLqgeMAPJbUixNqqPaspx5z2L6+
6X75MTLEF6XZ5UdvU+2XtU9+tKvpenwNKa+FUHykMKoChlgBxpanPUNMxFI0IQtJKX7gbUblVz8Y
K17/Nw6cgRgJtrPTkjpGLY4mLf0AcKs2+CsVfFMQTQQRkoN5CTL+DiKhHFKdSffzsrEmYYaygtre
FKNWe8PfX1yW4oYRgj1n+gMy5aDNYnsTez66x/xctOxLXsDAVurPnc2g/23N8dLJIDMAq8DDCq6P
d7bviPJ/OaQSUFicGgCFX8+/+jacDOq7bcxa2Fwkes9euSSjOnwS7Xik35YXOV8IOZvmaY3g8m1u
08ty7wdziPDwglvUNdmdEWmk1Flac9ms2DlJNZ3Fxm4jGWQqe96V4Kt+o8kp7fCQJQJ9wryiscEF
z0Whc3SK6sbWFMy6lmfimzE2RPFim0pEtIYwiCYChLesqL8nspqFqbXJKqsqwQtwRyxYfugIQMYp
2e4mHoHTJi6V8VhmXIr+zcLJDbTZGdGFp0V06H0NNnC+yWfc5sBdAohu8IZoP2BviRw59gLFHrQV
gs8mVCnE7aji2fgW5ggNPbLyUzS1TmwgKh1Iof08Nh4TYCzL3KfG52cLT5WyPlYE1F8/0vUy9v75
FcWOUvaXejHh6bT/M28xTlpJEubjPuwhzmZhCl+NyTs/rJqtgQD04e19m5kKOI+ETGBPEH7mYotE
cRinmPBNyBsH3ARtGYnOUlyiYkQ2fEnfJoJPShKvHSEIYd4ee8fsCYybFr/0oiEEJxxvs9Rg12UG
skelrxRqPTTA/ne3PNQFD8SyNuBvbxZSpSNK2Sycb8dLxy+iTSfvhOIoza9Xy864iwoU8SBmGhy1
XwTR+vPk8TqimolrW3+bI0EjtgaK2FJH9wlDkmYXDJPO1vbxXxHQcZr4jA6X1SsCTuUpW8wc6N+j
r8oFFuuaTjD7+TpEEM474GkSsgFJidGVFZZNPtd5yxNhuymCgYwDWT23L4BaJuBDr8abdt5b8qJG
XNxInLd2amMNGMj96F3bbX/v39WJq8EY9LM7W8+hqM5mU3tSF1hnKCwfUsfS6I9YEdm4dGiKLSJ/
1kjtseVyoXejoGfmZLgBdC1GV5UclK5D0mwZCvElSB1yLzssvd0XVnq7FPpd0iaa5SzjWW8kncqO
BF2D72V57XGIYH+NgIjpv+KQQo9KuxY0gZE2j4/Z3sHuKSY4PH5ZROj7A5VolDvhQAsF9x0+RAGj
droO3lPK0pIAKWURBXqvB7bNxLFH1YtxGIHgbvA78LNZ5cB7iVpLozF5W26g4xq5jISSAnJMNvuO
FZIDbux8YhY1oZWXtSe7V95sWLmtD/4WLFZ0BIz1dwBabGVmYBrr4kxYrLB+dI1tZuONO9vtOTlz
oOlDnewQQPrBxZFu8ICEsm3wqBVPXjmsi/JyOXQrDmMjOHTMAH7wIi32oS2Tz/Wlbtn3RixTbPEP
wjwORW/pbcQTPIdZaMx2GHOvHwhClxTjr77Ogj61s8sanzYegmLJBJj/fOMUAkssfCikrRrwTAS7
3U4Li9ZRbYGoBb1M069WICfdsvt74qVZvqNdqFGiTynwQyLCCb1rDGZlv5oUWSXgq0canh9Qca3N
DmyEPRaI62HWFQpPqx7aOxlophFEixPkIQttPe8dJpYOvzvh6FKJSmklu4VJCjA/Q0+BHpKrNgFC
cAZELzW7a5gd36/MMmsUxZ0FKZ8BTQ1eovQCY5I2UlOdEL5e5Q1Az+kzWvWc/NKjrDhsWl0QRvXj
hT5E1zDjxBmOaiaeKIqukL1Vf80Dfv27ZQ8DX5hGmJ3h6qgWLfGNrDNG4Xvu6fnkyHDQ8+Ck5sen
QEbo8YJyE1S7W4arbo5mVVSHUZRY9rpZbbfrmOtw2VLBgeq17z+vlFGlTyLRY2goSjTzZkapnXUW
r9F97TCFqlFyz8ME5o/IFMNUpjfi0eYvY+nDE6p0FSCmqoZqNxu5PRHGHZaxyAQSmRAe4hSdcvRE
vONxFJ3CBiW9CfjsgJ8PNE+KHsMLHYOEb6WFACNdrTqW5Cvke7iJ/CX9O/TWqpKHeOXmsP0UCVkh
LQV7TeDivrQsS2gCrbsxqLSWaBHfQdPb0ToBPBZE9hiuj4ZxnywPgJ2G1eEnFdxy0gLDPUnkfGv+
3Lmfcrbp6wL10NtamEcBAliGWmRKvs3HrBKgwh8KgjcBuL2exB7A3uTIbcCFVoSmh/sNO+ChTu4c
UMiV9NRJw4MWx436QwPHk0vtBmJdge+cFKyAo1rOZkwx1ZdPxAuw6iXplwiRZ+738i/IuCvuzil3
r44ViRxIxLNjyZ3zT6nDIolKYH4N1ifKZ6m1yYE5PFIWQcD7h820Yd2mIn9FOa3lq2Qr5oysx5i8
pmpcHW7qpzi2unWqk69P1B9GmXWTsQWE5tcXNlP7zEEf/oON+nplM4XvT7/4tDUkWblm/ICI2pKW
HCJ0UeWevXch9p9Kq9evlKl8ewH4IpfgEqQnoHrsJAv0saw6PvI9L2sBhQV0nwgjwZ9FadacjbSI
va9KQGUO1IO5zpyGj+9+EFpLJPhAQ0TZGAtmLVCLubB+e5RysRqx6RV8l7yvnFX/rYeiZpRKaBuP
1kKfd1RD6sCWlE5Q0+5xlf7DIKJMbiNjBUc0anz4JmxcVfQjU4DpoevArx+R2T5qPw60xWNfDsji
/mnIwUboumwNCejOGATycyBWyCg5XK5s/DF4wbxzc8PZe4P2XIrgkXeritkjeKZ04uvN8BAEUrBX
Hikwn+l4QIZIRhGKtjUSQWzqy/lfqW9wrACq1qNxl5mqdU5lR28vSs7PRwHyEQ/XpsbWVo/DjEzs
WUS5qkgA3J2KUGY8ZLqqB6jXXMz21GGJuoVfnzTKeGsCtRaG4IMlbspdmr9h0/sBiWhefv1vyWyH
5PxqafqibcpDSh654J0jaf1VjUvwouPqEBV+hMoWN1Zc5RlzlZAQiE3jOjc/E994C/JFEE8pcbVy
CM1ISAd90V6fenlHPssrkn002Jk89tfFTZIM68evVvQg+XbLrkn29KAcXQv6XpVpY6LhC1h/BAEj
YeUeQlIhG0Hk5K4cBrP4QvVoHjLf6ceq9+JWm1iYQeMJCSMwmsTSm79QJujeTsFrVVPFYUgv6g+v
fyslR/f9fLuMWS/xUdZCvG4/ZB1bpLowEId8pAC55+rJotvCyXtLNrscPaltmc9I/UsQvCwhY7I6
L1txeKlmaZJstzDcJoGUr61tkm1qL+AjUfyILWbN+7HkNyHqKzGP0UjSLtqMvPCGSkVXkNlxu0iY
IFA2Uwq6tIXH6mUA2ag3iFgNZbMd7AJBhZeRMpvQYgeqcpubcKuo7FGbPJyeXOHaGb5hGqazcSeg
mzsfaVPDILJEZPkNdt81MHw8a4CE5IFOF1wFQtXbIpg6x35WDdpQ9QatAcW3eU9cJORYN28mXgNV
4E0ise/yDoJE/St4OBunjPK+gxzisDrTnAemOYv/dd92K4aC31zA7U5+IE7cH/pkxB5PMRWWuoRE
uf4ItkRMFxWu8oPrKy1E0doVR9EHZeMSb8aVlGLcbZjdnsfazdDR7jMkJifvl1vB+/ZftC5OCpEh
hn7GaoApSI45/bJGx/PZiEymWFDhFDmWAF9ba/vjZ3VHLX+K5WX8F7JobB7f1FssQQb42IWc5iTw
exB6zkLoOvUApvaHp5EwETbSGaqHuGylIT6yWgLHKut4cnxC5gmS0eC6OMxtNT2wpHb0h56GD1TQ
huq6nQW/Dl+UwLJx97WHtETzsbPt2MTi0M8hHjKjECVVZVnnyMglOf5GXnVSdbfmlkH8y4VmSD3p
qhHcGfJ3n1zSQxBD0Lt+tqcjyLW2lXT0WTMSmHANrSpH3Wm3u65sRfAhle1WkZxeUcBzC3LWPQji
JXsOskoJoj3pCr9SP8/dqZe6u1/SMt/hWI7gIFqECMbLO3cFFYVXSK+aCY+5XDiotzpxSAzNoukC
PuioCiubQVZBTCt7JhNMN4dsoUuaKHV9TW7uX8zHm4kgV5UhkhYZBf1tIvdj0LLsETAFWhJS+nCF
qI3Hd6j+hJEf9wjXAjbfmfbC8S5z3Wqqw4NpSmm9wYacJa4F0FAfcMfpdnqB9+rnaUJQD1Xsir3i
PuhYWyAipxhPywHcNeSemoPIVlrVAPZv/FGt4uON2oOJO1Fxmf/1+fkxlii+KxDutWE3k/iEgPYp
eRfBaWW47K9daJ8XYxQuBG38PCrKRNm3VwJFN5A3cYdMoeM4BdnyTmuRlf+ytnXe8F/+eFmZL0Xv
bgbeNAgWSx1YhLOEnhNXN2Bd6PQwivuzjeF15owDnABDnYtWAjWuFpXlJ4JSLehOk/4VKTOAHNYS
P8mkDNouzbdKvhRDNdm2rZmhfHPHodp+pyDGFEs2n70Pxp7XSRUiIOXliYkVOeSMih5UGh9hC5a8
LapFxWgkqU2aF+x77Pt7JBbhCSQ1UTaH1AE2Me+mdeWCCNqQXfBHWoMbl2s9lTq0y2AEbLn6aEGJ
RTAejX1SlVl0Fgvfy+95O4/Qoq19LBAJPbmDoSD87xq68vCysMlK2ZU3ZyiwG5OhWPiU9dNkIPgL
TS0BGBf/QOn2AZKyFfS7P+Oy/qDZ+P3wfE5OyOzN0RqhWg6jmcrB5qQqy87ErURt1EdYOY8+DL9V
+CSE9Wgndz0Svfe5iTL0vDlbFpLRMOZiWa1fsWLvh25L/kG8WGHXhasNQ3VxK3VptxgTwn/mu/JS
lMExqTPxbMwiveiQZKSeUyY0Y9mCAwCH9JzpIZshpt+YKxT9IHenLeJVtLb53MoTU9dH266oxV+y
aPqR1XkTK5XBEmApfKRKo0uWWWnrO7lJQ6Zjgkk4mOURG3XpaTWZ9nb/qMruDJ/in2KkYmslMTsd
mgRr+RbO3DNbGlT6lmCYRjyXaKI7uRRXcuq6lw4dE4OS7BdU6izpvsBQGsjQ4eChy4rywF5CuitW
Ul7lAx7HVZLPXn49QV2JkZqi4u8OehT+CpDYnnVUj+BJVtQPS6edxsuiDch/bMLol4Nczl8m/O4b
iC5dvSKuJBo13Lr84wpIAg7xQJKziTVjmRfP8TmltpOqnugO6PDJOCCx1vl5GRCqU81c2SfrZKyv
XLwbBNjrJNoyj2veZ4JsCIs73bo1/PAnSsawFyDUC9S8BuMzifulyL25J3YNADqqhvudPkWLOY61
MoZHLsZNVvssRbdhmdGgEuDZR8X70IqIgPX7/p/1PYcAtVrBTyZw/85OGH3La9g1yy2v6Wi6UPrv
DC20PyqXsxW4gAU6jxLlr53R4uWl/HxKrWaTEbBedMIEoLLwdCKc7C1YqNk1aIe628IwlhF9Khby
fyAFK1X5LSj8QOuuET2czkb7aOMJgMjIF07PrRUzIIOs6IxhGXuP4V6WeMtON86JuK/fp8Bntooo
vRK4oKW8MAHmjfV3y7VioBa1k5d+9VKIGHIho0Om3925tlMq+yvrHFtK/ak4vk75dwxktYehp7dV
UfFkZIo9pah8QgT7HnlZlexNhUv2eoXHEU7eqthIhCyhPXhZjUtI97ZyiecwaDgbxJUnrbKiQMba
b2i19K5nhB09+jMgz8OQlyGTj5XsOOwTizDALiM7Etpi3YygknyeV/sZ+xJ3aVEewWUlfSN2c2wL
WDnj9LLO0Cz0unrQjrZbvqmUiu5Rhpl7Gdoj334VvkkXONqCHC/W98UdRSsIfvTyXgD1ZzfZYthH
kWonhVJiHFdVDOH/yAi2IZKa39Zmdu+MWt+jJiXW708LlJi/AZubY3M1hSGBI6Kxxfip8Jl5xDDR
NwFtOAhYgrCqwCMxvkEt3E4SdRuDP+LwpTF8R7rfvfFQXtNEFmhmvPV+GdUfzWUYJatU5tpAKfKp
eL8eg00L/Azo7CAWVwdY6GB/YD60MrupMiW2LSFiy5YOMRR19dYfqyZJ35yjKuF1X2WnDfpC4Stn
UDim+GmWxs5h5PvlNceC7+ERMoap/PqMFsFs1eo6nAvtVZ1fBd0uIdL9Y+6uhdHV1CgmNAnd+1GV
kctumjAnvY0K6Wm+Ppb/IElY3rktZRwaBQZLgsxMQrRQko25Ny94UV/+zO6CBLH5asXMzX3seUv6
z5YXEDo/JrGZQDed+90zznJTmCEFI33yFllF+BCDgIdJgmO1R4ZYlE1h7vZl4IdzPw9iz0o1ZwuF
N/lK2GtWgheFB4vFbAiygRo5mZ+pnLuA16IUDm6AzZEG1CPwBUT3xeQDLsTlxIeHij42MBTfrV2S
2j88nepBxUH1eUvGS2XQiQaJ/tWAHqBn2r3NojBsR+//tyLd5ASTgKPwPSnNc6x/Ckz8I/Sit31B
hHhUpIgP66Vq7pX6xtCsL8EaP0pvk3Sn4jm91xQdx2QSeJ07Bp2S9f9UgxQ2LitvvgA8x3Sq8n/e
8OZxY8lMuOqKZX5nbgUMZKV6u7+4DdjWZDOYmaAGjjS88eW0/4/3CAjxca3569ZA5+ty2PzoGRT+
uU5cbpwyz0XspOnYx7ll6hPSDyBx57uGVExVkP1BIZFtmnhQwbJRUUIPPni095KTi0ECepqxUJzB
16wEOs6KpXaqmOaR50d5B3qQPcuUOaj0HbrxLGWuaieAdx8eFrnwYgUok5Uzb+0MV0ewK5DMEDgw
cRsnwCcwuNNZwOEXOUYbp/NlTW+TIH2jCzhYGYut/m0pLUVwSWXX1lEMohvisWJ0XaGE0FurV/Em
i10Gd3ofxuTcXGb5wbpYqUWiE3Kob7UBAcf4HEFYmAmuHoy7Y/wMuLlSG9uwKHyAcsEqWG3Em9jT
lkd9dLnpEbUQSiioE25QLzoi9eoma5RoegJyylYRZ1kKaMPBigHCxph0N6Ssf851wj3+p+98QL3Z
9yoyKrdgaxEPYQOpOgkrIIsD0WUMbXT6dnyg1L593+TFRyxOzGXIER+Q72piw52ggdifDCLNF8il
Rc7FK+ipFRkf6BtOJ7lSsG01tjxFSfnUW3B4KfVRdg83b/ebf43HzyijHcSes5CFJMiArQVucw+t
ythtYDgEhuCgD4YW9ToNESE4vccgAWcJtREafAV7wbFNHqtT6hXK2GfZQIdQvGzOsHg3gMLci6Qg
D9ROjINd0kPBatftNBXEhSeV5KjbEkIOBsrlI2JmqMJ6X/u3dOj0xxn1/J76AS69rxq2h3k7K06k
erPUs+zx9/AGGvJFwQHp+0hRXhtQH8AF57weINHXh+r/k6Aa96+q2niSYg4AcGhucYe871KIb7HT
45u/UQj4Jvhi5/l1eJjId4VEVioBSD5n2GpEMN0g86E7s46bLlA3wHhrAaLJLqHsB4jFCBAnPSUP
+nuBQt0rkBScfeZhvmYZyGa1sJYAYWb2J205FGBTPuhd7qJHEuQRx6/C6YkU4VN4czhIrxHAZ4zy
j4S/YNm5HlkaZnK91uSemwIKmUDzd7gOB0ghvtgMstL0zUDVLVZHMxFQLni10aanzq0OJFeupVNL
CahmI5L0Mz/TqqJqWLXjG4EfN1Z/Gw5mXNOFCqeLRtUjznQJ/E0foyjHxDYuHONGukesfxJzm8qf
/Ht1IO8+nhHVFOcC/DvrR6tzh+vXulkcode6fLGrABhnsxb5TsoPlIuxhPrIdfMS9tOsarQ8QVJo
xtAyVK1QvAM5w91koI6+2mtEcTJQOWrbHu/Mperp09S/EtRRu7/bXmHqQkmOoW9fthdNzwpVI6Y2
ggWvBaMAW/5nnnpFHq/6yvWUlPhX4ZI2lwSZj+U3ygWwKtwWeSkHzNjd/uTfbE+a+Y8wjTTTyPNh
oo7gdQxl6IG0qO2cPGRozVvrSg2ZISGokSWcmdoMhMQvhbe89Mrsft5X0dTIZ9gbE1jc7ryXSE+d
3eMdH/jqq0hWSIBgoUK0IUZJOZNvBDGDJ60QucULjcdujT0YsqMqzgap8tMln3mF9sEwzT9iADtc
vbw/jAfjk1mM3uU39ncnyfWXTDdlplQJwcqYFVP228NMUnEI4oBxZ7h/JWgD4LLGmzdhLkMirwHq
AA5Mru3i7kphELYhs8mjxANFNZqHn+eVVNmXtfPURnTUcQ7XB02dBHBMvs/XkKMQKh0Wo4T5Ym6F
aT9qs5vY1Xs98mc99IMRD2MTZL1WJco81D9Z0/OJUzJfF7qNAhnulyKgtwXqBCDxZlAgmU6pE0nZ
MXAEnwjlT/emvaREzrsFOgEARiivdTIvRU2L+vLzcWygAdInKENOpXTdcr7Dl4iqMyUBpd0Af4GO
kh0ppWFDc5Hutxufb50m0pHnFUr27p0Gjd9aKFUIf2PQXqvqAMBRc5KGoxA/Ct4Gyf0XAQP5gO9P
/2Gs36Hek8RH/7PKk5KUNLYMLjKF9kLMGl7c4Hr2yYLqbSdMAEN0xRkRCz7kJTsRxBXgnhpvCRmC
3DMyDWXm3qeLoTqtp8B1vtFTPCdJasSnRzLwleDBCKFySEeAHxboTb9IP76VM+ddnnFNeXMFlV3b
QkSwlLh6RV2DK9Tv4IuJAsjUqFVsO3VIBlC32tF4eRAlvJIGbVOuZDrFziJbdTjq0vkLAlVlyybN
eCsqVGzNDUPkF8HxPowgM7MgKEseU9M/A93rPL1TSJP2JKEQ6crZRPvfrsKrW2Ov+3oJbdN59tge
ShI76IJ4Lf5DgllnUSvw8uuuthT4F+UsIVJ6JsXRwmyqxfFm4JXks/aQVNKPsp37bievqlyNIety
+JNXNZYEhotEUQ/YkdWBxQpPI3EczPbViLN415Fux8ZTpFCK39zoOkrFlA+Cs8BziqNpBOgm3mCc
U0lza2ciQEdpzclMPE4tAOQfDRL7kDGbGk/d1kXvXy693ghtjD+swaiubJxNsqB+/RTI86GCOwaQ
gbHR58cPoBZ8dOqy91Rj83bMLzY6JtOkIFj6mxPFkwuUJA8uqL+9UbNNlGpow5na7gDFsPCUDuhR
yaB+8XhfwW20pyHPlX0kSKjbp90t7QM9dMI2iQ/pbHQuY2/5lV05VL5YE0qkmwry6bO+zysP9+hf
mUUOaNdKAp1V/Qkv1B5Fs+OYDHGAb+Gyu6JOvm57cx+1hU/eGHLksykgR6RaFZR4Z7+N2VkP4N57
sziUBdRrPwS2oKpHXl7uGI+FEUutbBdE+U898Qik+FMGoZ2L0RcQJ5CsI/EgJIggFBURq47DSs4u
PdUQtyYucPQba09HBnMSlBvCB1vST1AALDQWonwa7x9TJVtA8erasQq4IVL7wPYRbE41Hq2brRwg
eyCvVMU6EMcd8CmCRtSqRx0kxo4PmCP5VlEhd7Vp6Rtv9XGfqzAeEHedCV+fAAZJe12wcJ8E3qCq
x/14LrSU0O8Fl/8RLs2yyP3+WezgVGtSVYn7SwmarSqS/AR1+ajY0Ukzr/WLzQuUvBdirpYefPoo
Ys1wj/ROvMv5aJ0G8TBSV6MV5V6V0YkpkujiebjrwSrKGHYknW/JDC0RYgEEyB7rNnuMRX46deVg
bUlTvONFHQVNSF1t5b0fwAZqHi7NlVlrRMyH7m+RyOhUWC39z0mwRZVF2H3CQp9+7Prsn2BLZzt4
tpcXBPE9nSPfTcA4Bha4x8rk2q7qc19ffO8P6Z4NpJG6RItHHroJtWZwrE/QA4Vhk6yKtNDmTWEg
TVb9mKyBM8A+RCrXMCePD9pOVv4dEYfEv4gbcKvFQhjcQWmCqE1w8J8XMOGJ0jXOirRgO7x36p0v
p7y9dKtb0nVeYURJGbInB04CQLawdiJPYjo9LsK5SciYvsjX5ig8W1NvRdRM7wYsgcVyQq1NcJz+
iWcNh+Qu86/5dTF9DReI1vS8edcN8WEZveglWZFoku8++VDzhVOx2W/IRsQkB6sOGXdng8WFusUo
8bSlYiD3KfNm2MB96sT5X/R5rRIjD/LAIbK+LPHvClBnlaziJ8xJa7Y3b7at6Hoz0jIXcWMPc87r
Z+vc4lSHWvGomNm/tSeGzDX/G5z4wHT66XMvsOTvKlWfL2v1HRKiIShpbQahYI8FxiPo0BGnfVS4
Tjd25JCIo9E3WJegA6oNoC3He1+h9Dxs5qdd/jYBYPzuOsfxqBvQE18QpleVV5SDAG6XtAEjRRgo
JZwB+Jj3+01q32S3Y3xaixNspks57Zk8iDUmScsCe0FLwKj9RgNsuwk1VlmAmctsMfnGiVh9Ov8+
YaDN6hgUKhABBvQ79qigymfMuuVe9VEdO8PHstYErOn3ao1hyE7ieLzEtWYz4WlxEARZLvTRVjEi
+eHxy5F6Sa1JuzS7uGGkpUY6Vs0yii/OxDV0vv9XdzlojqMwhlFBn7uQ03nlvdtAdmPalAp47Qqu
OHZWadyEhkw4g/Gv6uQM1v01ses4yAL+IwjVgUFa7oiouXXkqRYvdTdK2eLHC9z1bTdXHOChD1ws
U/ed/s3krpcTy5hmFfHF01+HjJZMZ7aIpBEoEyOko0RI7Jdf0Cb86lfdCOHhOqJJUO/c/oKgLT10
a8j01rr0MecH1yTzXyEFGEbWRZtABw7VSjPr+6TRWz6VBrLvu0EcniV417xPrn7wFp6Os7SMxlR3
pIxKyXs6hZSnNp/q/NL6O4tylkuMjhiFm4tKkyf/LPqhEl51tAqIw/Uw7gLlsIy3PuVfL6JGkFRA
/HMYkDu9jbinMO1f/r0TBDeVq3M/9Xu4rNwW//UPPSTGWP9cxNtttLka6wkdabbCJJzTwXunx/cy
cn4zV6e4sBnAjJhTIBuVXeMmmuRfG/BtD25iVC4Q6nb/lpFYHp+pHSzwjtGc5J/v7VM1eEx+n3GE
HoDDLuXLX85WzygaQt6k/5dFBrtswIeEtoYbwTpYIkpjRSGVd7HrTQe4coUUlrnB3jO8DVM8ijuk
PPQoq95PmtNhC/ggDjSdhtJd/SF1RRxb1LyyuuvgmYyxGzHJAcm527FobNilvhISdTzI5+3+9NTR
waOULoDREn0jgHrxyAhdFRRh6wY4GeYIFbg/IxGrrjXLZmGd5fooQzqG2f2yCScdnaDBFBJDJS3f
h6lGOLNW3bJLtwZANrDfYRk+Fr3JkJSchah9q4TD3IXHNaW63q49iD/ROvpKsuF6egjIR5hVgaI8
U075uoebdabD5Q56k4dk26kW55ytXWIehI2G+6okXXsPkPuPp2MnmnLgTjttaW5mnGO2kq2g7KhH
wIO8vPg52EUeuA5Tp0Z2pyqKqwZOi3jl5kar8b3CmNLjBrjq3kJ8P7RpJGQzbM1ZaGwvzxQ3Sqxf
0Dfu0vkJ5PZ1tfq78c2NuD2NzRtKFhT2TC5S2p9SzoAfntdbfUvIZ+4UO+qMb8PwVFwy5Q62KQGu
vrjoa8IkqqgoHzVXFvrwf1mmF/ps09C/KvG6vEPyDtkqNMLJGT1RlcBegztG/fZONLRRwom5tb8l
RuuTWmb7wStAWPn4ePTTewNeqfLQsIo/WtFK42xnD2P7HdrxVfVggaowNcMX68qNwBDeROYXN7uB
Ls6lV1iSu5z2lYFNmT7kaWkZJAi98wfzER0v1fHGAF1eQ/xtjjt3PHd6S8wR95efSvaQiH70AJDR
KKoj8zkpskCpBOBIW/y6PLz6EnuxCvuDEErfJ6+kqQR/9FK1+VlOGiLMYXYiuwT8nvcsFqOtHGe4
fyEBOwmeT0ljdAT/XIrXw6TVJQUcm4JSPZT1iRZEok6KK2al3cC80+smzRUMU3EZLGuxT5zM8ME+
jsZwb9iMO5hcf9+Yvvax/A4jwqdw38PE47aUlOSE3yaJaorfX6nOeHmeVKTAfWmP+pNLFYVDlZYE
/UMEnQzdnRaEONiPpiqDVFc7aQ0mx6o2wPyDQjH41pHxkFhsLu0rqHFSgkeijoj0lgGCrjbOIEn0
YbMhdpgjzQXStPBucex0hgJhfmC8TUFhIdzuOH7KT4KLW+Tj7kHhUExnNG6hJogaV5lTdITVV+e1
O4D8lhsPVpmw7wXzzopl+m5wcV/moa2GZjWJFConVonvBZSIUTGQmNUipw03w4ZwSrir7I52CEop
Z53F08aIki+B6O6KL8Vi97S/fDk5C6PzHN4cHgfI0nYnVTdfOz+7UDF1LWQSvi06PX5o35+BHwPh
XChfjHsOYh/OL5Xi2ND///8iVEy/5L4C8UNRWPN8oHjjPfH+/3nZLG8zJVZxZdfcYX589BPP/PRy
sIVuq8hNVpcLKdq6/t2/n6w4WWS94PcDmYUyPHQDEf7SCi4pSX8pGecJRwnrDbUfp+rIqNnv72cz
f6zKzexsu/yqofVWg7gsdEdtW2uo1w/pMmo4mpZjLHoGeRiz3P/6swcefvi9xVM64uJzapTjBrp6
qVvknY3CynbyR3JqKEkQxrGTOzs07NpK4ayVV9OMB797hXqxSZgYNapH9xatUxwEZA54DcOBw65O
8ZAVzCSHiCG4gDfo51OBQByiJAJgddlNxZzzeWTEa0ed9ITlzEBHka43V//p3xt4WKEsALwVv7O4
1L9cYo5i/ol9TPAbM0vyO1Eb19T/abIfUYw9Bj0F3y1l1c7xJSUIoxGhAHdJs8vA7K/ynHgzLrSB
l8sXfcUbygLRfKte6aonjUc5bJLq3u6tAn+91mUETGacWYX5EwFUcWKgbLSCvuhH7pJtihTw1t0B
3YiJ7JzfycqgfJ56qveVHDWWVijC3pOTookt3NVYc/2Pgfs9D4VmhHanxU6mOsw9M/h140vwAkfd
FgEWd1bSF94jwsM61VmYBp9abeHeR/DnDFpD+8hTmJeq8tEY1ikdm9qaathKYbLAWR+MenXlsyvo
+HpEgDSULnu0ady6GMLPOx0DhsfREha1VSpX76nnzVGV0Jv7VPtUkdEvdINGrjh9QVxRc76s5d3a
3ymP0oRDitAzfj1KEdXQ9NmRp3drbc9osBp+Jfjb/7arJv6t+4jU+zbBswvBHLmOzlEuQrrytH/T
jBc0L2fKLSCw0BXpjJ0FlpLZULq9FszsvECtSz2lcTR5kuf/QPotMAsF+g8r8sY9PJfUEIiOJ9Nc
NERtQI9QvflufS/90Z9NYS9UocOp0qregpCLpPjntnBkX0xbb5QNdBK58/hnjRaZo+qiue3MXQn8
/evdPug5egC7S6TQTdmt4SeAq1oUhaqReYtgH1S1FcPUF9MFrOZrVzrLyXEIJSUsmxSisSOLCHXI
8UsFMjfTtIrWqBvQIPEp8MPJMGQjEAtN/N3b+CwDJD66LsUS3ypGtWeuebr6E7LkWWk1oF8b+2+V
zPqoeXA0/H8HXkjn3V5Wttkp/5/X9kmRR3C8Rx3ytSbPSylwdTsCL0JfnVDVtCbkmcwGMMk71IJ/
iTwl8IzZWTS9wv2Zfn+lM5OAahEL/xbZAxqTHcInuyjydhUkqibLM5Eo8j0da3Bsx951vAghre0k
zqmzuKKJqwOXX1LeY63u6ILsyRie6/rMf6uEZXZCxfVlFcFPyyHFNHQSMfToJtWP0QPchx4/axyc
Yo9ec31oUqpOL31lLIBZMdM489CWA2da8JcUhYk+zh1JMVsNtzrmnt9GUM3/CdGRwpxBaR4VKd+c
nM2iiZTJwFHU/SIYKwH2ZG8fBuOvPdap2w79oxra5et4PqKrQdigWbuKVra9koKnp5CWPREumPVF
LCIbcM5vX1YYk1r3BAzVco8HqCJsLy9f8BPhgzUBy065+mNDxdP7L7khUU5nzENczZ011OVWHGNc
nqtEOzXGIh0pHANbH6eGMNyr9WgRxSkMiOM4tKfEkxQGFxckIrmyBX3tg0OsD7mHN5aZN2nGAfG/
y98wr8/oYUoiROomnrHcwuiuknJvIXoCt2zoGKAfoi9TmxbK7iOrwq794noUrbBRnHylcpdPemGX
jg7L/mYu6dCdd5TGC3OcKR2ZlKD5X8Qu78VGoV0cPMiB0xtFUq9TuevKIUPmY3elt9BnkUWH9A0v
AE1AM85QFO24ZqQCIRj+bTLHXNBxpYJhPlsfiRC5GXKIcBc0WkTVuTeovDl+icvN7sV1+hN6F/Bs
hgNkjFTDAFSwWxBOK8h/lEUzk3Vhl6gK/kty9wrkuJ3pVGLJRIApYngddWcP7u6XjpNPeVYRV+fd
448Zeh4q9Q24UBzyN75vtpsguVpZ83kzvIlYvim43OknAFfIhyfZ4CsE3q7pcpunKa5pXfnlKmjt
mKtWsiGJ2qlGQk/wufrb64mt/tN3bBBLzWv7lAdn/GTW2LIheE41dhfuweCyGnG7REuNPqfv/rSz
gDaj7BLTU0cyfUPoOf4kiuMJ2gwPo1hUhu35vXg/hmagkE39UXTYRy/aJYMBJFeoSzOp5gyP1WTr
VW1CC9Cwl36BUtMkmvnudeyq1EAEPjfOcrlkcjCN2VfwEdlp1pMOgtuVxe+3dRnBQB2kd2sP13wV
WSBzDXzLU5+iZGbG8FKkF0mgQ1uFnkbvOJEoRwh19rKB+1n00rmqgd3+WfugwfbBoFFTkh1Ucdtp
SUo9OSHKHCe7Oaa0MAbHqTUuFcsf6dCeyJmVQuHIEFwsfBTsAYygjcNVzSGdREc+2+jP0aKSzcOp
Wj4KGXyb4Y0MvSY2CVm9ED1dshuHP2j2eZQEcuv/eNJnegOpWP7iz4atPE6hpaKlIfzTS0Qn6Lbr
1U0iy3xG90XirwLJ55QYKBJ/Ni90jbh1iBS+TIWe8ws9C/EbDaLLxJMrZ8WkGwSK+CB+cbzm6lg8
VLsj0LJ5HNl72JUnG0P0ZRK2UhwQeJ06lfW1bJyyNbBBQ2nocSLwsBN4IVUA3b39VZ31uboO7eD6
AY3NdOz1y19ihayIRIT7vLQDkPNpg52z8GQHvGo4fNzTNVdHtt+tzIxU5pltMg8kZHteWCZbUjy/
p3rQNPLESwRTA82QoB7BW8AkLPT8OKmRQA3sbyEbtc9uBIeusDKWiBxpCbQomquo1IjtJmnjOiNy
TEoFO7ndjtFJBkNg6RaTqPzmZ6hqPXyeejMgbPuMDiIOVd8XnB48PkLYups0RcUxbBR6gYMaP0se
zn44rBIcyTaqzs7vggJzf2F0pf/QBf/O21tkqJu0RYZ93FsxG7zt7NFyh64Rpm/HASowKwOVz59N
ZlSz/f1wVPMbmjLKfHaTmcd3I/mBucw/4rWPWiZgW+SXCdcKZBc1s56kT5mDDxldHUafiX8Y+hsM
Mmak8TS87Ixor8p2Rg07mYXtBK79E+YExKnfSFy4mZqMSieY9sAwdc9/B6weouJfTo71ZbSnuYk1
kjWoxvA/JyBF0E0ORYyku0oudfkqlNR6Os45krlE525waYe/REXocY2VkhyGRXjftEU75tTa5qaY
kHe5M7YD1yX1liy9lge1xlUPXmwhQTz9Wn3DIdN/uphq11Nz7yi470y2kToN71kZz4pW/D95/7WY
t80nL6y3vzrPIoxO+anN5v9K7S09jNYHXVshc/dI8EE0o7lolRB14gp0bd11DSmQkkLfMH+LaAoZ
R8vKSIOAo5p9EIEcWAvHziXuN7P8n+oDIg2eupygJOpYnj1yChs1hEOx0CUiLxXJmpi25cq6qeAh
fnYImDIJutm8zUB6PpAutqKHRT0cMnupbaruAkJ1KE3yAdEJCcL1LLvXWpAoy7KBlNlyhihsKLt8
zHnAwXagVqrskvluu0aaN4gRcB9uKgctBh9IMsYc5JBPS4pjqReIKQQn59RPEnphxOLbWQEr3/iU
1g4tgUo20sA32eNsJSig9x2Ptxx8GEvFjKvrKGYKpYCP/dnorecU0Y8WrurK2eXNqmCbfFRfNOP3
/HiFwFZxt/gj8CY0WcDwMSL4GWbGW0oB6YNI9mCYEXNtDPy5rVgTtFp9LkdcZIjBpdnJSV/I80Bd
7QbuX3eRZs3sK9QIlWJaWXps80Z5cCTdmUCbSe/WHMTjewdroMDvW6cRr9nuwOm1SDoZaEa0L+NS
8Zgn3efuVhAL8E1TV0BkOnSNrXfsU7xu4py3/1DJ5TPm45f1+EaFKcdEC7NsV6iNQpCM8IBskcmT
V5CkfvHBSaPF2YDxigAh+pf6P+ng7KhrXkxuvEXy7t0Akh1nQkASYYfikyEeQX7hXJzW9e3l9Iyo
AaXZWiHTjTRqHlmXXXeopSghI4YFC0L4exJfhdZyxSyg2VzRInk5y3xak5QwDK5PnZ9u+enHy9tD
W48eepIhqRzAEv+SBTLSsYKkNxmZwT3b4syc0WWu50sxt8ZKsqH88EKmUDaJKc3BzGdbRkQ3oC9U
gnHagojNswt8NF8VzLUoLz/Y9J7OxYLAgTLdUkOcVtnbzrrOeul5+HweHjUCCWej1S5736CwMkDY
Sv3RWVkhkiOL4RUQOTsVTEHlXvqqTf7PDKG/VKuvfe27Y0jhEZBjJBnplV9XtmuKHJs0V5JjU6/M
tzJoEJLY8K9wT2+zJI0B2p7ZCDNAsxxU5tlyKb/9imZgB8WBuERGG2fQV7UK3NkSgcIbX8ORZgcF
3OQ96G+t7w1/GSUJ75ft0c2fr2xxVLhyG7f6rh7aTM9PybnAYLiComCoOR7XwmHtdA/k/4Yvvx/I
pX5KghW794BF+60o6L/6QFbLVLtTE3RbScD6E398xsGRztzBAl8SCJ+QuDbvEoZ4KE9CCt2Pxl04
5VVB8XkUXgv2EkdPkIUodn7HLc5bCjqoqDh/GQMZskVVKka/FRVQDQr6z9PbiTTLSC7JWiRWYHgS
LDnEhKBQsX0A4isyLUerDhGQb4ORTsrBDlGZZ++jYCj0JzjAl5CEzzeA19vV1kfP6fKZOT0l1vuA
9W/mSZ8rKF85acH023LDHxUN8caYDPkJFFwSv9ISCqz8zPo+ViKAHAoJOwzyBnGkkpE5oWv4sGB3
Gw51xUtVz1Zl6XSnxu1bA3sxxTuREht3AVVKXAuS26BRs0y9dizYQyanUavTMNbxZKXKa27jZGd3
9W9EKqCrHlc/dB2pfLWsO31mIW9ivbe/ARGHt1qgmGem0ir8KahC8/h2t4ryy2pNSspcE5i2Gk0s
dJOMz0GP36zxopPFKhOXCWl2s69+c5lbxqM69vSeOC1U4lLKcbQCsSw5/+MA0GQ0jj7FcJARTsN0
oWxjNK1lB6Z3toZaMlRktoaXjQRFH6s3U+gbFBhY4z+/ICe/5cYMABHxRGiG31ycqmWyTCPEAQbC
Ru+fhfI8UjJ3eCtNt0zaDtYuaa2mtFELNWyF+F0dN6TaWbZj0T5WcSK3hOwvDwHGXS1ncC271BjM
braeaXiGltJtLp5LLqlvZ36z9R4J4EBsWPRvrEP0gjiGyoG2tiMjzfjjoF/F033T56+BTmdqbt50
jOuOkAsUS9YvTkw3I+ouTebyotA8auUAR2/BWEWCpAf6ARQujVl9JuvM1slmHXzFykF69rAFwfP/
rjl9YvthonlnQ6zCNB9JWf+FiXE0iUuvHYinW2IJ+Kn6Hy61dtexyBqHxeYjeiVUt260YbiRyJIi
wevCrmYeuXSH2mY7PYdYJKiSBtE0lkeQ5Qkt8iNhZhiENcQLZcbA5FtLPAUfCzannKl0hR5ennSN
QtRViZ12IlOTXpXxzQyCuSEXyr2UsQfusd36VM520a/9i3PTesY8zb8E+1kN4PPY0w0V+C6zRUAL
7pJhiZJtmb4qFXMvEc8S9cvL52CFjfRs4YjGEFrUtN+s6SfD6TPuQx7U1DI743/s8pugQV2RgzhK
RKC4vBm3tQtCg1A1iGBGYPvwv1/D7TPiSAHJeQiMWY/1jg9ZylHq4n4D8dYRV4TuZo0y2zeilc/Z
SVrAfrrAY99DsaBPZPPNn65ddN0qONPhKnMZC3DkgLU9PBYIl1dWz78eRIkcfd9vvi33H92++b34
kNHMIMPpipjDu7IAGLGmQ7ybdM9HLu/2xbMNqKS0plv94Yc6DalQsuCwLxsaSFi5KbJe0Kc7LxsD
ybNEpLpGwdA2YZtk5w6nXjuewyb1647iZJm9Gr9hbj8sWPslZUyLVHFTgDvXBzJLM1JjGpiml8Un
F8C7E7CVFdQLJ65CtQi8jCQV/B6Kt55gZ9QTaFOJCN5E4x1ybkk8VFe3rX5spuyV9onF7d4A+o1S
cOWSY/QoWUq56GGJID+uj1PK/LxzJuGnTP70khijcwokCr6rMdQAaRD8arpU9pwLeK/shqbJ3qCB
qESXi35Uk8PzRN9QPmdQK+VS4tmc12rsKzkExt8FljnmKEMPhdUznF+xm+PLh5lUXI16Uk9WXsbV
Mhh5MU13s0BwKsAEU8lNFKYoCXRIBlB3W301IHSZL7hO8VMmKHdUD7HHpqxu4thHRJcOwOjMdkjd
+XFQEfAFW2gj/ccZkeRbFvZvx9I001Vm5qzWTEveiwV2+sxd/7DXRXfbyqEG/HUopztmwy8sl/ju
rL2FL1rugnRyGVhTHMaEK9E9SyJc5Sxw8sbSDZZrrZ6j9emyrI+dnTZrUW0OVt1wkuEhWbCj6Jga
zqO5dFNKRRFxyyD7kfpCtkVKO4jPjKNPMHxzpIsSy6qpMxCG4SE1Xb7c7feuSUA63T4iDaQ1MGvk
iGJIMg0z5Knt1SnvIHOp0nWATKA0LTZZZ6SAKrRXgERwSyCZg+8YTALwfodOwuWLhRmvTv4F6B1Q
uJHAtC4lHzFBlFWacyNN6I+qu3minHkhpZMd5y5Ui6XlA4Ltu2XxHAHxSnr77yk2e8DO8Jm3krNp
w6SRD+YbI+6w0KwnmjhpGYfmVDlukaMyV435sYgBiPGrynDCrZ9YWqQLsBVNWP3yJcub00niDSIK
ovrwSOSXPFjTk/SXICYb6FgMd6P4fF0KsltbKFkc1CyPQkPz7fvwe+1Wdrbjwo2DCyMxzNvuf2ak
kipJHFp8HNhxOy2CZvsJXjmF2L2GXfiHr1qYy1FB/l9NkIzIpW2YmdSM5d1KNYTSSuJAGX1nbm4C
jGHJ7P4BQ/M3RLbrDyP2vGELyiwUYxQvMxur0HEu5XnFx+wA1gYjFmhtxs4i4amu013V8ZFsMy0z
G41VKNf9P2hlQRLyEYpkt9/TTJ8+8nfBLldaCsp/vc9wQwEz0lXjZYgXDUg7CdRwQn0Kq+o2F9Lp
KsDxOweGmn4UYKyee4DIM1NSiKkD/pr8kO6WL106Vl2WSxsvmidJ2RTeVt3t8hcoNMdJYIoAkKDP
rik8PvqHqtp04e4P0/E/dP/7QuyaGXX3a624EfdDMddsQxPcJi7xkXwehTfb/wLIGtyhULTP5bjk
zp3F8SMmIucqave/aIe/Pnu29EZsA9WGMyjzTi6s9a/kI7rGjPkd+YISx1F1dTrKwIwOGPYF8kbN
agz2nWkoNDrvDBNQ+Csady8R1vwoidaUQT2M1zfShiKkoI2QTVfCvOB2LbQgvf42dugrlxtGsGJI
TjmEVjrRXGN2za0ie8GTfkaCtYkDus8X/TFmxLzVfmLUxYsuItFIlm0y7j2dAtex7W84dVTrZVHe
JnM0eaytH0e+lxzxxZNt4LSI1J6OYcvnR6FXvF4oY5Wfik4CtASRXSaLyI0emeHTagVvGzUL05rO
laXbxbkgaCJXktwh9+QGLt321EK6IzQvuHzSLHReYyD0u4oWWFbFeGB+w4+Db785N8M0LCtRNq/6
wUrKb2J300zVL8xjEszCpZ+cJAwzFSTZdhJwRja/OqkpVu4azdaonZI2riCTVM0DYKFkhLuppiyf
oAtXdyADsCDSKuuicO9NlsPjXAhUfXjLHseZjHzblr3LO0rfzfjjtihKry2hLO/zojLQexwZelZB
M236Q8JgIT+eK+zrbtAm3p8DpDOg6dhTrj8sa3sk0tJeKVcWjKz69+i0u3AK9wnCJ9wBgrNGEP9B
rEwBBYeecGo12TuVwtcPfKrUw8Cn9awf/6i6QPslK7wdmLC2xLPhz7zWU7SLQf5vTLihlE1Jws0i
m6ssnQVKGzQ6Jn+qsUEEvkAJSL6pj9iexqGITSXHZtxQYuvnovQucirdiuqG6NNIBaJD0xOksRJA
cctBM8FOla7KmykAgIS2gjiO9NGZ2bvHrM1VLfqqRpF7tGEj3oJXSIJdPzAtL1nTeymJKHuOfKGF
RcJxjq7qZOplDqKUYBL+UE/L3SlJUfs16WpRe0EoCIJbM304fQP/mXkUm4hvB/C/RoaHMDPXRAGS
shpcg9rGRXFCa2EtxCvKJ1Gc6fVjLK7Oocv31dVKiU3v2jpmghqK5hSrT4qKVLbxGc9jP97ejMxz
HTc/4mYqnWxYSrAeDtdEagBFmqpah3nChh4YbqfJ8ccT4bBXaDfZ/HdZ/oGtT76SGcs9YiArCDqQ
J3PI22t7Mujzk9NVwcNKskE92T9lFgPbvuzOHLt3YSE4jjN0JyeE5v9U9FodN+5vWJyF6VbzDO6Z
vUDvYFFG5ZPUEwc45iOhsOxnphIQtgBJacpMPKuwkMh+RR1Q+EaqZDcTZRtqEW3tktp4+Sp8xu8A
iavME9HkKGdySyKCA3cSn78eFrvZxrj0dAQAaHSeiNvxBpzes/Q4VI8UkpZUJaN6lTZmVyKvvSDH
OQHuKKmsXwtUfLprmXEmkI4ChxEDGggyh322THQMb7CXDLaZeWTZFCVZGlotjXU2WBudAUA+aav0
9+mJ8pdSxpnwH/IW1wVjbb+GZ+SXvr2WnlIFrs5zKlP1qUpyxFDHzT8Hbr/9jRIfq5AYCZbqsu7I
zAVnrboTC4EjLgETTjCdpltbYZkBAPGJ8LQ1A9pmyt+4AGWPGLQokyUDUB/SLDUFyo2XHgpwemIF
YFiLuCQ+aw3EuE7Kd+P2z1u/8Ag/fM8tm+Hi9vq+61P6c9dJbMjY1eVjQcrFiyhGwRMXw9F+wh2Q
Qj59aiwsNRw/hzLrObWlzSKupc9MQGow0IJoO8ZkNtjg1TSS6iKl5EhMmkqzX/RkA5TWeWNMCMz/
URJlNPzV92dCdC2qRR5FXTuybp+OGO9MYBazLuFmlEsM7lZ8wx1wuzg4ipLMjikfVQZbOjKEEWLo
9tpJQU44GsMSUdmxfsCoCQSN3uKdzPqPJUHP1d3rf5fEQgmpMfDD5KlAYhQujjkBLfCBEApVSWQu
KQ+ISlNdrGP1qAVRn67lPlKdPUJvGT/GCa/WcnqtIBneg4JRw5AB8C1HV7bPnTLoYLKjDwZzEgCv
kNEjHza2LXXYfuCtEYubPPnsXsCpsxZPE1WXEUZ8iDl7xy0kUhD8+XUHa3XGBz6OJ5bah0aZO/6n
Jq1JSo/WIygHQKJHrIbPlCcJRR///Czx6InpkpkFQbYmmC7u0QTJCgAUMqHBQ3a0YHqmYbvtI/db
dO/xAuJgCD33USJnctSaZ5YexJQfJ2f/jH4nmaqbaMnjdRCVMbpytlHyDRYlCtNvtFonGTYKuf3N
rgBThXeS6OIII2J/eB5syFziKfvdMYp+4wnU8H92JJ6iwKMmBTRU2GIjXPNsyzopajXBwoC/BJsW
qYNUTLNjLNiALaswwpzGbaKbGYgVxyUFukstJWE00ZYpBQIcRrtruDhrAt/XotUVDlbH7/nNIJxd
DbXf9gTpkXurc8tec066LdR7Q5TknngcB54UomIRrXe2a0nbpZZPPbu4H/4Rl1DnKMn8VTO4PNjj
/4yaXD2mIaGJyaoTYc1QN0bbBBcjtR1FOtz/Areu61aTSwFdH9HQ0GFXI5ofEFBKmW75zKzJWxvG
XErCA00hFxiUH/aUhzXq3/9NKtSiBwhy2heZEun7HDXT2XJsu1EbQPTeP6cSMxOm87fXEMJ+YO9w
RdAT9g7NMF7h2CO6/Y0KF2QyHtY4jNgAzLmZUr7C815udquJbZh6o4GAbU5ld8U3PiGasEZ6t84X
loFWBJ5ZC5psI0Yk0UTt/k2pSdtmSFnv9CgGYULrh96RRmMBc//HNR9Pp4i6s3PZYGOL72r39shg
8HTvwndBYfEGetFy8Lik8I1nO9pOd9fzPjkyxNkLFfc9rsn1jRbWbeNkOKN+4N+DozBRsoh/YAtX
s/NDAuQSuxb3wqMsb4LrB1TAT0yQRw1VTAIVAMFTIqj/pplfzI4I0NK+R2OKEimQDrUHIHYuWgJH
wRClHgriovmwdDeZNEqW7mt9sLQpZn8I8w4sxrfU+gtsDqRi6gULjFBGyxua/77RmWxlz+Z6ht8R
B/l0fSLMaITkm4zEgjgRb0ROJ5CqZ8kmgOa3hJfWFxYmrzrk5iq/pULCxE1n0d42xr0OwrR5I0Oj
COAJEX3NqEDRXeqSqCleDeaWhEXfoOomsmuKopGKjip9S1shjz97Trq5hlBpC4c9mB5K9wVFJY4l
LiRsOdMvQS764hYaM0+6eNjQpYLXSo+YiybSn5KSCO5nKK+YzenzQXYKmLKeEgYP9iv4U8GXeq/f
/3+c83UKvyfs0HI7H6ZCL2iTlycSUL+CE63c/2LTK0wzAYI18V1JNc7sxgRUw8NxL4mz0rjQ2yDO
Cakv1hzyLDKSleNoupZn0hY0retzYgfzcVSpV6AmIQmuuqN8IAogATWHDaY//SZvmMx7P4tvgVj0
/0+zLA+viKtqOlaQDgzN8lwyIZ7OHggAfPl7VSXB/Hu4o+QVsvt/q+7NaDodOozC/Kr874hv5G/m
lqpHTcbPZDA8xzMNjfxnjSQ5HW61eIs2NDL1ibRlrRoClfiNzqb/+YwiojiHXK+be0Mq+hRR7rZ1
VfehCmP9bR/xKBVh9vJZCgma9Nto6esy4JQjELw0V7L9/vAYejqLAs7aczp/EILQHR0+5Cs8TMb8
T9OnEjKjcaY6gJT6PiRCpTvoxYlBcB0eH8nCsIFWq0uzWfra5W/XYXX5/XXkztZyDUUdj6HMaD10
Q24TIKO7hobKQdTQ+hh2bju2PBcXlw9evQ2Mo8gHnbaIf0J6ZTH6ZtQr7FCTe4E1c9Cvd9R3O9Ie
KTEQbwA115BtcoQHI24m+lpBIwkIXRcevO2U+f5fKVTjpqL3LKUDU7Dt88gV95pbaExtxn8mc0lR
EEDbx66zEteTJG0OlgnyjcjHvVkSo72dg9Y/P090FM8UiNgy3qTfHKw5pQyfD7uh+FViJGUEHEu7
9OdGnaZzUV7gl1S4pZuGjbHx64OBV+0XqlNV/GVlQPeCogRXJWPmJbqN8ToRr4RgnLxTTWFApgEo
zXkShIq3HHo2GH8VVn6tp/6ZWEeG6OdVgvcqqwzf0EOAencmN2I2hEHI73JVzXE266uEaInmdthH
/BhOYmqFTmbKv1GXMm7x5Ke9aCmXsMMS16N4aGkSu9YeEtVNB7m5Cj08/9D1qz7ruaCuURpqlyDe
oqDLcLz45lUrZudcrAtBsBSrzzrmH+uU35/zalB4f3qbnNcmYbrna73tbgwvA6fcHH0tIDkuO+mO
XcgGcat0j2GBWhvjUZBZZtoVWVAfHK+IBAVv5hvh0Ar4rLp9wwOUcmu6MWsqDdFFePMzvGWkzGov
qrJa1qjYNBGTTvFZPApegE6GcO8cyn/jgkZ8R1ZhfZ529urKuvRfQMgHE6TymS/6cCoEdNtUb8fG
8zitU489Eidxwj5hewN7TYbfvuDSNYNnbgaSwq9KGZp+FscaOiNWQa9FIwIEvlSLHU3FGeO5r2Hr
+ofLl2FHHNwoNrPavx4WHj54mTsxT/vUTEfSr+RzlsOEU1tDuPKM1HBfnTe4+6gFQdIK5FPv2feP
KY3dDp8MSHvRuIOvsLYNQY7IckPY7a1hFus46Awo/Y1qtoCV7spOH/yUmbNA8xQZRvIm97NVvbkv
bObyDt2OSXEFoKhNkzliw+y9hPYMfY6JvpeKIn7/J4CdXwLe1YfRO6UKZq5ejMTm8mXhqMFIDCfT
Qjs3IBQ9RCIpj602FNfYV+ibj0Xhbq4UOzl2UdaJphnZKPixP0zbYAY7ExwvdGXWqgJNW6P5f3ey
XGdFmVb57inJxEpuTG2bqTHWbK/KQ9WnitmzMIe3A/pTX5V+HOXUt4c30glg3hSIsbRC6NWbecPk
NlfcGUypL00+sSYZ4G6AzsoKTSwPxg/enhORCWsED9Fm8E1WtldWg2MrptBLq2qkyov84tKDAbmE
GY5qJvRce5ZMbc9xUG8LsvSvt6kgdu8frDj5lXX/stGPdFJwUcFaMWML2J+RUUTiLKkj68J05Blf
WZhaVLaax3kCjkczvwgf5OSwH75K5/w8d6B49UqnZgaLRwTRqnc9q8tZ6g5onB3naRjWsyQ8/Vzr
AY6Wvoc6O37Vq97L8kwm+VBDhRsK7rg2fq3okxkofb1UT8n5K72DzVfIUDST87Uzqp6cJW+WV9KO
YgmhGNVwn8JXkrx5Fweu420PNiccVtB+61a6oTmlbYdlklzpJX/2nslY1GLS5pccElCH8TGkPoBj
5uy6Vod/OFH/4WqgcJsl+v3kiVpPeUL0TyTuCZxwLEQet/U2p1iPCp5yPFVqVOTihxM1Dq2k4JNR
yWtlLeWA+kzyUh6m39U6mVbTpsZC20gwo/m/F3E4UNeajxK9JJlhQNwpK9I2goAFS1ZppL+jSM//
iRvilxomGK7GmX2lDjMnPX2KSaMQa7r7vQoMiVnl3dAB8q9ky1YlKqk/Y1h3LZzdZXYUXj82vMGl
a0EgU4E/Q5SqEjzc1WgyHxiO1t+u3hI+3VZFNcKH0Sp2AvhadrbDLN0ch3ijCWfxEv5zrhepDuWU
kZ8q3q2YHLRWKlvM0GJDU0gGf6jyBWIdPRnAWGyAp5yh1Ive8XqHiZHeilNGoBWZ48Z+DK6HqOJS
HBAGVVf1Bz2UY23oLqDxL/QGIDSzr/kvs9++BFsEMqDoosEFLigo77+w5YkhpQc65MkaYseVZ+Rg
gnxKUv/BIeWuzigK07ifH+1B7mksq+RG3FWIIc4OEcsG++P/idW6mIZs+5ZH7hVAXmduTQFy3Sc0
fVP/eOE6uW9twzrIdHner2ULgZduqy81rUlOt5ZMVrBC4ie8qJhSwgxV23dQcDiKSodirNdQhvAx
+GOcc8EJ5fm1qvN6ii2waIzCgjIfENVHGl2qfZTqDlFjEjLsoyYworX2zl42H9oO2BJZ3u6PYOst
aUiRU4SwEB43B8eE22tAf/IVMWU6MuQl1S7qpvzxUSlH8sIEA70mQwgtqYv+d6fbYELTJSxCrLYp
PCb2uTd5PJHW7YZsga6UK8qW4QjkMzt7dZMukvnatiXzEm3RUgwKeznH268cJQ77TBXnztx0i8tx
SakSgBD8ss2mln1KRcgL8h20zEJVcS1DCA115FHYV4+0P3RKli50HtWkXL1xjG53SynEUYl6AKTA
oQewquPGhQ5FKMVqh3iFt11x2LErkAlIf9LT/cYb+cNXKPUFKLh2SHhDroQZiC6zAl5yOrJ1hJkL
6x9AIRvB3SmCJ/cI8qBJOoT4fwYpxbmz2zA452Mqxi8pFXzRgWlaqDH7wqydd3aAUYncDwm+X5kg
MMlsbovwFEO7rHL5WEotBbS3c34ESvYEfxKqaNGlflgu8w+JltnJVOiqv6V/uYk+gsBjntBKUWg3
kXlewUbDk1sxOK4sEAM4ZhRLGbKpgXRh0lwLyqjoig57MxiihiW2hS6VKllGjjbceBh3MXiTAWA7
JraQWW4YvkMUPJyudTWr4ePTtcTiFysoLOw4cpfyJhR2xuM+L2BRhXd04v/mcAXwCx0CfuPylcfl
P+PWSnQTbXrYDgNXptXpiMmC8yOmF770Dn2wQ45US493LT7OM8GHEJMEyBlLO8SGeRlnoMUqt+rY
gdQhNnI9rD21RTBJFTDDDyxACI8CfXxi5b/Myqu7yjRdG+/25l5Iu28D0bT+jAzFkeuYy83tnIHS
HqpuM5g3XoWdS75AiFpgdPBN3Sq/lOUXrhEnSsAwq5fMGZIbKQ0Xq7CEbhPGe1rZz9SGPnZx00LU
F+5QmJuqwRftaLt/Wh0hpvmt/vbUzLhJ8lZ4/3GpbW6DuHGiEwOTrdQ+0V4AE+obkxyniILoxe+4
FkJECHfbrRmfDudwXaSPhQSrXOpewQosZZPISTxBdgCpEF64793zUhoi2adPmTyHLyUoo5V3KLrM
pUOo4BKI7yVlTWvzrWPgEG0diPlQJw+OilnpJlNnVVfv4Wcso4fSnhizN5uEx2kh6l9AxpDkPOYF
HDJMKSFc+xxhd/16lGT8FfIcC7qq+ZpiFSnghXwEvDAtbgWeeoS4gkBWPdS3uI+JVrmr3GG5AwyT
nAQ5MZLaxJHqjenb/fxz/dyM4cuLa/v8Okmv7AuNCGt4EEtY5HuDZ/iG7of9WBzgtTsVOjaqYaxe
jpmaJq9BpMMB2DEo20xpcq31aHwFTF+T89v9qCs3tjeZKUXzEVyDhQn4lBW4K+xa36P0QtkcE11R
9+/UEemQ8SO3hsrbXH3pC1uzpLMIyYeS902ZAJ4Umw62RYT5Z+14R4wyd9/NCe6RdrL0I8zWT/gD
Oq/8hmBA8XBOWfIg7RQ0rnqeOBVQCEXti0OPi7FcxNtt6ZQgrj0Q9IQei2R80znDJFfpU2JwJWXs
3zxx7z4cRjmSjw1FOPtcX68kzLsq/BoseFsJ4c6+eqhft3FBdUsSb6FBJAlg2SM1BlRZvdaBQdGc
LVzr4oAK3Rza/x02J8JXxv1FrF8DNO62Ck6aF5do9mRF8cqma7dmKUpN8kyDHIea5n4fcGwwXqnT
pecDQto73cHmpCEeEnVLeW2lc3RGzUW6bhh9zfs+oShRtNmPAnjnr2QkxvI3hmwABg6jnIJNEUr9
ie7qiB59FEJKMr5Z/Fti8chEVyole7TVEqvmEN/7jNt2YpaEzk5LKqYUPgxWRQnhMMv+j5H2hCGi
ncvc/HYFrwdeg3rhESzDZeUSLDW6OdZGCvMv3VMm1kzMxrodLpoOVsflmYmhWTPPYvIH4S+3ke0R
9q6/LICiV+Ri11wa0KQ4SvWbkI0OxwW62bXkbwSQ6LCKyQWdnpx97+Kc695OcJ/QpD0iGgH74qtG
0VstueAOa5MXOIP1sTxmenEyxsTVDccJwAQ51ofqgNz8JmOl6WDMk71J2D11ZvsB1AhcF2AgJ/cX
UyAAQdpRISXxZTqI59KBTG4IOp+cHtgvcar9Q3UYdLLJ0GzWLDdjL9Q92xo/dXg90jL6BB/B58jF
4KlX87LdwrpRIxA/zDrRQ3xi5P3fut+QCCqlPhnIZo/NNeMihvZBUY3NiZZHgWz/wqwdBIPiE1XO
mGfs/JrU/Qb0ayvZV7Ev0DJRi9bwo1a1pG6pcp15JIc25f4yxBYkgPiaSJNHIE3bJ2lwkPZQZzfk
PtfNZV+YVL5IXW0umC5/Bpb3BJU3nWfYdYMw+nqS/q7ez02r8w3pjyinG0241vpmr8VbgK9jCgNc
1CWCGyB8V8MNJQhhob3Mb4K+wWsvZXrZ7U4YFdGip5n5WL0Yx/Wv8aEE0S8Kxs1oO4zIBzXmDzt+
NQqkm//q6OWdbPlU6nuA5AM1xT2x9VRISVXVcZsDhzN6FJXXyA9AIdamqmzsDXQt11uLpMGq37ln
Hfr2oE1/99lnQlRR+Yuf9IXvsUNszgVS00tUyqAyy4MeijHLHazEjZElUDsmJfWNOMce4X58I59N
eSxjwvbtg9wVRpHk8SCQL8c4oPq7S/H2r2qojsq11ARJDxzV4VHJI3sJj7IiA7HuwUjti3lnLJxU
Gegjk8buzoxVeQ4ZUPjKKUJAPkjrTtUS7iWnPNS68bR0WHG4ktsJA337BL3xhyDf/gtcqoiDquNW
YMPpJKgza07ktC7Dj0V4zW8sLzi/udgLL61w/NThoWd9O5NnWh5MovG/wTo463e1qJGs6YSqtWrs
mnF4bajTjVhC5qcoOLLPDwzSyoedrQsc1wVFOgf54VjMy8p/hDXilcuAsshJtwBJg+n8BFvHcghS
bli2fUDZoObj8mF47z0CFjuVuF1DZY/V4nQgYm7qgZIMd2KPsTvP6ElBJv8Xh3QNVSD7Tjos+yaI
XyzdzcQyTNQeJOInO22P5VxCKtb9/ukqVM9lfuAmd+KXFaPIdagK+Xs/PaGDaCyhIMIUPkNqcYbf
jcjz6XswJiV3SCxI1UaTWkRRUFeJWq0mJde8Ww11g/J0Z2aU5z4Yvcv1zjXodNc0X3T4Zyrg6lnm
coKJKatD8LTgy+OSp0l9q5fyqYqJkVmzyh1XMP2aCopJ7cymue8FdYvuirfrbmsFinoLeMwyGZxd
YCpw5J+RJgpvGQB4c5kmlNULZzCnjPq/y52NjtVFoWV51pUQ+yvkPYuVlSTO+fCToFGfdAHj1N8T
gWUYPRGJ9Uf3N5+2sBBrv6sCwzQ75c5aks/xgKrdmnKgDJV+lgOUtj3YkzCagSLMdit1KOEO+eUR
2U+qULBert1Be/aJD5W3hbhpqAO2pIhXC3D9cQMyYuwW4bJBbXuP+3NBMTw1Gf2a5LePMRRQrRKu
4ZScV6TLGizxxnJqFSub/CSSUF2M7wIGrTc6JnjhpOysy+wW9VdnqgOS6dARQ7w7hdZug6YuUWD2
+2sjiTKVb9Q7/O2FACXnj6R27mFqO5iSewWVRedDlj6Y0pG0x1ErzVKXfpzGx+jqr8IWZgWIJIPG
ZtzwbhRiLdhJB/6UEv5WYzOCx5hr+oUsciofnGQ8sQCaSl0q8oDboxzyGgEk0rh+ffkD3TU8jx2t
HB480b8n786TvQhKkCgt/D9TKEPqMCsKDKb/foUrHhRKSEa1KMyTaF01PWHBSbtqR05L9IzmdA2c
WyNqIA8mxvTLLfBGDry5HZs3skeTtA4h1yL4FahWIjhj5PmLB2uIzG6Tfdbq6wJNsqnDic8BwgVH
KjmbMSNo1ssrVY4aa90WNP6yPLpn1JuXijSVyrM/cu3keWaHNV0IV9fQMFiYNWs4h/NGS/iP6rxi
WZHHjG5UUtcn9dOdFnbSBfs11w+DG0MZpkPDkEyQPA0zA3YkdyLm0fvWUk85r6COBIyFkPD2dszE
PJgv8CtSVsdaPMMLu69ch0xa+uP3BvzpKpQ4qw90feX2q8LmrZ8N88dsWc6qdR5YJYdfkpB8jzmP
fz9iej7mkx86r0ACN/Q0UrYfTM9c5tgTlHCRdyIhiJUSaryPyZ86Jq1fYkLCcx4BmdAHB1bPW0+d
46tE2pvcDe/em3IJ146VyfUSFvDBnrj3ejVTtmos4FqX8YtS/KHWNsEteEJMSffZWg0UQ+e4s4cI
/5fhvVkz4CjP4+XO6D8OOMsYmxNRm7fozPOX43HpoBpqSx+tRQEuKV9xRwUYVy22w3o87zfP5a02
093cxmeRgdDezza+4wLQnLFH2ysDTtwTdbz8FZI7Xe4+OlZ+kbGMbbtMErXDYQvECSL+gxGOy2A1
cPLKV7A/1T4BcljWzfiDD8doKz9G1g8qZjF1AlfTNa8zPe1YAUjE00ZAjlo77pS9jPIWQAjwvDCT
dSvf7XcDjKNrb52JHRC2Z27hGXoS6nK7mLu8h9oS0aCU6API7Xclj4osps8MBCH8+oG1+R4xbzbC
y5u+ep3a80EgYOaiZ7T2EBMbFEqn3uL9zp80RmV5jUVMHDgFXosBXokJlxh8c5YGqXDLToe2tfC7
5JvE8mCKm1+b37dFojTU39ZIqQiUGSrMxBq/V6h3VMN7Kg8LsXOg2GU6nACLfNm6w2DiurGoLEFz
BPlJQZD494JXEUpnRr3hxyihj+BLahQwYBGvMx87Efc02/uULyzOmCOLgUb/iZDas5vSA+mn3mQ+
p+XOp7qV/DRBTezilIHhpcn/PuDnn6nL3x+ehRY9Imd6XE+Q5O2ULV7bzx8Yxy3aMqAaTjKE4XAr
QSgaLFl5qpYtDzPyR67872yTn5NSx9OJCpHadWlI9SUsC7lFRWVbex2knW1KbbQZhKyToX8NULJC
Rwut+oLVBe9znQFv2Uq67UM4jHgZBBXCGqvS205IkNsrf3E3BdivM6RNGw/elh3GJSafIp3l6Z70
QIn6iPK0//07IdXcqFxtRpmNeieVmCM0ZfVqhYfgwYjwruyjhonmCUqI3RunFpEp/8ADxTly+rcm
zBTfljo9PmtfbmszknkL0nQN0RRddXrlzTe6Qn0C1oziglEnuZtmxGmY7sNmPEvFgYx4liop1rli
nA/8iX3AlY0MvNXYnT4DBrKQ91Je4Cp0tkMCpXXLmcZByN/qkvO99uNpQAxG4tj4DTXlhlrbM4hf
ssVPmFqaDFYQKE/CXS/XHzX2ykt4Bxt++QTxUZlxVJkTR0yATZ0tgsur0VPmmh+6EqpflWQeNggo
xdmzZ9OwH6Aqj0YwV6iaGVkLhrZv9tHozM1YEBY58uRafMhlab9RzNcz8SHUIOeBrkgFcCt3lwFi
OJPSEWOkMAEMxNxUWVNhX8f0vGgSVo28l72A38R//9t3qKJUngHqFqHicINvulXI9PxQQdhj93wD
G54+/1IcRyOu+rtMsMnNgCuiTsXDkd+6P+JmOYjWbIC5CIAF5qwJ1qCafHyYY2vw2uMYF8h+yhLY
52aWl6+ziMt9K+2uxXn2jgse5tgBt113UZcj5gQoFtK1dsUo6g6//t+9aS4x1VwqBEHLzBnNrOSl
XjiyLcCMs7WEMPTCwRWXsIx68axibeRRkGs+iLjp1k1Old+IgnmZALoA1TlRVnWCrDxLMeScwxE/
it7b1tGKsGeqJNUnDqqpv8auaZS6pO4WEtEphSpQZ8+jnWRutnlJ8lia8TFDTHz2BTXwGZxtukl2
7vwWjfSWQq/1oXIyldM0EXQVvE7J2LrjY/yxRdaqE0NB9JsaOlJTHAWwU17AJcuLRM+fP1G4qYjs
Jc5Cap0T79qEJ+J7u7FnpVl5/SHdR8xW+hDVaMEei5s1gW7AAtxMvEFe4LZzrau7e0lm/b2R11Y6
z7WiD0YXEApmsXwI117z/0FUkWersZe7O0jL5IiWroJqOQ2G+b7Y29ZUL0WDtTnyGuXsfRa9maMU
aBaUZy5+cHVeg158DvwTVFissN9+70Q/1/SXcXX9gfbhFiuH6vgYnTaRzcxrK9OryEOr3Mkbe/pZ
Z808l6U3menF73BJ0GlaYnMSoa9GMH3Z3c99HDZbWeiQB2EY201p4OoVTxJavS6JgAzsQqdzScpF
Dv0HEDUfVJgj3d3Gr/4kFin1tOsIniQvMuDIDDG4YnspBuvspGyXIApUNfvOz9p1g8eqLCqANAMf
Ewh1riNNuzRgYswHkhYHzEnBzl2AvrCxJpXwcVl+DEwkDrcwmxd5WDls0RVeLsTUCNaYuoSZonk2
6xLS6gxKdRrqsaSMSQbP0zLQk2JC0UX2euPgOK5jHu7yUxM8meHkmD6yPtzdb6fnirzArW9JQokL
xzpaF+c+IgGsHb0G7fNb5E6mLh774CEQySapZ4GZBJ6QURHRt7z3NX25R0alOU2xwRRizooMN6nA
Yd12wFw4nm4y2KmQuqC0ztjibOzdtfowwH9Gpw7qSrEJmLHEBbZUbfOh+8+4F/sgVe2e2ShaEchw
SxRwZBLsxtaTAgydf91gZvqU2RTRuYjeW743dF6ncwR14ftyQugYysmsdp8OiHk/PRZUvVo7RLb6
P0iSTk0YQR3T09UcqqDYtcrEp6LLdSXp2YlveuT3qXlFbFdm934T4vZJr4wprr91YKdI5xLHluTN
4Ib/uxBj4JITmDXM4g+jxcb3j0MvgJJA8NYp/v+mTk69lgYOuJaAit2IVhWobi2485nJRTXSQPy1
3QDztghy7Ub+l9+jjR1BPKAt83ANLYI0hDJGM9GReda3dfd1Z0jQBVu2m563kYIwNeNuWyD2OdVm
oRh3WjEq4FR+MrNjfYwOvq5yi6Akfwbg5rYw2lBzQ62njHRCYnexUlU3ZdAs9iOMVymIY8F7MgwA
USnL1HPy9pr0n9fMBF08/nMdQgWEkYMKPwSQbqERorVbIOmbnEOKL7ZlrC8qw8E8PzmifGGr1Lcy
kFU75gPvompEXS35j0/ORuUoxWoFrB+NTdb0siI8ldBYgaqOTc9dA2IswS/Ak7e5o2lVl1GKx00K
TmFPic1nwNbuBwlw1mxKDhNwv5Z4qFSHxl5UhElTEBwt/RJlXd3FBDcbcwR220AM7EwnpMkpUO11
Z7UDtqcYSiI3c3L1i8JpjiRLFAtRpNu/zF5S4/ejF6rN0P9F6Y4iF3WlXXe60+pDdMg7zXJ6Gr84
UQqL6mW6hd7mmAsYPNBrqvIacIwWWAzVpjbxcD/CI2tM2A2Sj5edYVyshgoldwjJdNHtlNbSWpnF
dosiUAAU7VkwAgUtYQE/5eHayFF2LtT12DnrTyZgw2q2oSrrwYxscosGjUssDjcsIN9Ngb6ghiS/
zfQeUbKxDtfNsT5oQDcAgBdRWHjZd3yNYxhAQ+drb1cugVqoCIBbEiGEgyaud5qKeJrD4IksdeIa
lHd2yEO0IK+RLb1jU9SdZ7hSFg33kGtORM9EK09t+6yOsgIFfZKiaIA6cwRZuEJvbKz2YbS85Spl
KtnLAuKWOQecGlsYTvxQETj2sC7fIB1mFw3aPXhqIfDZUWGBYMxIb4VM8pyFzHl/dDM836fstW8W
x9zkbaTsXyXaCBdcjd94Mrw7wO+qlhYe65S+qIne423Yz/rJMN8WIKiTd/CbQJb4CAa+Q//uVD26
tfgZ401YEGIS7+yOAnIu3lGZHqDuU7wFCw7UD04Ux3WsL6o6X35XibFpK5OBPY68zzY2d7kAWEL9
kERWy0ILHwPVfaJYIrPJhIfFCKA9XoUpxbaSTfqZQ2nw4m4RVDvzHKLv53SgninDV7bCB25op+89
V4zL/+8uLCg0Oz00D1jHRkL8PR66mj+sYnmKWqUrc7m4UOJIOMhYIn0vswwVojWZ4QoGI++bwcY8
jtpCj8u1p4XH9/Ic62EWkGGmM0EdKvMySADd7ftfqH6Jc0KivBDBjs4yjSzLhfSH4f/CVVgNqInu
IN0GabE0GWFD03q+guvaEZJXegFv092Cnff1lDuZxLNoNSRmgfizwFA2mnL45M3P0tzRb9NLUR9w
PRlCjbzTyqcl2VqtQ6Gr1yx1d4/cPPHvNFifBq3wkpuxUwqlnHZWVnwGIVb90+KfFHzK0pg9mYnY
04nyJFiEmzbkIkeTKs2ufyxIRWR0nu4xoDyTX4Jn1gVM7Kfoy9xAsTn37VZOjdEGecfP+oV2WEe5
eISK1/0ab1Pi7EtagY8UoEMSMJQOoSwpvwhwy9Zmxd3ZPX0krd9G8udpdCjPnnB6UBWslajixXJf
gIj9frZutCYKYOE54lXzdPq59jmNbBEjSnnNhibbgrqVdWlsintZ0EqOm2Rv/9pv+2a7gP/GeS3Z
/8SPG/0XAnjikgmglIj0B/CWqlD9xHZu1ALI1tq6XtBCEO0jpqppUvcgRYVZpL1dbQ47DSRVvqJq
x4QoSKpF37i2hzEnfkoi0fo7oJCFJrmR6s+NsWPmFIlP7u4W8wx21Z6JackCoTg7JeFnpYokWj82
0i0u+UG2Ir7Uu6bojIetoUxAvkyEZVwS3iCn9SO/1tIIxVJrIsog4j8MqwbnQ+lBOALklhVw0ofA
+/0QtritOmep1I3nb0TqeR1gIkhP6Z5C29fIhBrk9hY+G64grQ2KOQU/VvzK2bxgmvW6TNDqM+im
qauvmDxEkR355gpRM6E9wak1WQ2PVxYfJMozFghLVsLvozA4JEc24rdZ//IYqovxr0F53rhtJXyV
00Jefu36nxjsZqn0Aoy9ysYHGrKKmbvfRSj40twlxAod1ar3v3L2C1nVhWIhSOWtaXU8Zux/gnCO
HiHQrBOHqGUhCchzZaMBSXTcjZOz+EaTeiqTa3vK/kbsPuE8z5CUmI9kIPgXdjXio/a3gAGfxymF
8dVPS7gN+2bmxZiFqMpBmTY+dw+xZMa9DcqCw3lRoGv4SaNGE+VcU2oPBbz0T3D8I0mnk1dBDHu7
cEltH81Yra8CEHlQlwVBpujPPjAX6hghMbrf3Wsk7zTUbl9sWmeeiRHPvEfMVJAhkHZmqp1ancGq
ULV05G5EizhkSVuo1GkOwCjlOrBd8KoAfDUitZxqTue6DspO2Uu0tQ8qZgzeQh1cFLMNncaRb7F0
1v18YYjE81NVkYk2R1GxWSI6IyS5u1Rxpx41bA39HNrPG2WlD8b8uXl97xxq8UjAovwKLFoWcEDO
zz7nphwJY8zS4U/EYtN/yTm1I2WrcT+seDhX7aqnmgB1ZnL7U9TG6L3jEVPtCpLqCaRxsheopfqu
j9FqVg7gWx5e1FB4bl9rmRNRVVNRwY2uel9YpO+RI04fXaaL8R08BEnNd759iWPcrjknEArsvEjp
++yP1kM8L+oyqBmtlzs59ulnrQ3sJm3hjPTYs0YRSJv1T7mPXsWxA1wYkVzlAZeMWwdfjfzODJjh
9I0lAU0TqwEqa7gwmVpB7YOz7x3QZ3Cqoe+XgGoyfMuLvRDFm/2OJqzntdRoITwXQ81H6jOhKssx
3i4LARtXGfbcmqDQlGFxlVuKZberu67plkf/smEvqz6BxxsceYsVPWJjHLtsJvwP2WRShRZxIF56
PYUzAOBP/rlEpEsqVDQHhICl0rAQuJEj7LDigFb+zPJBLf6NSubPzGKmYoHt9xYmwSPH2TmlBaWJ
nZPYW2SCG2YJ966nXqUBG7KaKNhZF44qZo5JDryGf7OqL1cGiEnJx1WSSltGOSqGFnoHdFcfuYbz
X6NPgngYphG7UJEd5/f1Z2tjkcei0Ix7ouviNjlgNTm1qzWS37NSteev9E0lU+OLfESFBE2UK0eO
XplgkzJ2PHrcnJ9t8gVokF7QlSG2LhvoiFbItOL+aAKktRuc6u7jjfC40UO6TSYK+oiHgnQsdrbl
s4eTs41ibsYP35cY07EwHu6b6us0fctFFzNiWHo23ncE2wSro7zIPSugs8Jj6hH53rAGPGS8z1Ok
imxA7fR55BrzD5oLEcX7sPAaPrg0PrbMjmb/E4QRktAh0eix25Xtc1Jb/AY8QSV9SBpOSLefNSGH
hjrf9SHW3OEr/jJgaI3Yuq4/0CLQG4YKSSQ7qRNwfe6psbwoXsP+K2fjwPU/nKF5Euy0chP+bK/I
oEJfKm97Y7kGrco42s4FBs2r7BGztgZDdYkEAuaHcpg4rcyU8/CMbCPtBCD0hQc4t+yRGf2O0ak1
Fb6gRJ1OM6fVbAB8v/eGWg8IX1XZGEvCfKQKBOI86D5Uuv7IovOqksC863iW4qPCVpUM0onWZH12
38L5OiXnq9Ce0A3VwCSuEIRPQ2pIslp7XZyCHkbl02JQ4fV9RMQFeDmelkuPZP3+njAcQcZwQKIw
OgQie5HyNulcynmFgCQyyyeTEPn0OPNK+C84zpOIq+zAXlW15t0iM8JIW00IRnX6mcxDyjO1wkkW
JpGQhBY8Zz+OSanYxJQUbTg1nGTOTGXRDs1gsrtafiDgTpbV94AjDUIiqg6r6XLdSpQCQ+6bGQxr
2S6u0Ee30/txJnxrGplc4mTicqmVLPOI8h4SpArP8X2BAZxWyUY4plF/08C7EDXF34+Nugmxp6hb
TclfhQyEGP+TOEaqICNh5VFItp4++/86vkw9zhRuCH9Zg91y0W7WK7tlgJ2myeYMkaAiUZtrCJt/
5b3T21qTTgfMjww39SydT6WCVvuIAOv+I70CmnDtwq0FDbNrNECdp3j6WNMFZcVHF3P3j9ZCXgzj
NHgcXi7eJmJsvx8VohDMCersVzBDY6I9RV9YKzlyBW3U2Tu+Nh3U94H+32KteADBV+aBCrB0k3Kp
F0Yhw/ukdPI0B95WhUvG+PeQ5W3e0wi1pOVwNRrm9B12OPbzbcHfTAXE+5JMIzEG+IKmgkBQu1n8
BAw0PemwubbgtL2kYkpiDCAAE44KDQXFafuHzrxnu+dqSy7lULvcyBKg98muHejp5hDKPvgCurWe
UAuZVFkY91YJylh8bc3mFS7d8JqAPsXSmH/c92NnYZ4Si/Ql1NtgTv3iQhUwd8KaTG0kJSJX+K04
02MLxPuhX46z/jEwYtitaJnA/3KLwSky0+gi9Bl77AIKSTLJlf2LVi69HrxaWE6VnNh4nqL1enxN
TKRohuitD0Hqupb7W5b0w55/xW+1sXCUFOsaiZ3pmb9eKFX24NVuD2Lh6lQVrzfEAjslJxVol2a+
rrayLKAqAgsM+SwW/qZJ4jMQrVFnu1xrTY5XecG8IEiZxpzueeAlYTr9u1YtOnXvRHjE6xJJA9rj
Plv+XDxdd1UBNjGqI58i0z4CLcdxOO7jRRrmWWO9Tkh6PLDGhgNO9/y69juKtiyf1Y193adnLtji
r0JfFwdEQk/uj/7MbzaKEeozNUVJZIfT5/wBykQ4ysaMym4vQvyaAFyb4GTy9HWkHv0yalM8+oTw
Bb3PJfKSUKDgTcLXmEqiOaOco4qmEZ5Mi+K1Uj4+dm/wn7loRG3pACgQpXImiTEq/bW4RM4pl6C4
Lsnhssd2yl1xEp3AQP5yRrEB/qfa3KXTk/4RHcfxH6MuCcMpa6uvB/rMK9unisrbEOq6iIoHPclQ
q2oM791kbEh+xxKtFYaaWifsCiufPQOm52/O9vWBmhJXUKBm8hwfOjdSVQLPdDZAZ+JgcfhwtNhP
RQWAA2N2KwYDZWcG2cz8ZIwF6BV1LO1qiqSMtuxPxvkNrgTPrP0XVLuAThUfCCOa00RAP6jDBUPv
Z3GqG+UvJwhqQHVF72MAydltmpQ+Iy0lYmowWSkbrp85zykXJiKlISKY+6uddPXLhVhKge8qzqg9
6OV4wJztHyvuPWLy315nrsTJK6iKWBQo+bXniXTqLdauXI/0QSo2E1WU1uEw4ifrR/hGD5NguZ0I
Ca7DNMzEfknsky17a78X1iqxVLAjmaK9yghBiL0ybhmfZiN/3YZxKKszi4cbNBQmRSTyMSfK+Psi
EEhYZ5Y0th5S9k2NlC6yExDY87YoshDAJf9xniRnE36QIDzQeAfG4nz+HLUa2ZSw2uDx862DRU1B
sapIcjO+KADnmSWzC/l8jZ7zBu2RJZk8/mLpvKH8YyNP0pQGD94AB76oGTccAAQXpkFHOIEYLCB7
xE5nvlHF1yiN0VAjKhIQ0W9Wb3YKg7Gaj6i62SXaWxVh0gLKHaSpOj08rUQQqjDq0Wqhf9y4NMMs
V3LJUkE0IvZl8Ndv73ODXTFWWhz3y7eUpWDyKOLANmDsg6JTbnIP+UuIR/npkpZpfuPZYOuvsWUI
JKUGJR4VruoX4UaVDEWGVc4E7AEBEJxXaWuOoOjWzX88jMVsYkDsATJw7lo87iI6NfO4vcjLqkVC
pWgnAPZFagDd9CfP/d3W6UsxixTL4vGmfKHAe5Xdyi8Cdmsope6XpkAM8HIpIjU0JHf9LK8tIlDO
ts627hq9ltDZe4jlHqDosWBS9MO9quHlWmCI/fZ7Mz7QT1dzP9EkuQ/O0Sw0PxHCYXjZYnhJHKfX
OKFebboNOx+EhkLfHGErZZlxThqJP/goxSvr73N/fBSMYOnRQFjeI9Ca0MBtEZwGXJqvMrCm0oHg
gXyTCV5W0ZKkh03lRE5lyDjo4n64JS6skWT9DlhAz4Vk5cHvv8NTpKLf+gUgpd2XnX6LtG8DCLuy
yIVEpcCyLx8mKE9gKxOxTTkdbJTrfo215Pfkkion82HG98EZKvfyVtoNJy9YZk/saCF5l/RpKr9K
XqM4muxMe9iteV7Eo3IVUPKt68mllraPlCrb/I7Oi5TC3k2kYd/grNyxptMY5GZxeTTWanQUMPzy
2+6w06fX8pW/ChfFgtfBQfh1KAuVeL1Pxg8JXkWlVJSvjiyEGZbAsHtgtzpkCb6QJoG1xt+1Ly+Y
kbRtmg//x4QtyeYJQSxoE8PDWjErLv4SDvl2lHtzq7wYuaGyFt1+0+DZ3XhlDhctOcueYgUptRX4
DDQOE64iNmG3k7TwgHTewk7QmBhZCmhJeaDU3v/YhVPYyP3TdtQL8zG05W0wgqmM0n3htfMjnJds
2SaqEGLI/gWT4axEmmIeXlXLn3+iyGl5kUkADz/wMADxEXls002WDf/blvQSXKPQW5h1gL3cNIFa
ynrDEHWcPo7KIrTNv5XmQDfxiN4834p5tQV0ASN5jQXcTfIYHyVjV90/kDK50ldien9yHWbRv75I
353hrPenthFS+NPyEvcUPy4KGQ5WrZpoUJzJaDZiXXzJgCZbPkgKeUQNONfBloml+UL2N3dgYTHT
DutSRtgM5tRT8xrLBqWpuWmNB/6A6dnqDA62lWlOTqQma86oK3ISrYXB24mHi1eWeiKO9aVKPxfc
YH6iMYtvhkbjWkbvWhcazxOB+jIueEojQw8V6NrUNKc/thBLNZ75e0dscaOCO3rCbaf3VgYpK/dt
8DB9q5OafXWEUxy9EfuYg9JQQbFlSUU/popdNJaPagLY3zNM2K5aa8Sl/4iLLlWlpDLi+xBt2juB
5g6yGaR3S7i6TkMKUGugcbYcPrb9XyvrApbEtWy2T6YmLUj1RJwVLKtJsizNY3sEUh0RY8IR0cUH
BwAiJehtTiMLwatxQmghkwPWGrx4VVtPLVJfDw8P5CHN30ugecPSOls0uy4gL2BTz244tzfc6qrK
1gZiEa/7wVkz3dontxMfoRb1696rm2qv5WIjpPgwJt/EAKs2lyxGiS+6ynrOTaaAw9OIvSR0r7W0
VbX9yJXNIvjcxKXfjLM37oL8Zylx37E3xwKfLVIJcyc9l3W13QC3hOaQuObw3t/h2UKetxfG//Ju
52PKhulABGJ+C4IzoVn+rre6nAsHcYreXOk3ao2HBlxvJchvYK/Ok/b4Kwc2Vfdu/eD4xv7wQnUu
CfByoHytq43zfW9pL/FSbXgJCBVOCqT3v6DXi2N9o/nEkG5VJXQo/o6fZhfhh17QQdhYvbCaDTw2
1QAcazt32hxsCfdvjZFUe+x5sHP/ZPKNbkO/ZL/Kmr7jYX9OOVv+5+Mt2NCBH9VmWJMxtpqJ+u1G
4BlhbOTWpAU3hup+IWAJZpvVYQ3KkJTV9flSzWswdaOwMYkl7S8rBJPXA9rlisIaIY9OxIXqzUJ9
hsGY+bAnyfIiEdB6citPdYILUtZDhqUnxPCsxUbKTH6OTtE44p1FssgNiaY8/+RibSjx9GOkUx+T
19FPCs8u7PVnihZHxK2+D0Bcc4zsVC0ZS0wXBzSDeFK1GiOq9XLIHaOMYC8yI/nRk7pPhORMKZlX
oebAC8z91RQJhkuNSbXNbLgg+J1HpAuycH7czHl4OHCN3Cj/0hiWoaWUVJT4XB5OKqYIfd1Xzj3U
e2A/t9s7yT50cRtyToiUWl0k94ad6wM2PcnklPdZBoW90JVG5VcpNDADjVqHeiOEf0mrQ3wrUV8d
NIhB+2qHObw48FQMO4ZyiC9sxUtDcBbW5CwU535j0tUclDEtJ2yAdKl8VLYkvMNj4wLm1iHsB9ST
XI5rv4O08dfzgivYNE73OuM6sktEv87qC8jDffy0bFOjJJaUdapWxm/2amSZCTuDttmt0ojVXTuD
ZY7P7npt2CclHTR61sSeJghVtobobIAaicfol6Ozh+usnDzgnSI3nmMs2QrMZg8FrpajbWNtsNL2
XSrQKx89UD/lbs06itb/5iHCLQT5RTpGJqsMK0reOugE7sQqyBNht8XunWQn0upr7rRznRebP1Cd
bxZ1XT9qlfOQiZFfJsHZ7By76Fcm/yCgWvNV3Dg3Otg52ApmAHeEZl5xk93MdN8iMrL8oCvkllBf
N7G4+LvgrB8ItCesfG/JRx4JR0yfPznvEqLHVzknLJSHS3wfcJ1IIL8XxKN3gLAzIOSCqPRKJ8w3
Qo5tT47iDEbf9AocD7vWcQQ18C0MGo+y8ikVihs/ECqxJEDEsz/MBOIvHV6mk4FSn3rnR3rX8al4
Y1jGTQK/nr9NTzInZnqsNTnBQqCFEuh/CXCGcx6mG2f3SU8MW7q0Hj0xx9o/T6srI3lq7dGAz82d
uNPDNOhqbZ0WDUMLmuB8MIpCwfvK+WhtoczC09aoyBItKTNSDQ/1m9DSGq9A/lKlH144WjE0Ovrc
1ojzDc6M/N2OaMlnU4zJMethBjC9LuLVQTtvRoJ72b8lZ91fwUCT75KajUw4+NXA+f7vjk733Ld5
oD+5NpOiHnBSE9xjgLvvPx8H1/pL+w08eMGJUf75NbdAx2e4lMLw7I1ClYRgQWNvKI05tJkzpMUp
ZJYi51nXl+3IPkU+AN//8dcB1+WVup2IIbbP+Q5vqS19oNXxIWRRmejy60DeKezERorRGqeJwh1W
FqnOXICnawSvoVA0005MQIS3SuuFkEhAAwwvYdsGSEBcl9WVOc7Pvmm6Z3Ji7/lowzfiK2zMRZM2
oqucFfTEHbiu9UovF+7FGQH2vK4GFRRipsNqCSHKYYI23tBPkVZBW38Wkj+kR9VB7qkjAwIO5JcK
s2gQ5yyqSgTa6EykQMNxg8GE0zbDLCrHSl/T3iAPv5GR2OsXsgYi6oGzFGBT5YZ6axviASwJH4fr
QpnR3Kp/9PUFffXbpiMd4Ntp2Nk3L9jGQ6MtqfWdoW2SMXHtba3dhvb3qF1xQzRbCjZi/1a+Bvd8
NCmjQVFJ3/77ptScrrLjVPBhSfqe2pL1pHImSykHNsK5i6XZgpKzFojTwYjkk6qid9m5BHkQ4Lqf
c2WpJUtJgamjMcZQ2Q8uOUf4p0gz2BMpXcDiZpdtIR1wp1vFYECuhfn4lK0S8SNrhTWO1iPgp28u
3IPdUiNeYyNb0XXYO7u/UGF2vQXhbnUWy44bzMdfXcHiyM7K+CAPjY8lHZZmEuQhGc0GruXTvHbl
D77wd4K9anU0itEFCyMPpuXnsGCe08NvvS8h6guIY88oD6W9RgUxiVvTZXujfuOXbPseUuhxUiku
SMvGmj9pQk0XAxAINDb37Vm3dIcQy2KtP8lX2LaOonqADaN+G9oDUGOQC2DdUEVh9x1N/yb3xiXA
IyQNDKzBOJ0f89aOT1lAkbto8oGWsU90lYp4B64nXPbClqLAn0K8Bj9cwuGI/EJbJbzubVVmhxcD
vKqSidoums9/xlTXdTUdubbYxvQt/6XoDp35rLg0hn/sqVZXQ8X66nJC3Ocsr4eP/Jw2cfq+rltE
B4gwf6pV8P7WOu+vTJ1u5YeSWx3gD74pS8lSsvbZiLQoWen+SJQIAogFW13+eBMeBMSH0WVP23eA
FzmyUdQx1c32jpXPSTetl/gYogCqy8qqpb5g2FZcIG0jZYOGW/ZnoewBiiZoQWClM/ox5qNLpwUv
Agfg2LhoQeQ+3RH8y4VC4SK8cLLHHfnpzqXI6doebrZvSD1YhCsoYMoQD2/9v5EirjqjYkNlcLwr
Uqlq1a6CSFKpWqSGVYRY60WimAd8KeMSoyGSi2RtEFD26TfZb+26+2BiWi1w4ekca/3jn0pAzEME
YregMRg1vDJhIV8mtRMVSbIMQHYTsXaHBbqEmVona8H8R8qFsHNB+MKyshq2s7N69J1ceBMi+j2C
PslS7d5qAVdHjx/lD+TbxdE9EQAdD5sRSCXebRRqexCRGJYRm4H/KZuS3FbfQpHtSOu+Ai9OrFQq
xViDgARXBpoE5+Nj/lymmAbtdHlkjoXenlnV2mxq9UMLAtF3RyZDdr1S8sU9fWklFHLwvHy6hwTW
L9DHYuJJbSQu8nVvw9CB6zo0FE8TEjseMtDermS8nb2faNtAV9b0cJPZs5pV04xz9rRKXCcoHl/r
PY03HsyyV1OrK3cfymqZqzLIpb+uCxtLGGMVAv9zel63F3RKXXfYiEKfQHvPLf1WVVi3uhk0QCxb
n+2Q7EzCMf19SLTSp4oD3Mb7vYTj/D8ALL0BdjZRar0BOqjoEv5zTefpGP0tx6bEJ+sEouGLeCAQ
k/xLd3VJDYaEs1CUox49yOaXWPW0s4bAKfAGbCNNQcWvB33XqiRGsznOeREOy8iCm4WE+hss4lIm
K3xlCtSzYyQUttFNuoocM4wSzPl3fd3uOf7hTBbBhNSvadYxQwNtWY/UJaZ8gZGE3+EtCq0i64wL
glW71b2iYQd5+3hGgMrAn3Qpw1DvTHOMvy/bJxq9rAZGb0D55P+59UPZYq01zeUYcOAxIcVP5WS6
woFlflNaOtp2lzZvjxrlbhfQEg916iKYSk2a75Jd1SfZufmuTik13+UYEWUOXLrHHAtoyuhEwONo
/knAgNmS9rZnEkbQ3MDWfrmiy2ilOhRkVK7ePijDSQaoSqux0V8iSOJLyDL2PlW4CQFnhYVxKVaq
DdJ3sUuEeYk2iqjhXi+PJIuZu+poU6CslSrowgC6zmYuhzLdumDjCx/qQ/tw/IUmZeQGKaUlUcyU
dmdS3Cc5J8wQnE4Q3SAw7WJIUtgLpxridkIUGv7H1d1t2NNMbUprvSkKhoYutspPORgZJcDAOHew
9Mr8QQyq/SvKGdDth5WQX69dfmHXcqLsfhvNv8OVa1/jCgX4df9u84yoYxFHBf671bRKSGYQzWlw
hc4xLtXhyQETFqcYUl1q7xjFWGFhfxIpbuFTmlPZF1KKYo5e38+0s6S1Ok+LAi+KEcGH6YEyG7RR
gmaT9f0Fjslk4T5PsrNwZQMebq9Zok9Xbv4znwOJk8eBb5orsHxs0emPlBpAihxYWXGUROmAqggO
LIsuLaWBlk9fIIqf2EUzxL5ihlTQ56wcI4ljr2S0PJQu+J3aBC1y0oJoFHhfVC/keA3SEzG5j4vx
g2TMQYv/jlIzUqekyF7WN4jYgAqavCN3mxn45iIkVmRpBY1GtJGvIgtx12qFsabDLlmDrDPSmpdP
SDbqsw88ra/d0jqvF7bzwsb/gWdgCwbYaUiiw3jGmtj/MwCqqL5Zglj3zZnwOIJHr9uucmGyAiUa
XdVkwuhCibZg//w8M8LgrkvLbOpQdDsPqby4BvltqV3INmpCi9RAe/JhzhW3ahLZZ+a2M2pIMmDl
Kxdazfo66KvrwuOdrCJwutrNkxd3TnrHBtjYmOZs/k7vQglUTV3tslkSQ7KZ1zeARb6Ook/X2eGF
eTC0GiGwr5Uo3GgU7S8hlaE/5pV2+J7tVk8g12fUv9/rjfmRN88ym1Dks7DtyDpzoVnmwsPCuu/F
R+Xi7yDYSm3RTjFzWyARYJ2oOJp48oWkIL8aEavHJ3I7Br7+ahF1G1SQxr0heSST2G/Xbwmg/MA8
fY/3/Mi4Y4EjwWZQKSUDBKkQowMAgB9+TLs1aLkKTpNvj8n/GT3kN2Ff41Dh6uYfLGl7u+Oz4lxC
FZfZUq4/X1MTqqMVgiQtWa8kswVcj8dSF0lDWW2rSL9EuqHQXUrHWOa5EDOTGbgHg+e6AvJy6Aey
9oqguJ+kvUdsPB/rhd2Ru4CeTHCsptOMtSXUPk4xX5iYuzN4tHH9dU6BxxCaX8Bd9Bdhk9y5OUa6
YI6MByWJo1OVPxxDVptzFjAxvSMd8y/cnonNLAUF/44qBL6OEMtqAwcvI0Nk1OEzT7tJjgZ6J8Qj
QCCWzPjgSKHLu3Ld8ZVGZOsMzX/BZhPGRCw2cGa1EMSQBY0j96xN7n/7RxiTpSaiWOojYC/e45jH
Rs3RA1aAMTc8rGl82dm9Nba+7Y2Sp6NnWnskGDjtW47mjTlDOJBZPnLvVIeAcVEzw1eA87aVvQ8s
5001VE0CQWxDdhCQmsZeldfpshpO9ys+cffmUp0/Icdv5tCEBc255iq0vA2YOJ12w/BXr228trsY
gSQ/Lp1v5LIYoORKu9dHpL/5cAnNp0at8j8/e8QNvOvHGc0TNcd3tKvW5lqsAmOQEl7EkUZLXUmj
vGqnujMYqgR+ZftYoAnTK1HZ72ZccrTyZmWF17YKW441FHFzpki4HIUEl7ovJ4Kx8aUyT6ougvlx
vgT3wCWaIcu/+vgTLeI7SZuK2OR+yvv9JXWMhFkGCsNGQPsnlip/Nq3+NA9trF70G7Thuvl/BJv2
epG/GWnf5FgviXLrrYdXTX8mw+IQHHO+fx+VusiS5SB7ubyaGWThgrdHZpwcHYARfTt0VtejvcZU
fKV76phybPkx+tOlioGmv0NuiuP+u/zqPKGK94PaqW0fZGKznFPlFIrOMKqh039R48s4s9pTICmG
Ucx1ERwAkVX+AgvmWlpPtUfx5gUDOpQwKK4PVJfweKy3up8QODMUXyHecvmvGttV4CosF3WLWaJF
96BlTxw0HFgOGlZ6x1TY0bFOc9CU/4sWIBlx1CT5Aqw6vMtDPWoIGcnaOBzL0MHkzMYu/Q+frT4S
r/LSc8zc3jYv0moBMyMlNWYzdB2nrI3WrtSfieP4hT1nmS7bINr1nce7uPqxEjjyX/fK8NpSpQMD
NWKhHBVlD+D80yB7vJCzBAhXWE8p3DFxMl6xiq4kwIADTQ7IaJhvNZbxZ4HX2eUf3P90Z+EbQdKC
UrUY3UCPk0iwaH49tsq09/xIHXmkUkW24v+LQM75URf2EUsNQGv7O/SHWmInwpDrVlTFN3c7DQZq
bhrxJA3Shs4sTMkxFnf+3H6RxQXsO9y8ML7QM4eJ57IGoYa1TYhkaMfcDYqMQC8IA86mEMXCfXl1
dvxOEm5WXaxidbNbQlTLwhHRjiP7/7mLygqMAwTH2gYZOxrmek0xIEhYLrC2E1hdJEhPK+m5ATKC
Xg65uYAAHkRGRdHrE8hIXcRzw7g9vg8xtTkgNfL55/LMyvvYCWd7ycM8SVRuvD3+fIMgjw9VKLeJ
IE0ezkll9LZmFZ/CRAwWNBL/0ShQm5aSlxyjYPZwhPLxLePBZoJEFOfaUm1tUEZLAkEZjxd8SNZ8
oljhRwmPjmcDhJqqkiG8lIBpOZr7yK2AZ083paJHM2tY69aOa42/cgxAJRM4SsXcDnxuMRIJl0Um
U6gVzEFghziN1u60Kwf8Rwe11F0nztTglPzo8Kz1LPSYN+EgjLO2NOW0BnHJfQGHmiC6Z4OgAsST
rPrai76CdA9LpHI/IWHAbcurqBPF71tmH0Xx79Qf3oP689OHxwIFEhVR+pOpc1JHh1kjklO+qzNC
F3c09ghuJ8X6ik0EkPdeMu+yJGzldxDNqHLSwhrEITHU+Yd2IqIV6qNx8oZKwy7YvWwM86lyewzG
PkjCEOQqoIeXLpotQeFVy3U/J+izzSgPJC1doQZenqf8OzhFZfhzEImYCFkWtiqGQ+stmh/OWIlR
anP9k/uXqAepIEE9xUSyqJNYeZkNJnlTTAAHOs5yL9HN46SV9QyduCX2aOOl7HD1FpmjJYmG6zZy
3MRNm/IUrY4tpjcsrjLcwJ3W4t6twKwOTT69Nl4zmjTauGowSP4P3XKhdxuC9cYZweoL7hAp0Hq9
xoZkFNcpZ+PInq8wtmmBek5oCeQMq/slA+/AGe+boUc3/pcgq+QvBOv7IiK3rWSHpmFwViXp/xF1
qgrNHgjU5xH+l/17Nfccnw5AytHPtpAa0vQboP6ak93ckc2iRWan0xQsQ6cSxuJkw2Io+Djgycvq
M07CKrox/cQ/+X9N+y+5C+cu5ZKFxXy77XAdvL/Y2AL0AzAn1Ucl8gaQvZJP0/8R5TmpDT1TRt41
ECkOdhVgLrG1Jf2rH9J44TwGoKCf5Bm1dwcFsZlgdU+QdswhmbVnSeSJbh1GOrAXfdBApIDbc0pj
LJh9Pm3mF7nAyquZTnInK4Gxys8TPr/Axzx8kb3u4clX7zfJ5Rkhoii2Z68g/SSXGJ9A0eiHvS/T
8ezo9ljBJ9IXW6ooLHVezaM6R7eqhfZtBnvpAm+qIK8PfrNoQ5qQ5AN6C3n7NEyd5/rwCdS4MOFn
LWvHBxtEF5KxgK1vB/V2CO9glOY69CqVqymTL+62LrqjfpLsHEn+cofVvlf9YZL8h3xBXv/NU+e8
7a+qEt10qINLkE8cSysd8wWeWfrpdbbqxI273hO8wR3+UmS/llsqqDs6h9/a5wcO8yygNITPfNJY
L/aUM1E0GQg3GML+1wWS4atJ1wHpSblP9beDmeddOnJZSb+mvFAxjbbb9tfD+/YxA/svbYoSsiT9
vYG8MPAgXioiCJG08wHGkghK90+lFfz154fUeovhLCfoO3csdiJfqZIKPUKeMLexjLICJLdft9J9
oBHwmuN8N5LOvd679YLVmrhxXywBMJtWRean5TfXnFk30xnSYSqhi03oDdZI/k6LDAlFsF3p9nqi
6OcXi2kNKgdpto8YklUNabsvQ/qXg26St/ZScJW5iSeyGACikSBZj/RcvueCK1v/HeJtAERnuNGo
q7h+FOeALOc/2KCkUmqIBbpPYA0zsZM9gjsO8Z3UwPqZQ1uLDbXDag0QUMZ4ttCj4D1DMqnG3pfj
j7WbiUIuIhur/HMi8EyAMKoUegwtOxRfWU6/hvgMBQch73RYY8jAIPUltVf2n8Gs0xOtysvrJ1Ki
bg3e9P6YO/PM+t4qZZbhmUjYRg+WsyX5uVHMNO/jFtXqAONEf2oOrsJ4wegnM2V7kh69zt1oBde8
WPFt5zujv0vdjtds0aJOq82vZRA4oDYtwYO0YtKR5q0bfXcomB3ZMHrXy82q2n+hiDGNkQRy0X5o
guJP07WOqy8T/kuiVs+6qFjEl6Ek+vDwWP3ozQs8wV8a55twzBa7TBI+BxgTOcalkvGSPvDpLRA6
7hKcEceNOqpGwdCvMamAcvtLPlP0r22Bl2QtekO4yxckhiU7+agcWxIACQ8pKFolUu2NVVcTvxPb
kQfenoevOIZRmYGj/CIibN+m3BYHkGwX5klsc6SRcuv4hjVyfT4ep6CiO8Vtrc6QAcMNadF2bu0K
pQUkHGxMhb/AEZkZuubM/WhaT0Gvodqq3511YnoA6PcCfO29BK/3g2W2+uyNFnkuLs/d2Ktw2atK
XzlHBpKX5NDCoYS+9xnr9flvFSAWA/Nb5YXFERfwddm3LlfVs1llLVXkJoIn1jjGn2nK54+iQlep
tiVb1K3uGJVNzIccrgKGserDlhPWoAYCovQRayHYnsdTZp0MheEPAQSFyDNaoL99Ff5ZrWQlsFYB
Ki+VNCYaD1Sc6wXjwAazwNJFBLqMyKVNqsj85ZQXmH3j1hMytcJgwZvt2cKYfkniPS9R1GfF8dn3
eAu7tckH1UGduvGtjZkwpwW01TowI21Nzxr/Wai69Icuy7QNDu2g44hjxgu6cgAUVpBU+6EFwnG7
RxG6KWYts6aSI7PE5Cut2u29HIFrRaOCQvRHTL5NO6zF8vGrS3HXDDy5c+6++WtFte2z+Wyh0uZZ
f5lno9NgdimUAHe2nAE26E+5iV3ilRGxGs5tz6sBMUjDt6GqPw0ejgJgQ7xc6cX3PuQHwPIF27AP
XVqu5Lu4rianiJj6PWKjj1SZWK+E5pT0FB0Ntm8/sZ7I56zxLifhiYOQsN07/80FYWmgxBViT5UT
T7jDnyDaW2eHvbeNn7gG5Hm3ceBp0s0ajGptEf2JO0KPEmRVX6L0GiCX58ywAKLUWFJWCgVrs6dn
gv5iEv8UcWWN1Nh1o9DcY16Srt5TMxrjWEVBef/wrAqpyJ5UbLQ6iPOTuUOra6tUjUCibZfXmCxF
OT+mGN8iWct8XrDZwt1nlVpriy/keKcUiTZkCLgaIVD831oKD/DQhxJPe1PYIjg6BJeFXM68p12I
LTViC8ikDXrLtCdI6s3/YScmAr68ovN0iBGuBAUgNi4ny+XL7O9OtjcURGK9WKo0ewCLWAiCAKO0
6zR02fCTQmm2fPuTRDyXlb1RYPcvB0Tzj7uqs7+3cVCMn8f5MBA1SB1YHquUkohTEFPC6QizsK+5
maymJF+Atdcu1/fDdjb9fIHOIyOutAyPSphaLMG5Ob9OFA7qn1dmjf0qywpl8f7fP3VismVZrf5S
INBmACLxB1o5sEV8i6WWZdMWCoFfy+J2DcS3LVzvEGePRGOwBFg7dHq4R4SPMZD4otb/yqlXXEgT
NILaeu9uQ2Ly7w5vGzTu9FBai+x52fKKiYmbHP8IDlt6bIWFc4at8U0jqhej6uWqWUiJ6nOIxe2d
3nbgtNMax2EQKWPTqEJTd3VR5cinqHc9S9tl+WS4nHpC0PYW8wXH+ESd5qP91ZdrPFFBYjHI3o/f
evj7BVQPyXeHGiYgjSVNnawnxM8PVAWcYl84LqIUpBVHm5ci2GjnkhVt8GgxtD4I2MZH1CT8gN6d
7ntaE7XkmW3nd4dhikxAE7cVND8O+lCQ80rtydZA266AySqdtkZYE5hZ+o82EQb9MkjFCx3pR5ui
36ErkrRkxTIvyK3BYU915sw33W7OZJblJlh1tFXJ2SzUZr4QksIOvrHBzirzCquFLXE2SuZuoatP
s7OcGI6Az8Q9IEv0riiM+tlG/AqVlN2klJgLhbFA8l0YNIzYM78d2Q5xwPUQYF2htPKWKTjbH73V
VXrBKTt4K3JxNhddMf3f68gXSWjaRHK1k+jmRglfX2dq5LiF5vItHV+aYMW/fPJUIFtZFNN4wB4Q
pLgAA0XB+iQhN0hwhNXlR5JdzrkTPfcz/6CQOGIk4JFCvAWWBlVlXtMBrxI7ZbzwiZ632fFDHZqY
kv+BZcTJ8gY0tKMvrdmXAs0Zga+iRcDwGNILfM3ApLsxx2xvE8F6YQtU/tzVgtb+CkQ+fX5M0lH+
2ciaczZfO58UlX/T3REAxxMZQ5ZnHXy0AqodiAWmjHfH+l38bs9/0rqoni4pIRurDIe1z2mn6Yyy
0GzuVmfSgYazS300AI1OMcgZj3Ioxd03gjy4of2//IXrONdhrlC4VeMEum6g+X8kOKIAAys/RFFj
JmYu8CYd9kDN9ru7gKR0CcXpREl/Kzboh3n39rm5yoWc1ciE639GPjUNvegzkeGJm7blkmrVgFfr
fW+xXPeD3n42PfLEfn6RdmNfwSG6kEU2KQl7Ga3iS9LypMob/DzkqJ7iKJCanreIaF2CDm0mwK1r
FosXRDIJSt/OVD4SmbHXDKvcHiqrk/Kc/Jcc1eALioGdxMZgnbmxYkbFbwnX5qN3Wqkq25Yz3Z/1
dw5MZl9JbgnaP3VA7ct+EWqTv75y7QltxLbWo00zdym1MmVWLkZD8OVaUTzUD8Dfx/gC49p74qJM
/ROIy9S1XHfgU+ay4lfYY0QyFwENT+Zz8zaqCR0s2neggK/9ShDQoVCPlmtrFXma6K9ACTCpI4+b
IoTMrCjTcSpKzwDvSneIlFSGlZ75VpN0vJIrccAutWrttuwsDeF7sqDr2UZW0Wzb/VJaQK8TbEm/
zn+Pxb4R0bmcbpVMtKsBiXCknixMvN2lUYFUb2E/9cx+FRGvy5jdMWPCrW9rRVkroZ6fv3rdMdO9
dfFicGNzktOm8PtzQogljy/birwBMNO9jHTRs0fslDSrd/joKk/PokTrCifF5xZWe+EDeHuffG63
a5Zu4/iC0C11iVooaWxP7zrqdL5HJrXsAuVrbcyfMcEWTuMF3NmCyw1q2MICI/OwbY31U5vzl6WG
EIAtiQl3EKSgr4tv30HjkYQ7zzJ7Lp9m5wEDhnOfGqDOQFgigLF1ptjxuWhpni+EolgZFqY8bXUz
U/noNOK/D1OmsdI4Ka7LZievOWmePaGZEzrG4/LgLVU1dQ5tx/sug3NbjqICQt9o7IFxiqmRU31a
5obvRQUIAFvK6abTWb/RBypKICiHdGFO+9lgay4qkyhKodl8DiF6napvUEep8850lLbEyapDPesX
gONcYtwIysG6D9VJ709BRvpbNPyHzzCusgSaevbWE4dl1qVyJ6l78TafDogwemJYLTeI1/zHGop9
Ew2ynimg+4SJQjjxpFx8UWvnKNbLqvWYW+enmw60J83wtemOwAUOSKPLFZ/90pEhf1a7+vtAXkwD
35UzN2/DKi/eNKl6aFZtRKrg+H8wJCJZCXYA+R35L6Kdwa+bTdi9GTcXOMCkG/7nNspz8xMqERVc
yNn+XRSbCA+VZ4knkGQp6zHWkJeN3EGQ7GgmmDU/ss8a8w6/BhD8PUXXPqaEXxPoBPLNX9x0XEM8
SRS08q0KSlX/m6ZTxX9smueKVPbx7F8IOn4FxjNiK5KBK3IMIpj89T9v9mX3mSpyGjCBfjDwkRNX
eJvhWqfeFFhROHSnn/fc6rNSvc6NLV+Z90SuEuHqCxaqzd7Bq5bcKruu/IyIAHcXcflxUBx3Bpkk
V4jzGZWS50nbNtkaEGbPxbAlv1V1K15ALH0osRULtLeqIDTDEGQ8KhCGAoVfc09kiwFI2uDmdcD6
VKcM02UB3SM1VRq4boIMyLjodeJPygO9SlNqk2ZOCn5F3hjBw/8dGdcsLgPuIt16DQtdefEsgWm0
MUgIfjwavut2y+WaqzkXD8qiQQCa2vBLz4uYhPt8Pt9DYV2pVlU3GqiI2DsJtDOzljxXEX26aF6m
m6OeRw40vlkaImXz+Xuix3SwqUSPqufOJP4hkVMVwoG9agtfZS5Wzhtfo9/GUD4YIBfr06o5D6B4
cc/kPDxXRVYS4zaGbxPJDu013OSzQ1zlZyh78+HLzrNYJpvZzHPfMnOYXqS6lWAHhlfVUcAaz6aO
f0X4mBudqLwgPuzE4FU9SlgXKEh9zxRDcl3scILRBB9FbQ/vfiyrnucZ10jLa7zsq2mYsZ6NmzTR
v8GupY+M79nkme7aUdN4xd6M3uQ87hFV9LUCzFFkkMdgp2MEXktJ8rSPlWkH26QEKbYbG0PQ2A+3
lP8l3E48aKD8IBOHadncjJt4c1ax8UdDm4ygyGmafJkZFsAisecimdlZ700YPVcHbLbhYRrrfdMC
8b6TqDGrxRLpQZDwFHOAAqWsBeYWmFmyIhRCimNketiMmeqDg+YgK/ZyfgCOCi0teRbFxpuHbIIQ
wtrWDtn0UDMnmfReH95+IejdpMqSqCl34B/zaP3QTdQXcHmnakn17L1TGMIp17CqU7hNF7tNnJ0g
jK5TMTU1+c9qp5TXbdNts/cysu4qcsWPbzsLFyDYi+KsBJvThlcusNq8/G6F3Uq02cRFYHhu3n6H
Qnirzewl7fovDu+w+YfnrR4gsr1krB/3tJgYLC1ca2aJYLkzx4KWft6sl/Ky0uraSkeiwIObyYQE
SC6NAtCmE/RXXxq/EdyRSHpuLUXjUbsxEznWwqD7ui2RjryLk2Gn80UgiFjpBiRlFIGgbwc4INGe
5z3yZ/3QWm6GqSQXQsvTlwRqQMr+msrLu8ZgJS0uXzi4R2AWL5Y+vansKT9uazGKWUqn4F2lYjw5
gjNwcPFqHH321B+zfQz4brvRrlfRtK/XGZZo4lbaiY0rTlnZ4fnfukoxd1EKAAXGt2IMFTtNVZ50
iXW+Crj5MvAmI/bq5rs9r/nPlXp7ovolJn79HAuRP7HD9Xiae7J4Xu2QpZJ3GYdKyxRz+zGDjr1a
FqfHJL3hlIO6gnzGgdyAiHYD3meYrTD76Imqtp4UEMSBw9Lc1ZERXf/0SQcxcwFsmZhACY7xoBXt
qsrT++F/MKMsVqOwy6RGlh9brv9SQjFNhB5ZLMCVu1O2+2gm8RJ8yKbyJxSTis5HCFLda/I1hOS2
HtQPvGHGy21cCJO5tiN4xND1GwcKCmNEmT0c4LYMi8eaPHz3mQDmI28qqMmCm6UAL/DXgKom9byy
MnYq6kGYf9kdeDCz4DzKposR8XzQdeKPM3/MwYEab9oGIhN7QAoeEonlFtWj5VzUFH/iB6lwxcUE
056LYPY3Zl/d73xEcEFNrUzpyhkpGessJCsVXcTKYM7nOT3OctdhyVmLHWgA9HSLmfvv2A1jILcc
j+G2CKmIAXP+Fd0qJ6kRUgKuRYiur1rQMPBmFhUazCoUeTdR+oGzux5a5779doZaB16kwnOuL1zH
DwRemo++iA6fXlD/T/+SpQurMYdfggFMEvLmZOj+rXU9USAKVkkkpOzjfsueMYH9ewElo+6TDuFL
LXKBQxtI9D+liRR5rJ0iGsn8vrEPf5f6Q76I1YbJAGbRSnQjg8uG/nvhi7Fp70lcjQejNAN/xqxU
MsYxqmN/ZpF0MwrTeNxOjYvxah1CpjQJwVU2Oz2I3zO/ZLW3SrOR7GfBoVw6k5Vn/XRaBvgOulOJ
/OPx/kjc27M50XLwOe4Tjz0l1ChrWpGyo40r4KLQ5qlDrF756LIE4qhhHoeryqsLr+XyXsN+Wh9K
rLk/TzuW1LtNjMFIBNcQPQoK89KlvMWw50ko8K31ZobKCmrmYuPdr8BsXJVXUG0hnsjjiIrC+Jt7
ncQdiYSEmAOJ6/fMrJgFOI64AjVlBjkBX2pzleGOJzBN42Bo4DiF9JZVVTOdDsvXcco96kqbB8w3
QzjlOva+MoVcHBE0d+OINFmupB19Z0f8d04oKGyvG6olZdZ8GoV+N6Z9/7QCTxv/E5h1dY1igoaB
ycP3P6B9ogRp3FqlIJUYjT99oMsSkxdperBS+mz/hjDSZ1Ye16IbcfsvhjozhxY6JT63KKxnkV4K
RoQyvozNmwzzvQTtl9HCDqestP6fJb2iSzsDfWDRSBQcoQP0CROPwtbS0X3gw9YfuBDQ5fvK2Kdm
N+79Q/q6e7joUHPy72SPdhmZJ2u8NS+7oE7WV/6aDq80AFA6xSji7+yhpx8xuvVC1LYidKWUTNf3
UCdFQmhRA/BwZHhuWonEjoVGA5FHFfo8gn1flS70TeJ2Hrv2OMbmj/tZdP8826UERc7Sx/yMMUeG
mF21alFSOHulatC10lGDS9H3nKkmweLJ6nGrBJmL3CjJM/7UW4hND8dss5r3EzsulJK7kXnULJ6k
bnD6TlakbjaLsPXzsP4mJtJis2b7A9qwmzf9xbQao5erpew3bOj4yzS2AkT50ORx/j5lFjzoe2YD
BMEgz/LHs45Re8UVJxdlFYCmFo8h7X0cRNeNKl5zY1DwEMxDY2R3qQ1/9r9Ol3J6XgLS1lZ+/oBe
nipqxGQ1NWIIjFlFYBgN0j2yXrTwARR4KM3ShcrJc0wtien2yh8EUohvgoOu+qkhk8/Bc4/aHw9X
0C0b2qBAcM7n8pw65KPgDqTFvmZC4s9RN2pfA8G+VrlP59/TsD5WWjyRsq5+Fli8ayszdOWBelg3
yGZOcjSm0KHEm1YIUrL3A3ijUgNyJUBOZxmHb3XqYoV1KCVRbEpA1hHCJOxfmHyrkSHAiIw1/Ic5
eRPiUr6xhCDsw4z3YqUoO5/rFBBURGwf8GJIWpPzIxa36g0PBsPcCwOmSqFYrqHFaqpQBUtF0Rlk
rkAg6uJfuR7zEIbGBo04aTIKB6xyLdmytMwE+pFCASH65nq4BmjvIY6p9PtHwjI4m3xG3a3uNjsS
XwP8kcGfhwPta+q7Pr0TaDzdHNXTxxlqhU1tSI8soTZUWaEHQYmq94wvOxIY7/H2LVCzPreKy1Kz
WhegeI25pHOv2DG8Dl4xhZY6kNpQjZ+45GYVJF7q1cbD2C+63ccwjpc3XjWp1cIqoAxPHowQaj6r
QPzAOOz/V7+2JNi8hVdOVOcNKeTQ2sR2RQGwRP+k5o7Qx9EygYVlIV7gpcCAa+ast8o6M0SfvBVp
7CE0pw7aEfoNaiF8gghdRysur8nBkNLTNdjos7KzGwTNjsu5EATO7g1GFC0qxx0YfBxEHCdBDDQl
q8F4CYMNuLN9DrFhTuoQEF/n0ijWezsRCii3DHFWjiqcZmna4kGGREv7TcY0j4blNQdRwyAePZTJ
B/aw/DfeQ/r4ijp+EUX82h8uS6rXfWJhTz7QMuUnLBGoLledX2xvxAHFd71G/CtsYCaGhgFH/EqF
LHq4MKMwU/GQBpmADnqo5CtvRK098s9NmdEE2N3ManPqRPmUG11d4s8nk061g1/+H44UhIcLBBma
rhdS4UDv5SPy9l1JN5qmdGsPi//Q5z4cptjbkqD+6QuX9djXgeCiRJKF96yRUOD8k7+3vE9HH3U9
DJKIS0tSemcBcec4NArZoN22wwPf8g/5Y1eUkHmP6rTKyxVmyPGspN8E8bSpg5mL0Hkxe0lDistx
u8WhNPlmebMaTKu2WpU7JaAajfFu3eDnu7Qht8adEFl1cqcF2A11McMAAjWxuAhzRXku5V4HW5gI
BaRo1FoAl/+0XgxQStGJZy37GnreN1hG8JS44eO+ua9wlxeCSya774nB7ReOgvs6h8nzbRHZzI6Q
Ew2gzl66+vcPOx1Acifi2yot0vFMoaNE42A+mTd74D+u3PKILkcSCRHyAi0kz1OFtcQkcGZiaWQh
rzDPjwzST5N6/9JuLM+6+JJxTC/ULtD3ljOfpBygIGVZh3fjYWSpGLIL6AlsYf6bOBymwB7Z922t
xuwCH2VCOzu7Fniin501woleHV50igVucA7YuQIKLsvqqUq1SMh8QkS5Vbby+RFd5vFYVvYJuy9l
25jGaH5k5mE8oJWzF7HSg+i9FXLOJWDVjoJvv3FjiNQzMrEEEPoc7KEc5e7woXX1Anii6wb8Q70L
pKd3yqViGERz/AdEoXtMG6nU+6fsfGK4Kg39noIHuELpt2VlI7e+khNqGWeJNpVfXxfEIcymkX7C
NUAEcLNbNXjxRpQu+zLbtJNpoLcLDZxdpIZOoh5MKIwYWYl4aLSq1i/ct6ESt6W0YptrShRHjZSN
0n8fSMC2aJchieJ8QkhLsnXRtN/2iyOwvCaLuNTP64CdfVFVf32hIr4bIqZS1B5Cdg6eZCoyaFpE
G3vkHYzGLlG8gbBRKhAvde/je/yhnsW673JfQLGF48K03nK2jbosw0yFAXUhRi4gOtBqBJLJ7IFg
Q4fhZf1A0iiz2J6O8MK6O2hRRHLvUSCfxmrA7UhjfgA6mdVnYSOOoZ0q1s8K7Q5q0iIYPJ9BX+Ts
Vg5/zfkon/pS1RS7QXWy03KvtQq+/AhoQqE8QCGvLxvUFooSe4TEGyPtD8LgTewz5hS6BA4dS/an
n43ToT6CQK0/2Xnv61aR7AUQzB6s9NZ3cjUQmZ+ltrxOQ9cKiweAzYdXq4eAHpe7TDnhdSVXCYxo
Pf0Kd2HtuvzRalkG+HCYSEzECaVHfRcl4R03kcnQ8nT/g3yrkes8Ovs91dOFSi40t5FC6x5FiAmb
uUUcLAa6X63GLGYocBp8voR77PF13LratUXXqJanqoNQ4evYbcYHOH6D0IHmvke4Rd69cKJkChQz
0/ImKVw0HXhj8PBmfkbS+bBQ6FCvRXHFvD2UAWZ9FMlZ0hGEJDJDmv3HMUAxHXKH+Q14rgzNxqEB
wVTxKgffXyPBqXFjZYPngh48mErvGUmOaZZal2U0XPJvLm7dv1pVNdk3H0+GtEkchyTgdGOVNrXb
cYUM7uw703e75OAfHVuIda3UHC5pqoT2AhXP8gteCxmTocA6CdoMLZo001lz6PzEDpejLJFHoQkG
avqh22t1Gt5sumy6++OENPYdJcPfNEPg8DSE5QF9t7Vt/ZXmfXE7ZOnDo8hqVo5LJlQ8oBRuupia
FrHm+bUM8vNc3XBEqYHI56LF2+7zsMBsVLgKPfDiZ+gUR2MdMnvZ0R9AdRDJwUzZB1XAnU5qw/Sm
jbXOgfGev+6UN1RYVmoNtRlobTt8SGrt6NfJT5IjbGZ23dRrx23+CmiMdp1ocn2es6X1i55W1wHP
Jj7ndXIf9KQeuQQ6KYSpPv90eijTcQ5GE/V6+CEXrfZ1R/0LX+zz/2htHjsW+uac6QN56VRXfvrH
DSBj1icLsIitVQcCE5Ul1vf+Z/Izw0PVOtAy+A4CKdJCyN0HyKs2swna3Z4nfhBX1O9xAQ2Xpj8q
Bu9vHfjk396EJ38B4PNRcMXNhXyEy0q3jc6BGKeFfGbaBONhJpJ+H3fCwur8m/SE2biqZhs2li7I
iNcV3LaYKjz5zQu8zF1ZmP/w3tamfrTcEnc1wC3tSHMvTnLzm5ngGUIAurm84ET+D0WR9Xxnq8jp
zF3iEIZmzrgig9f9H/QVepFo2iJ3X9shKXe+Upq4NUk7MNZHneSwd+5GAEkSQN37QNIK6+TYL2F4
fAmXgLKxlkpn3N82xo9JsqpsRwsS6IiF3d6rBp0r3smCIj96RKD09aTAATjiwxzmHZBlBNVjjJrS
YXSXvZg2LthLokTSQnt8KdG3lSytIHDopaII9SLRjxDx794FB7DIktbkmUoBrww8Q31oT/e1NsBa
XyY0JTjW9boZiijwrqFJI2B9+jdzlPjqQfdiyCIsf5tKCODvMc/miqQ3jWAWOKepUTNJjuAayI5S
Z0MX5QLPZCb2zXf8JzbJN4po+GIbK2CW6pX7rqS/hzHFSV7VJmqFgqVrCSEfi/sa061HDOi3v7Va
b4m8lsqyNAiuvTMr560OCoHX09VkelhB2rBu3D11oMjJYa4k7p6cSNKg8Qhu/60jUwkCvF1G+BKx
6+GXvHD6b6hAcG5qvBXUWRMdoEUsnGPo8iGtUPChBIsDFgAKejX9wbcS7sMVPR5cKLpRFKgnraJr
Wz79bhhGbvUOC44qMC8/ckC/lVnWEAF6FxzIc6vXx7QFd9UwqUG6trYfF8MQjryttZXL+WZYbw0f
/xwPHRWVjgLySo5XvQvQa3ULlX9cFcsmMksBA7404fnLUJb9XwF/truyNVFrHiw+TOd9wZU8Mh4q
3GNZU0aenYoaZRtulKEnsbU69jyYDFe7z5cRLx6b9IrerlTzA/1nRq9gK4GdIMxNWMog/71/zGvF
Y/tgYhed+tmNL3dpMeEhUIh7/DYNQlLcP7Or6MXyu7hE6Qv9Y6o2O5Ne0PLN5khnzSifAKZvKg0B
u4SB4MzYqedu3u6NstP/LMyt6i/l2rtBxYoAkD9++A4TBWqmMZtL8fTKYTIv1kSBAn1Nw15zj96T
Qs+IzKDxjVJ90GLZ0zwNVQ5p2hfzaXxCP1FPPp4K+s3BXRR5R4bQkV9QFAnqeZl5K/Mhz+R8VvOV
/1DIvsrtCYf9V3UbisfZLNiEQMmEuZwHi1xuFhTpne1BK5PRdC7vzSPv7hElFhzidLQ5YJ53ESBZ
Sv+BsMbTcKa0Zv6UYKV7R0ntzDHadei3eT+AZP8VmdsmNZAedzNLClR46OCBYJAqPVoWkJhBCi4i
rSASftuxWA6Gq3OBkFy5p1YR8GQAfA1TMwo73eVcJWM39XnqggX+O4/XND7xFSsRARSNY4YqM73J
5+AqQa2VQdOKQChddH/jV86da62FLB5l9RYg4XvTS/1/PZ0jc06zjy49GmwH2NYVdQbKoJ02+Wcb
9K8zTwE0J/f7bJjcw4QIfP7T5jmBFjbw7x+/BP26lq/6742Wsa0KELItvktZpTWqJzfUhAuOjo41
L8nT73/XIUCbITl470A1fb1sx8Oyu7LbIKhO0Jzvu8WzHAun8Mdk/WIWhUOa4jJZngSuBnzKFnL8
uh2kJ6Dk/SVU8dgK8raoc6IBWjYhaDp7CD85p2d++6sgt5PopXS0hPvIQhidodEbbvnb+FpGWS7L
gmj3DGKM/EWJSZNW0PyJK60COijs6Mc7JCVevKd7oPjsEc0ignM+coN3sO0ueQqIn8IG+ZH9kVo5
pL9ADsMSDqn/eGqjIQJRzGZJmLpwObRX/v3AD9YC9llRQccG611y6HefIW3pIqcZ0pSfg+9+wIa6
0CLtZ8wQaN6nDFWrgYKaNl0osWl+LoscmUw2it+holoUlKiguQhQxzNGpP/JeOHH+jW8GksNQhqU
P04Lykp3YO01CwL2O7M+wlqH+azvkLXPHb0cpy5KeAq44Fc5NGt+eyml6U8HIILWQbtwf8kuXJ/V
WoKdZI1Vj1VVThhcOYnMKoQYhyteWgbFO85TQu5mhSblUUfOxhaBAW3hZTvyBxgutvhAqaHcJCKr
O9BI+niM27OwL2nJMZ98rXDFQtaZ6os18Goqs2wMTxUfXUQNrZLLIiQFQWqI8fQuHus2PUKms9UD
uAHfu8Wu2vqlWTqLMYD9l2z+DN8QoGMoSd042qzcZ5dz5eHGghQexbD7TsDLGP8xssuNsgeLc685
e65lnn08D9LJrVusHY7y0mgZ0hZLdU/dTlT6dIdYE0uzbd2WhlqmITDmddqEBdu5ajcbSe6UyxRC
bXCfXi/qFPTkXMrUyo50y+ZNPP/HEpW+qUodj9ecKy7CSecWXAlPo/yDLH6DskgR/p2gNTdvQdZC
FzgfNmx044iTz9cNDS+OOY7mx/dM4boLOZ2JbRBZV/6sV68YRtfIvW+ehOxQT9zlYRI7oIOM2pq2
3op/2t8ZlmbtwnpxokfDJx2NYnDKoOmqnZm9+I2BS8OEedloCVfHiI524Xe10CwCb6OpR1AQDr9d
apdC5b8LlG42h7o7ein7LbmmPNhcBZQhN8FaZNzVNXi8fK/9xCzra9HH8w1fLEB8LFJD1X5m4X4/
x0iHTR3K7tuOSv727T+ylmp3L57ssaqfCdsZGDYuEqqp2dzxxd3Wnu3F3J5sGL9ED9dpmASX4h4o
keRIRUI/GZSRoazmlfEiU0BkX293QVJfdncv8Db1FyCSS8+QCXDF9gyX540gZkf9yaj7eCmfmeQ7
2mIUZO5t7Fon8zLbhCuuq8LP7FgZ2nBcuAADtWZ7b6VceNpmBdjVOO3rtqJGzK5R/gRXwOYrnix+
gex4eBLnU4ktw8IHc3KC3/q9SqKR5qh8pNETAPqIKtk+DmTs9H/OGRI+HSxSkVl87259dCkXoO4g
dK1n2Duy9slZHUkysLrAGZ+7fB321bBEFhbdwyLImksnpMVb2S8sLQxU8fKsu/dsZQoQabFyKp/e
9tf67U45ZjzW8DLxecOqk+QATMg9I+dNSY1RV8H2+9kUY5UcgTAT8dkeEq+AnIHPD36tGvUA2cs7
XjNIkdZDQOM3dNdPyfFpA/nKNsiETMc06izZu/Rq1O29TzianAwi1RJCgD3p1Txd6VBO+Mn1bUI/
fZDC0SicGuNEPbT5Xy2mZ/30VEyEM4nNwiGG1D9d15z6KSVtAeAIKtLf4hayflyn4mzaPnovgMzb
WiqB0O/d/6U+IeXHZcNbPf2s0RJL9yU0xkkH+6QaVVnshis91AxK/Qhd80XFnLl4K0cnj/CrrQXs
p8itMaXeLr698t2Cx6QNmfGHP7RC8kt6HFttRMXNHu2XbHy1NUAn7Gu4/56RDnz8/zVP0in6P+vN
fO4xrfCp1nebw3by3NLPD1RGpokHPBUPphNzPitZx732XDtr2BXWC8Wb95nYUDDZMSecSgNAO1Gz
lA3QkRSSMIdXGhV5dQLHTbUWBWPFEWUTT8GBvgsPCoXlHIQJblS62pNpRGCMu6Gjj/isgIMNQfGU
lr+PM3Y/pVRa5NTEaDYToXqOVO469ImtIviOHAtJ6uGAa4LXd5H6Vkx+rJ8k7+1qIuRDg1zGbgvp
fnd8SV9sqWOaOitTH5OsDFkYTt/V9fDuPHOCucxXiqgIJUM3CwgCFtCYCfr/O9zHxBYAutJd7NR3
iMVseB9xiLkYlbMi78GPmj6yEYAIZPMAJ5mDMnhmuxvRN8N3hGPpZHp0BZ24aeoXKK9fXtz2UAMC
Ojc9eWvBUiSAa5NVuJ9lhV6uB4h1q4YRwuKn1OTITCCf+jN65OVI09p+1fWYWN+Ut+QZed/M8J09
I0BZV5ajDLIa7ERcyOQtzT0aRKFiED6CSDgLE/ckd3+UgfW83qJzj8oHTNHYTZOnCKYYFImEde0T
F9aNmx5KFA5qd8Bx4CFfMLtaSXmwfYcGozgFkPFMvCUAGodsxF9ub5TNATsF24Ca4vqHZYF14xX4
rQtUgAomYkFaQNdwTmyon12fViL5eVUlEXQqf48Zasbf/vY7Gr88N46VHm4bUQuua0ZnLr9btkU8
UbUIUyktwkskb5DTR/0rpIYyqcRd6qbyvY/6PIcs5suWsIVy11qK6G+5TOtc75Nl50Fh3QWvF7ZU
kCepNFEbqeFMsrwXf0+1jk/vNV5mMV/W8hiSTJmORX8uXAk3IpHrW1ygslQXLap68sdXEjsRoifS
KeXQRffvkOlkJbp+6hKH2GHK8TPpaIB0gTHsyvyrbx9QT1Cpr9owhhM488+ES6rXgsv9cFiYuWo3
038RhXWALedO9yiwOlE8dfTiKtdNNMIDRU/BmZA3m56ud6hRbS0SSEmM4hVCFKP52zeCxVchUrs4
xEPTtw8ilk46aLTZGLB8a8p6iLPxebG6l+fSOS9QjYGDRcj57vs0WPlNruQOZd+PGirJidPtFLff
5l2TmyLrSHyoZ1ppMFpI6n16vPB9mpUoubWgB8qA9WTHXp2QDjzdk6WurQeGnY7TFEHXJ1nifwpM
MYNmzbF58iS0xTJMWWa5zR7ynwxG7Mlh1dE+R7wsMDtDAWB6TQfD2LL4QfqNsbwClazRYW3blbiw
DOW3kwUb9+JqJZzinxjO9L6kyiOpzDHT7Wkq7HuHzu6HesOBB+UorbW43t5jv8HagtLmnx5+EixX
XMhZ9WUd8E2EBL7tiTzIy6cA85mRkq3cQ8kj2sZ+ieTnWSWgderU8s+OUWf3wX7ZuxULX0wldHMh
5JljwSXFPRp5pS828h4DGh2nk7spq8rEd4zLriuU8OG+32vGrxf7P3SwPaewUdo/0RrPqDWNXP7I
pz4qO3vp1beffh0Pe6FiXvSSU5vgIN1LLAoj3CAx8otjAPzA1DHKssbWU668eincuYTJzfL2lxa+
1pJ0vvDbOjQwD2NFfHZK5Tv1wWUjikRwiC5/m7ilNbAORNcCmZ0heiI82UFD9cXNGbXOPdYhGS0e
xQfVVi5mcaxsr7hxlU11//OG/ESEpNAIezsTsMkLKcSX6BP+CfIZHiFE7H2augQgtmLH8hNdnPza
onWGB9I+6NXq5XUHV3h4e7WRnoSp03YDN3JC2cvlisN8z1J23lk1mAfRjQmvKDPUXGZ+WUcvdGC1
5GQ+UCCu0OthnneS+MbN3jPfGPkF6KoztNqyOWm7CYDkc+cqgVqZ1t9AOBVliai8pte4rjWjoa12
OC8NmrC4FLTyKUsaK6qtm8GEOA2CKoCwup7bgJ96u6ZZw6zK8/HLK0/iQlOqfjgpneyG91FIkQEQ
L2yJvdl7vH1rn1xaaRL1jwS40UJoB11xFrJt8O9LOe1EiUcQ+ylTcNWv3vww4z959xd6xtw9dEjc
kPapHYJw8nghrOqXEXdoohHhfGOC0Ks46ETVEC6lP4S5LpDfKaLHWU2Sck8T516LawigXgP7VwoE
LSoMWnkvrSo3HfIDWzzFABvNI24ZH8IXVgw7KQ+pya+x8HkGMTQlC5nE4fnF5c6jNaUAbLpgSnDa
Li7gikHD//8+NUu5pGjPHupwzL2xnLrC7VQDigDa0FdK+Scweqrf5VpQt8eG09udsLAOpLCQQd5R
JmR1NBKoyT+z6azSTMYg9RUyf6M5E7p2LWVEMY6BDu6a2AEC2daxo+lidcmM5Q7pko6O9LjgUZRY
VqqCgzna2IO4Q5wI9HLrE1HFhJEAoawxBaNEBawoRPQwvwmFOJXZDi6pow0pLduOH07JG5r5KDk1
AW/jGDFfu+BRFwQJgWpj8PfD9U2IzMM9l94cjEbjeXaS2wWQ3x7Nmq/Mk/SmyWReaP5vwhQqNa0l
Xr5hBEYWVA3TF/4/wskkSVwjsPiDfN422cVbGmLwW6gaMUrNz0Zm3wLB+Mb7dyKRHbv6D1W1Vm35
QDElOv4hEFZzy16qpgus+4whURqYg+bbzppgbfRTdtutaarHV9ImfwnWVYfXvKnZx7OveAEMYt7v
0CBIdmkVnTAvTizXh3C/4ocNs2+PqTEAjiTeCkjK0u/YI4kHx8PFhWKuPUjtDzrYwSLfgj1AHf0Q
ZUJsJvxeyKuSCLbyXhqaLwxEjSvhFoNpdplMJFxqHXhw85xY3XC7d//9w/IDwLrveMsRWih9HsYN
qCAWAw8Bi0+c5IjIApTWyEU8S+KOrYLBfqc2zSZhOPU07m+Kzd8jWQMFIJqPgJcFa7Wq6eOQC/V4
I1+w1w2SXSGe1liUNR5biS3yHSsqT0aWjGoFZCA/DKlhVSVh0w/aaelBEGc2FcUMOTCEH4ixE/Rm
cHzU14SMHAOwBQf9ysmWrSApEeHCX6pB46/KVgaudpRNJdpRfyIKAQ63XJZcQKZ/fDcXSIfbgMYS
hW5aqCTz0RXtYaEIX5z6LAHQ46FYkJv/WkPj5UStwqwl2TW3Yr86MbE0WaPnk+wZ+Rxwaf6MWFR5
xxDvO5MMYXSME4gEOKJhXW/geyUtNLjtp2EZ1kbWd0kA+qPRo2eV1cq0ezS6AdWgkDaa5+Ftmda8
IXEIAO/wGh1EW3eDNgQpC5whQXaAbRZkcG57B+VkxkqUij4Yj7ioT9kFtZUZo1D9IYuTvzZjylsG
6GehfPfgGt6u/4sXN/N27yMgo68BTZaVkxuFCwOH1H1wQVQS+To8ngUMjR2np1IMPK+Uws7/MNtq
w/Sq85RvhqCvHMomJoW56v8dpgKzL5NAPpHvsTfqtrLhcSO43I+gEUHtinLQ5i4ueu0SUlOrROVL
KSuXUkt3r5bnpXsrrFdJXqKaWSxVeO+3Td299vicMc5weZa5CCRAPq2yegP7gQXM8Ugfgj3MSADy
lJpBZhkzP4gYn+fUCh5hRWWevKiJePEUtB98Mm7QIZUlfrERAqa3wXIkRPpB2PG6djMX7cFXGWc5
FcJzNC6eQjBbtz1beAsnI2wQr8TMrSV51Co0SZW6O1RzVjmSZyEhbadDMR+9755a3/CjMlm/QLxR
JyjeovsWzlaHPbdJDPsKJbCrvibj5XRedb6mcYGVnIbofWsUJvDMY/48PUsk6W+JnGiUmVQRLAWP
RrJAZrS3zcGHi2R+8dmFtmnIzMHF8oWxFZQ2ss7tPhBS3kboZ7OUG2vKvHlPc2+DvzDsbuShyNvi
R9L79Td40159A6iFvb+2pJS2y6OkDyfJsj6YoszY7mmgv0RheB/PqhzXz0/p+VPI3Xr0Hrh9p6Tm
p5/YXA0pOMvvye/nmp/4BScMIeXKFlk8QYWYcB+jfGhjbEWigVYh42qd7EuNr4ljbyZWs15pY4cr
bMOuPhiwtWvpKJKMqJJ2p7wfyjdhZhJcAh/3zn0+ThsDV9LzylFbFl77MtiFP08VaWk6rbPB8oPJ
S7/4O9jJsqDSvKmASyFymM6Z1BaP59PuI3hKoj8gKJYch6TYHKHq/SewDJKv8BjKXWJwK9Iz6wF3
XbByU28d0kjJhv9gMtKdxCKYNELbRRrthhyRLHMrIPOrNsLQh2U5uj1fDkjD8WxrWVBNS2VMCq+o
AubZdGBgLIVx+7QuB0rC4nE3ZoJqU99JRa7qiL4P/0JasnaZjzYVwBmOmMXtZwhho0rjHDpLwm4C
ZJYMba8Gt0KIE/DYpN1v4hLWPwiHywzkwoBhhDE7VeQlZ9QhJdXeRLuJJkqlPrG6KylWH7kmdKFX
6uOkSLmu4D3TOOJZMp/HXJPGzKvTGGa7x4DRenW4o1e5Z7GuJpTfveivtSESDhxv5iOz85rMw1Mc
yi82H6oDsDWf4Nag1svdxuqIJ9ZdMsKdfn0uQUfeqet3rrWXl66f+hf/HE/wSB1NBQ6QW7SZDvjh
hUrBuN2ZHPHrVI3xjmh+p3/diBGRW9bc4geWtJCnsUTvmw+DKOKX2/qV2gIdB5IVuVnYreQqZZaV
idpN29dQCOQxfg1Dafsj3ZOSMgH01kbJefafOkplSnPw7IRI7PcmnxLwC4ql6QIljpFsjW5WjWDf
1uJq/Q0Nz0ge4/Qr43S3TyWPeycYguOXck0b+pVMmZ+NXDfS/p9M1nKxJcW4Z/D+UgR4G+cuicsk
ropwsKoBrocW8VCimWOe044DxQoghsIkbjnTitCY6qZGm04x1V5t3LjlOyKZ0nCgPotL8zHMMAVG
ccerRJVUgUm/JqzWqQJWYnRLG7wXLH8COt6aQdw2AR84W+W70GPL9foy0VJWfCXdETfMgzZ1IzK9
MLfAbUETok4d0ttgJAKp2/ADbZNT66L/TbkozPn5DzLhOROfYmrXT1jgZTWlOGu/ovmHHj8JPuWT
FnoPpM86aHlbBVkj0r84Hl3gxb274DS2A82b3FiYZydE5oo2SeqfKqQsd1OQwLGcilShnwCUJlAK
iOHKJZh5MoUsCRhMf3p9LRmxCFovCZMOoPHjhKxzJmRD+tgqvrkD7O3br9K95p4rtlcoGJYd0ZBA
itbbmc4ntocJhgtwYa1IRI7XKCA1aHVMj+UH9qXk/1fhOMpnGdHtWNbFG3K4ebl9c47aoGyI4/i6
8rtR7AwLT/IaG7PXLhhJN/4aPEGsfR7c6TkNhH5rSmfgO1p51zM5KzhUTyht8O/dzoeqmQiBjswE
qgeV3mlOqbUyeDXv9HWdkyE/AMJ8JHMwG9paEjycPXjhPuEO4YR2+MyfEXRUb4+8fM9LYJfyrjUv
8v9qDFDhIDgkaRuBxobcm6kAbkXiUqAzTP/VA2+KZjgvWeTpCG7USIziK+fM4ks8TLHqZW/kJjq9
zL4qwUAlOIA/oBfr0zGlGO1Om2OysKi2wTmnuixhw+v/CmuSI83QYoKSeCDEcX8+HR5qHv+lseku
jwChD1+xNcNKcRo1MPNCo3v2kAYcK5HUbNg492jarHi7OdBEL8nopnChXO6NkES7ox0PeLGhyjiK
mdAXpAfOsuJE6duZ4PAfkG7HOCCxxNw2j49ySAZHLip57AcxhDDveaFqW6JtNLGEgMf30U5mDLhz
lYwtmrRbPMTrQqbM4nmueszZTEkifinDYZt5wKiad8wBMovpGAgifkl6B1A+XwByjX9rTdnPVkUk
KbcrjZ4WnavDbVdtV7FcBposU/tM/psDx68SilI1bM2Yh3fRbpNT7/rZ9UXmssGYQKMPSbPB5a2W
4I0mj02Rltay466M0vvRyPLZuxi2De4tC1qYaWoJZpZ8eM4tA7BFOVTw789aNpKgpDyKsdhxkHSY
ZVP4n4h7XZzHJM3gkDXfpFt2R6Z7ZG/ESgQ8Bck0ZJwLiNzQxH6tGlFiQ+BS8sd+2Qlf3q6SFnK7
yNE710SIyLmJDgZU1iczgBRUpeYzeKQKVvhTJ4jHi7HrZ5kWJUMz0ek1+7OeB+DAejBE57xxy0pT
DtOcv8UFf9RayjNfrTGxsZ9tWnbe5RPGBPuo6xL6SXhAGDAIRHRbDp/Swi4XKFmfCztGg3UX+fY4
XHmjmlm2oND+JWZ4q6SvVJE6pWAH9HRh9qPtfSnVXOBVTESIqp1KV/sTGVk6lsb4ZgZxh6FjuHu8
Je1fzcDUAAU2bjBZUC5SC3kF+lrP8GoDSHF5JmRio6F2x5NDw0/Z968L5xUiZi4VgiSnDyMDiOsr
9YiQIdew0ujKYLf9bP+e4ndhQcd5bGnlVvyqYGOOT3A1z0nsCYqqSYgrLg/3+DfagpqQU3YxgpQj
MBmS+SQ5D7oqMZUyZkFgOjN1Pxwx1myA/CS9xwSq75+9Q2rnYpvyRRdhb7iDG3T27oiB+XfzKJHN
ylQeao9oiquozTlfNb5QERAlzKij+IWS5EtOwmb2Jzcci9xlDDV7iUFIFNWVGMf+6TXwrJaabMSo
oOKByfvuYduBERMpKTueFknbCI2/nW/ZsJLx724rCB+osCzYg7BL7JH8HL9bXpr1H2XE9BJtzDQ5
69KE26Qw+BK5Ux3htLX8GsvVq0Fio2on5k5EeZx/ivpM2rf9edmLIF2oKt8FBDWa6t/tQ9G4snIK
fQPoYsG0tHmPWqTOYe9wlavvOUCHw5CEcLBbzOmYopNElFTin0CX9T/+I+vQSqzXtGwPqEw2x1mS
WV2NO9aGRxXGEvtuliHB1pnlpdJOrUC6jogrN5Y/2pCd9Z7ldWHL/13uiTzKz8jur3cPRCD25uMY
pR/k1h7URgE0ujl1k23fqX3nw9ZeJtJJ8F2g+1izVylt4crpTeKkrkxtdX/DSkJE7jfQmxbmrqDl
f4yBbTsF8RY4xlbH3f2mMuO/lbXmgbQ4dkQNajFUn5cC4SFK8DuYn3EJyNGJm7R31VwthgRnBOPW
SoyQFlbvNybb29uzX8E4ew8ObzF7XFplnXhJGGLShZZ6qR1wuNtNJFGHhg9JgXlhpYob+tXXbXHs
MZg2Yf2Zb5Mbv/Oa4J+L2typVTPUBVP0paGCZ1WAUefHeyU3iTgyEVP0+i6aSuVwsQz+f90Mkmcy
GtHQhbBKCCx7jDF3hCEnyZfDhDseyMx7WoysAiyCT1iMjlBb0FMVvYL8rIIf/+HQZ5Z2OnX9wUnL
ACii4ebW9LLAFGmDDMH72c1ynNTMh//XRE6Uc2+YbDEqMK+eQGT1Tyw8dIRnSfZbGqHuj0/aVYnY
WRg24Hj21ow6EMXNhQQD7vyLzsuJOt0Gbv4qG1FyLiDo+t2ZW8pUx5KtN3JBf9nV1uY91P96rSys
7RPmZuFkUdNsk7RWxk+TC4GtRXzfuxSd8VC/homzkksAnuwibgRKE8rY86qPi0Y7PzfoPoPzaq0m
N7YFaWjkREmB5bHJGVrqpXN57VjIKyaaX+fIFBwrwL6L0EcvQv5aJOYpIxZwfvTq3ijuZVCn2fje
wpM7nGBqNSUMpzizzqryTMkgxOt+w6NOgn/wYSFJ/auXts8sD2fvqfl1nXdux8cGvzVHfUMj7lHf
8QrWgIT2jSLibYloOvtN3why/22xvF39ILFivu8z4CMPz/ZkXK88F6SnvZUsjoDl29NQVAzhUe9o
ZXNfu3negBrMHMqUUpNS1gU7fBTw8djZMSK28p1g2oS1IBFYXExAhjtg7Jjs1JOEWC1uFTH2ygY8
t6qxqP+LehgFXUc+tF97eXnSRwMa08XJ9Z0Hu2yGcyWISR1UNC3YU4Zs6qmUw8WU0NvWWtSti0et
XH7aFvYfASxg354CSS/nL+sBFDunAHfLMSHOQxJw+/SrfvvwsTwnd0DZFrHmKUNc5O4b3w0Vr2/j
G8FqPcPqieGH6kUpxdqCxtsiH8G7Rlnpd4AzCg9I8/CFgFiMDncyKhF+yi4MgSed1VFUJQd0C8Om
frdoLzjn/zL499DRv8/4tU5S81Af4PIMuNafQUV+Ah8XSr/mnZjmzwjHpLlGwGY4A6vMfG2gFDjr
pgpkF0fNc1zQnZy7YnS7ZUkQxvmu1x7JyM+na1CJFRSliursR20Wwo2W57H6Edg5z4sZaRDDNhkC
C9prxWX8umAsO8ucHBsCYVLumzAa0uX9xgQhNmznxyDpYmSIN/K1uQFcPAhs5bAh1D08F8HSbi+n
1AG2CPxVoyOQLG8HPnlXAm2a/Cq+uwC7NydALvpM+H7aUzfs2ZLfnBOQ6X5DBOodqwy/WOQRXJv+
VSvaA6f+Zp7jK00Zxh+R8Mbcac44wMGlIklGxkyMzFS56VtiZBu8fwFMux7VThewajdSbBEP66aJ
DwZhAmED9dwBF7wmCGHUnHH6rhhlQh9fgs0A7NKD19JgaIvxNTCzG0XdcZpYTEdTMA2MwrBc131n
QhR2JbuBJCTRvrytD8UgryacZlFEKdm6hGPdJMGHwFCpc5GqKV0f4u4XwsfbLrXODGw3Web0q9Zm
9Fu0QJMBMZLJKH9AVwnuD4CO3WcnyQ/AXjFKmalffwqOuUNwlrcshRKaAz5BLAAVl6/+jw2/SdDj
cXRAW8UXAc4x7Cn+QvmNDnHma+wpMDh8tCpNkGhBfGvtIJ/JfMCCwC7bc1js0c2mtSYMndQO3wdK
dnk+WUAmcYyGuE0Wvi1KC/XJ+yaD6NNQ+JTT/B6WjvgSmKR2dRZkrJo4uK+utIPpEE1FRBhfiYC2
ywgHKtTE031w3aPg4b9ACAByftpThcsxio6RYa8A1FivuKrXkYWZG2Vux2B1YzatslAlB83iBXmW
U1i5qNcXT09mBuwVXHszlr4xYvThwSzYOoCSPGW6kNyCOIJt4rrxAAYVXVG4IOtSQABwhrwIKBsj
tCof8D0wqPOvrLVNUAUqwgXMduXxBiUZLXz24lLsA9hItYeN22B9Vvl2qz/ukY7eycFBUaxezh6q
EfBGfFV3K5rQi7vRaqJ0pOjjB/9TaZ7x8+gjJWfMHNuQhAz86nhmabc7KphTX+/xhSLpnKigvQ7Y
p5J+Fa5iHqplcVum5O+NkKkUYuWWjbmzDYUcsRHogUYsoMvb1LNsZd3/nuo+Fn+oeCgE+b5FlX7w
xNA1i1bW8w0+HrGcHK6L2RuMgUd0o2OyN/od2G/tyuUL9qCXkHb+VwIBwtXVIsNsKl7SfYhuM/hD
Pz/6M1guhto9FYNjzS7aCxL/oBorYgd5X0x6/f81AxyNSlhZDGtNqz2UF4XJkDwogKfkQuUfn5ig
dH4nSMNhOSsRwUNz3l7MIoz+cTlj8migUjMo96Bqm5SxIyR+i0l2xdukUYwghaAd6cNq4yQW2ZFS
1F9P2b39pVpbHSbwd4HozZtgDrVv34APwJd5l2waBJrgCwGkEzzAS9cUzqQ2r341nCD9fTG4rLiI
gCT9st3GVUrhkDdy10GzCOGuyw8eROJPTDNnGsgXDI2lDcR/b1zq5oI0I7cAK60grZOL9bT0y45g
EJ16CJtibtCFZ3GeZujNv6QmEESO07wsetpZ4Lk+gw+Xltxq9FhhSUpHFnDTkcdV5URK9DezPDr6
0bjmY7Xfc6tdGQGXO4iSkxy2UMW/uUxo3N7WL/9db+PuUoMhozGgqIFVVOaXf3R0JVgN/koblQFD
vRhjdo9JhbuivAtR6bjgOZz13EyZ9YJA8BOp6wRakZ+PfHb5JUt2bCnkqHGNYDsNkTuNj8PCg0qu
IDQptymZJRkajE9Of2l4Nm+97xCF8GseIL3zB0KmGS+knRlNsgK3GCpGmZT1OqyPQaJJ3omBA5yg
rt7mTxJAUEtE6LFxphm3whQREpm2hLyaj3u27rtH+OFz40WdYEzJerxvdYiYo6RNNVFQwAo1Tagi
qrcxxOKclngzN5h37xLVXaKpj4BqhMVQn72d+nMCFDYPXUht8uKVXTNNeGJgRl3vdWdl0NmdYLX+
8YE0C3vdXylVSsY68tv6Fe6A8T0arICf3WqqSV7wegv4XeAeR2ifTLx3WjT6WqAwN3mNEtfliD+F
Sxcv/RBwCmVhnLYwnG+9qHlkb29QyUdDgg0XYo2JSTiTl9tMSz6m1X0BBQNfiraIOoGbWFvz3Uzs
I7NOXy5QKyyB++7spoqjbm6RUZ0RWJdXINllYUqO/pYvgpbKlvGwK9MmXJkmA5eq8GFDBFN3LJ3F
mCzIQ3fGkYTsIQH81sQXu1EVidIefaoccxJI4NoZu65MqbMlQFjz3fch6EM26iAvIjWwrf122Ou2
JmCRkcRBoaGnTJFWOr0k+DsXH45rNhogHOSo0Lne169ATtfN9BNU8oCNSvTZXt73M2UR8qc+hUsA
9JjSoOHGIGpgNJI/BCFm/EM79C3l2x8G3PaSaIGjwj4Xtzr5iDQK+jwrXybCOjhC/KgYfUPDi3KJ
ZYFXTkhqPdocPXhTKIShYOpqmOWHo0nhSRtjo8i0AlfHCA5DQgQWJArUOxq/8vEtu4BqjclGxxXv
h/RdIXnNvfUx/wYmr+UBTBmBcSzw1POAuHMgUi5grJ4goMj3Cc20XjWr/+jY5TjbKi2JLgJeJWK4
XjzFABYCsJ8ZUuO/iABlKYWRCY2Kn8M+//k668yuxv5D0zow1TVS18lvwtTD+HwsOVcwyocAix6r
xvM5n+yWytm++H05Np9okhHIHwrBhuAl80d/M354L+/BaI3WxaOcuzNALKeFBtdofUbP9cP0UJbZ
SpgqQ4AtzI0ibliWG8OhNNMK3KmBHvYeVRLUeBWaB32NmW95DJ1HU1eGvwDwjiiENN1MY7tAOO5s
z9rxo8IIz8qK0yqSsp3BQVoJstVo6g4xz/2rPNaSlAW35RIQkNKKdnfbbQw5cGH+ehU48yBPmfxX
c3/wbZ5Yy0CeEXJnQmufxwIfy+8NZ7QsN28KkJBpYa65ea/s2ps7GbFmGM1xXSyGtmCZdH0nXipx
A3NKYejEDtcwMYs0NvXScsfTgYzknAkth9F4CdEi0l9s9EjCIZ4UASvvIt2OCWYP5gUx6nsNgVgK
9xD92H/HWgA/X9HygVQe1VrKTAguzAlyHC4LJFg3WhIVayrrYnbvlvUVw89YBfHhIzBBzpqTEy0Q
dfcIzDDG5K2HaiSO4E2dyz8MjDXn5+nqBU+z8Pvr5EDx+lPfjjyJom/J0RwnPnMGqDPBBOR2KvBn
mMtWE6nkUbRQvtNBRyhdlzYl4Th1krGhaT2OEnoJU4Ea0Wd4xOM0ALEANPpeacYIEraOC06f/StV
Jmr7cFOnp4hTy0NY/S8P93shQJh38x6cDcAbQ9Tvrhzqm2FUiMGsvh9Yjz6spLXMnd0U58W2eHvK
EqmN/MuO9WhjnROcLsU+x89hYKX2lO9IvywAyN4koHcP5xjPGWbEXng+3kHv+jqENWE/MiZ9rqlF
BCi7MVt4YiLwJa771nivm9g0kG5xWivr1Ee/GJ0x7xmWQzbEZ5a56avsNmRhffnJ2JwbNU/1NkMB
tK/0wOsaTt+sw9KmQ5IN6ivIwdtT7RVzbpiDxejiovZigVXHpQ/nJePAl3eyt5k72UGZho8vDKe2
8liRi8uBANLPXqiIdgZfBegfYNBhiXZS2KlPaBpoadb3jB/lYN6/kmtUjVD+G6l/E4LeiIEjxceD
akl/3ikVW5W8ASRLk+FnuyhEbpaP5WsMMTP9Ew00TUjQTRTetXYMYn3DOrm/r27pLrHibzRQ8XBj
Dttx/qAVl6JQBYYiQywMu/JP0EkQ7XMgcSb1YciRSmp2rQasAUhWYmDYIcnTLqbyfEp2a3Vtzvs/
SH50jns7lyLXIVbkS+Oc0AT52H2NqUC4MeOlQJMwtHmltIzp5iEiwX4fzSI7LQ7HwMS4PwjRYKQn
pvjEE62eyxkZYkLyxL2IVIEoTQnJozRyVnnsdbRL7W9RyRiO1um8IuSScwfv9Xqa2cIWtThgKSMZ
/rb60/6i83aDQ2bTNSECdwbesAM+zB80gBgtGsSKMPpcNxXmgiMbUPTNBwPOTMj/rbsYwUcP4f3a
W257R6jyQG3PPUc0L1+8xTTJN7G5lABjG4iJkWk2+VcjNWjUsblodwiH+gzGBhrqvj9OcVVXXUqp
mi8VVja0+AJQ/2lG+D9v49sOcwrXTqbZScEosyeGu+YfX49OzXREfyn1XNuOjgq6tfTGef6RH4ej
IQXv99oEmRIN3Equ1FjsodEW+ebiC9KLfXsOg3mA2C11uLUQC6C+cqofMLWgiZd1bROrHpXQGGAz
urIP1W5bit7LrlvycSrpM+bmzccFJKPeY9vIvnBg1Z4ERFr4VpRncOkgFqaTkweFYjHEkdgvXCTf
lrtlVZh5YJhRCDVvclfk4+JKmew0jyvLgHBcj/KfqVJ+duAncfR6s4a5SHt2IoW49vQ30oVvEjqd
6H5Ku6mImVhSSo0GLT1uLbm/gJpwqZnPDcIyvKuLXM3TjqlWyfRC159Zl8HgI1leQy9JVQzjTpJS
0Gyc+TtPhpjnoBlehFqcD8G7faYb3hQnU4DW5HaBA7lQG/hYLH9ZQLHLWby+fqKPQlrTbErTUi+l
zjQQh1Gmr1JAFMgY1LyVYrmslesQ7NfBN4JndZOZDidKSGoog4+loIPgsVdKSXfFFUNWj/ZIIIzJ
DJY+HfV5P11aFLa01MaljQYLivTl+gjZjJAvKC/HzJS0MnCrWoOlN+Z53ON/i3z1nmpiFK623Rkq
y0MRIHUf0dRpz+cfJPjftSvfACK5n6oEBM5OaQWBZ9vpPU2dWvdO/32il6yE8aKy8hcbxnHK9AAr
ZJqlmCI7fsUBLBIMEss8+Qc64PeuL9YBAZfTClcL717uWRH5gbXu9CGmEKHYbRFofgMn17siwxMi
WbjyZyRSzw+URo7SA4/y7CaIqKfdTzXetcR4c7J01r2qH6S/HSPZlOQ2XE+tF6bFy+NwNxmRAYcq
Bjg77t1wBCe3NCzq97OdL6qltMVDXNvsXKEnf7SYBzWsclp/G2oQ662aEuK6oHxTuoE6Xx/dEp3K
nGTRxhbllaENBDQp0ymlUM6w7hkTj9dgsq/nkucK01aUKst6OlOb3ITjUHYB8ScY9QUW2UAbpnR0
21tpwQFm5LtR1WDEBYtsCwIDW5paYx7qqmPS1RFewShl3efG2Oo9vrW6DKKaoXX901nV5CdVjuoS
7Nv+LuDOVEoZs5tygUXP4xmgkqbPVj+6dFHYC1jlD7oPxNeBq7JIp4SwzWqnsm5/S01PB9Lox7vn
33Bci1y6o8oYCic/DybaV5Z7LQHAM0TFDAR25a30DRrCHR7FTi8CLYqp8GjhFYyJQObwAGyzv+Z1
tj/y+yxrc1s4U/TWSAU4dVyBp5pEx4JLRHi5Zimq49H1VWDY7tpYNXBkLXSFls/6BnxReUFJ1F0q
xoILNpz3zg8Lm6rA1NtDQz+xBnZMyex4wqk34eUkmv++XgdEvai3y/o25X0SLYN95Ij6ZrPLdhxP
mOp8sTiOUYXOjYNrNpFaOJiFcuVwrXBG0OiRZty9DigISMbOItk4ClDM/1ZXxNVWTGb2EIzLUPMj
XbV0wJli5chVyNIEJgoVlp/iuTRSFvFsmES2fEyGpTp1eytKFaWGnAyjBASCcg68mkzsjr55iORA
uFQBNmZGvcJWO0pA3J84gubiVsSdam4f2U8PV6gcllegxU3AfDrso1gsg2NcIL3sPDPgESbn6sfZ
fhbWWHa1gkzaVd3MCjEIG2ve7/CFGM+OJJPD82M2ALDWcp2vOX9qkZoG9j9fscL/FcLbHEEqt90S
fsiDFk3pegpQ41KCBmUFifKjR5Kzex1BduOTi4GNSd+c/aB/T54A95gm/WHeAWi3BPf2QXWoJETi
M9d0X5bYaXQhRZAmWiivggMbjL7u2UEisRFttHUa23MsPA5xrBPISRye5Xt7gjoiurHbZ8KP8LUR
oVAPspiDZIx1PmdZoNRa4oZNCwrfvP8jUwOg02kU1AvSDUG1eyrkC/WOqOP7QB9I+Cr3o2zRwO7C
ixelwmG5HUVI0yUJbu3uRHivgnqQ5JxyRvrhoUzQdIPvPU8QLYnGbPKASYR97U5jg9urdjVNMfgN
xzZYbcWdBDfaoWVxs1inpPStma4z9YE30CNLagS5SnMFkc4Lxn518n++kWTW+btI8R0Ip5PQgPTw
NLWFBgzLh8FzZUJbJfWFlkEbIvLwBxzI6DPYfrNDrerP5gG0mPMRmdYWRbkC+X06nFR+TPb3MdgK
f8EJ22yNuPwdWqq2zgqwzOaAweLgCwQvVTczYbQk8iwR71rFi1AQkEjU12cNR9b6K0M6JQkEF+eI
MHusDgeWeN538TqLAghNGPWo46Rwdn0EnihFplc5NyiVv2/CTJj80nsXiwd/goRbo11T7PqanrDw
AQgt7Wax/FCBwY+aTXhpZ8U3UO+ClXt2pjzUiXU1/WYuaTEmjycGx0h8iM7hAYAEi/zqeLhI1Y3e
DyIudSDLIu5nipSzLgjLm+q5/hYh1/fk240nHDM0mN4x1WcOKyg3GSr3cACHgOdXFHngdoiNTSr7
aYtSeOuG1Z1KQtqmvOO6l1iG/K2+sedjcYfP1guWsKmv++hsOyXIUTjZ12HxGF7bIVRBcV6CK+wc
pHitwObRzmSOhMtw+Ty1jhSGiCvqn8QVAB+Q1DcVe/c4vAO47P7HDBUOoTXS8THENCMNM9KrRpWL
Nclze9HA3gXwfRv8D8g+FdL0hwsfD+zWkNKCCsMwxp8+r2EH7jtKAq5bZ2rr3+Dmg7hhyxT5FZM+
CtW/uMR5ONBEI4r1iI/tCKpRkWxpFZbXoRcqP84JyffbMSirwVVAZO1El3ROtCvtb04PjPdQQp6F
qxXu7GHBw6Y15hn1XdRtHscgI+hXjDXL0tg0ANmfLo++iqWdPzPTVg6Fn6+SQeGFpHZqTUXPYhBp
0B9FwT2MtOU7SwNTqQNQ9xNK6O2BUKti41HrQTk6Zbv5aNwSKbbMl+huUq7EYKA6fKyIc2GrPi+z
apGD068FphJ45bd4+0KuhOy2v0pdEdoElWdnXFeEZuHRRMdZkG9FSS2jEIeSj3kCLmp6wmtRVO9p
0wSxTUQZH/mZbEH9+Rmnmi5yUOBwqcUtnQZwvMwSC07I3h0OagGD9XDrD+2sUUk4Oj/RKLnqv5xT
LdNjUcG2Hl7cO/A4GPdjcvOHXWPNjTb3qdxj4bYxCl202TB2U1RigzizlSvKbY0OuZBcbqZJBqHN
cmu0lDES6DZFsB/aGW0afx1IiR2xgeKU0vqn3nWE0yj9eY6MKnkyqrKgS7dYKSRm8tsQC39Mk8mN
eQF7130EtiJUioTWuZP1ggB4Og6gwmK3546NLQonbV6ytlUZDwkaJobA5NSh5cBWG9AiPcTihXO+
mqn997/nGMTRWgXxkqrXQMLv8q6cd1mTliZyUBegHTWLtj7QxVF1nnyhML1k60IMQfiapx6cJzce
oEPJwAep0mMHecAsvMX1N5WhvfZ7Awff7qqFoSDsuUDRXELC0gQjvB2GL9ncUvh3AskggZxtSfeD
XSBVT+3VU2eyq6HTixEwgCGxAYE8ca/SXlEFGHxzyTfm4h+nobz8XlE7LH1HXQUF+ZAIyRRLBHG3
JKbDkZeDXUZtgNjjpgbYtfRZBSFwx7x+ywnJtM+L6GZxa8OjawXvPtdd9/jJPGKcJM/YoLNc3Ry/
J/msOwsGeAZraTDHQD3Mh+tJLJf6dLSXEiImpkH6dAog6Amixr/1C+4ybE46Sn5ouuaNBm3Cli0D
isHpIshnMNvDZgCQrplTW6ZMUyO9SkjvwrrQogjynNrtJ1feeEurCAGAtP8BkeLnMtbkqAsjrtlX
nKrklrm2Q6jKymyTsSnN/kILugIYh5RFg9rk+1LSWFFOoHnMiG98/A9o74YEZAbVr177Q8uPBZfp
zbeWLU2rtt+wvEOopz+B9an4fqhPlgbS1qvkJ53lez7A5JQqqbbehRlA73JFttmGZtcrITHCZKy6
4nYIkDn5EC4k9ZR3rNTRMf7dYxUWZmpQGQSjTA9eAgwe5qNA6KcOuT4edOeUs49LC9jsWyFKpyR4
8q6RknTwdPpBlNQtv+POvrVxn/0ayKOip+ImbDE3hDc/Shgc0iGuP1WollbVUGrNFRwCAjXGH1XU
82nocWffV4fYKRWr7JSs2LkYXyzurhdjGK9FfgjU6XMHAVJksNA7IpnN5+EsGJTXgl5PqsNQSynx
thmpKw/hfBaBLHK7f2wR2V8/sAwqPO3XB4MTParRnKkSaGEl4ApH/Fo0CVVvk16s4uh79Sap2DyG
0IfRt18OXZodpU9rgrSLeDvbzeRv9Y0KsUkrB15KSeumhYrtfCiCACasF+c2HyC7DVMDk75sTF19
iKhtv17u683CWovq3w8p8GBR3OL+XXSwSEIoswD8b78/+Z8nWltddiDWsFxx2w+WHcPyhoL+W6N7
C6fpbn5/eh/qsePGPbLCfTuIedfq9YlqezilvXrdYTsyi0h1+h0LldekJBDLxocNE8ldAqg5ugwC
Xt27X5kAmRY7wcKR0hnLVAwynxc/FZRDphuQsfQhtC/km5rKOPs4G2zBNM1uQ1XEh3e7aFKs8cDY
GIe9UGqNyF4xI6TANRMBUc+E6Ni5SFhn/xP4Zj5Y7iPqNCjDwUPRS5t1+mYh47Ah+6eHdGKIntnq
i1n9lXERMXYqqIwWaVmQqyC4y3Rs16qdqPtKZFhQI3VvSxnbFwbQhuJoSxocj8Bz7cVnUtb48OJ4
pPenMyi8jYc5vmg5oJVtok0qsFMvmbJo+DSNYgOK1/dOmqEuUjxpRKTAY4lpu8HtapstCfjWqV9+
9cu1ApPkwCfQUbCZWkqe4l7RUpeIhWNV9ABWgzdMAK8EvGFy93rEhXhzmaVgMvJVTFAdVEMi2aWe
9oM+qIHsqhsnosTvJg+tNQPg+ePrOwoP1NOHouPo87R6GMFcxZnM8zwuwOHKfdlpk79QxyYV7IGL
J98Et2W/RNu9oiNdxJpBwJJAnqW80s3AIWCbx8/B8j+MTHxADfkuO9pRvniDhy7ifcidQFEdffoA
wNGK0Q/IwQ1i4ThseLxCotyXJJ3ehn8JSFhSzBYaalFqELpe/EgSX0J6iedWTw+xcxJ4QF/CH+df
fFH2wcGEigBiAVGOPVpHu93+k+89AjXx7aixTrNe4YSrjoc1iGZJ8DmmYOPgSoydwqWG2BUKVrHf
6FBadOM5iKgP9EPKrhW2+oaxZP/g4UUiz12BSWDGo08PZ0/ARvv00yawaKHaG97X2ZYHdH9S3QEM
cxa1rt0K+0/SC1kLSySLNhy1+clFSqduORIw3vapvU2ZHlJrXwsw6NnRuR/9834GDTVedaFSGshi
FnnF+R2I1sSUuen/cSY/wDthIaFBI/FbgF6qeY4A2754Raj+WbDtEe7OgS35NlFMSrMZ7urWcIeS
+j2OqAAJv1Re+t5v/Cc4wcU1T5AQkaPynpEMfcHRXEK+ANi/tkZLmIkgX8jYl16FHNQNy8yK2A/b
r1/UJemG9SFqDT6ivr8u946iU2mG75/A5wQCJY/0zJfi8Ed0tNS6n3/H/V7I5mKtvOqeKpbauE/z
zCtsb4ihpZruwXhUGXebquKLW2VI/9xN5DH3fVDQWsrnOVKqEyNUnEj1iECRP66GF3APhp3xuLzJ
j9oUo+xuk+rxC+r+5FFqsdBAwRL4jF5pmr7tQf2BgTD93BQZOMUcRt/aaJlKhPTlQ9PfljTCUOYJ
ANYNU63m5LmnfxeZGGAu1Om6GfziHIOY7P6vvfjKUQrpnBxrHufIOAyDdAhQRVKAkCk8p32i7SSm
HOflG18ZRvv+7frgVkJSgkOQ60kr3i6SKELZn0Frgz1H1eOKl7oOfwmfalo8H01RL2qD1L/fhKVQ
TSNJ1Ay1slXMBgYb/F2zMVbRvWY79BIqZlKLD4FsV824YibLfta1xeN5Y3VQq7/WIFzldxa9a+Ok
BpaXw+EugXnKirox7/5zHyhydygc9FpXu6M4dOH+LVcbqe+Y+TV+lOnhNlrXb1gQxyecgPCIVFcQ
gbKDu9dqbcixo9bFQPcbpadie1GsUbfCtf2Xxj/wWbQodUY3eVSnM0vzucmd2s7CfpD3hGrJTP7l
ZW+jzd7xNr9O4ahu6Be63NbgdJ9cJmxsnWBTyTke3nsM8qj4qHyA8JPc93Fst6IAtOpqSFtP9Ke1
Sxstom2geNx1pbk7BmMl2d+aU5vOv5eUYhCV+jnz211UYIWNa7/hT7k4wkAhn2hdbo3IK4K/m3Pq
CKHTxZS2VLa95thzArmaJEHdM5GlB/3PnFSq452DNivFz9KcP5ctjLl4nVQ91vwXfC8tXc0SVhru
F0e7X8itK5uS8UjwzlizJSLYQhu9x0CaS/7O1GANsADTagqbsgSvH4GUnNufXhWMoTq+iJJCJc/w
bNVLWa9f22O8+JBuQOIkx+PNcxMu0UhNS/yZ91e8zFV9Mk8riV7WzrY8dXKD7vS2DrNzPakFF4hi
OJQOlaa3H3+AOEu+l2OBvsfRszAdP0S0wFNVfpdGxYnHWyKs0x/ANVxqP35YUK1S43p+Daxjh+Zn
OA8LODjvkAeKYDordwP3HjMeVKe4Y7EeVafHThKVpzHOAvbxcyRKu90Rmw7tG/ZK2Jhc+KIgT3O2
acWDZg5VvXVKG4Svczi+uwtwDrcDxH2R4LLBAOTVUaAgycBertHECu893cIS5cf/Mi4VD7UlCXLI
Bmy2cu1ZkX38w1D1e200t/BTl2N4zVqqt8GTPROpPRfSZYj9QIV59LTlQsWUY0xCVaCJ0aWFzEsf
NwieJs+NZHt4HGsLqICu7giC+AGtwOwlRGrhgTAnBtadQmC7h13RmpV8ZLVahxJED4Mq85sqczZR
Wh3OAY8CBF9/Njd4kQ+JTFR/JQb33+aFT8g9AOryip9s1afbc6XMNd90ATrEpUmcVcHUR8rSMihQ
y7fgHnUDT3pMSmoGmPx5bZUImdSSjb6xLVcUBXNF5tUZU/nTHfRGJLXlUUShkWIyaOqCv9990y+S
naxKEBaT3rB8183XKcpCjqaXIH+jceNgrVnJhOCFuU01CmBWA7pnR4EucGl49fB5Cd8fXgFCybB5
gfloHseJpwDiycs1o/QytJsm9YaQLuRnzD+wj4tXWUmoA1j7QrYAAqIEK42gzW6Y0nSAdpl08m/R
TZMFhzv8s4a+N+qxwS9G6/1XG85NR9xZ5NUMgkFlMlvHoXj3fS+jcUR1sC9msJllCTsaNduOXPHV
KizZLf6AlrcRN+czd51CM+LKArhPClF74vTptUJs4Sw9Wb5hWVW8uZzuz+UMollQk547g/4c8iKQ
w0RA18dUGRAleUbyoUuVBQH7AjGWo7qnAX3PXmbNTzCmAZ8AgXb/8TtYx6rH7B2Ei8cc+Ad4kM/H
NA36IqL5CMrZZNg2aJWUgFWkMOncSY1UoA0SOv7K2dbKkz6f6SGeSXaOwrZlOUbBfQYiBaHt7dUW
tbZJvp/5Rqk4+8ISdDUUoB2hKRLHvpJr0Kzhnc0zaHp0e9TCVmC4Yjs01s2pc/ESZw49b/UtahoJ
N2NHBHXNn41ZCjIGhRpP9cZGUiEMX2Xo30iXryuKO8yc0bj6qpVHIYurRZUyZey+4TEVDpV3WIaJ
fpyCUpx0HLfxsM6e41ypU3uN3FG4Dgb7OShXbGoBRgbOXcP1euoT2OiRX9fWJU1bsLrXcGf87EZ/
7lPIWBRFrIB8UBxbXYN+VyWi53B+l60B0aLubyyM+ofxcUtucNKw+I6j2TkuqLh66JH6zCpPxa2h
1oT1PM8tWKBG0ulkPxD8j3B8V/s3sNYLkumy34OesqxUqDPVdLoH4skClJvs/Q3R0+wwYBdjxi+5
/buojGph0RNk5oxu+OzvozQbzetHUzGWb/e48MfxmnMdO/Jbr6TdYWYCFb6yDgbq6D59SRc2wxOW
9CFm5yrB4eJG5ATIy2cz5AKFzE6kQnzh6qiL5O8EXGBoaV+RfJJgtgIqkPTqJ2JkJ9WAggYRm8uk
Y9uMw79XmN041PEc5KxZP+rXJ1VWEQBBdFQoFqakHWMdPZAZNg+j3vAvhVw4yFFSUmnw460gV2ry
i8daGAdK2LGhU6Vsh/wqiYFUBiKjolvohft89TmOKflpzWYWzSvVryiYXXLSQwk8vCkRsWitOnPv
sbD6RbhEGwfJVToj0YVLpzO4lQhPQw3V/bvaDgzsS9FmwIFb7LclxeB2Ck6ugHsUtVLDd2Cknupz
T5HAaOu2lkSP6clRuUxutS2sbCAcY4LlwmKsmlvPJTE08iVTfyX2LFb28aSr9eopU4gwSonPwsXj
jDB74QpYe4H2trm4NQ/H8MAKgjC07mFUweIwcpjsq5l1Ii8GltmRHayeMeDCsXnZTagHun3+26/3
NH4OGP4GBW9v2FFi8jWChK7Ulrq1UndImT4Zhpb/J0dVjdlMU0DdpHoUbPSwVk/fbrLANqVjxLrO
5Vkmjty7Srw7zWDLfqdXBc4YybzMyKiVxM60mumwslFfPWHyHEjFxKQxFaiOso8MvjIf7OK4Wo2T
a+vZ5TVVv88+af7Xk19Nc50gSL5hkxXqii7BGiZttckBfWbCuk6fHIe86G6ISv95CSed/XauE3eB
zbcDMMkBWia0TDig/cQTmz1fYH3HY0RzQdJQNTFLPeLAj0FHGfwJiN13/KpljdvCy17WNT8ZTtEE
hEsEXw9Y1AJ1rxwPUdknlC81Bk+gfQGZx72D1V8OBsLNwjx8DDzIwhpNJi0M858QV+NZX6LPnJNR
73Cr+ecS4fwPZ064bkhNNylj2ms+KVF4Cj5jR7CxS4TOdG2YCn+g7p+rB+/hK72YVj0ze2BeJQlU
S058Cw64wQiNY2ZYvGNwc3OJSofQ44A8ApeCGBYyfL1QxMSbR4AVC0qr7lR/qhGCJ3rEUvle1Dxi
JHd3cZsuK9isJucWIeK8U3b9V+nL23yHfuGam1q0Ic/nsikOACwVqYsW2SWX0i+2/x0qwQnqM7a9
2UFWLt5c9NkaQme8zHM9Bgd1auW83iT7WvyvGOTqFuBv5KMdTihb1tittjJmxaLoNTzwrjacdvmB
1FgxXIQgLImFnSlvyO2oJvf+2syjhfuKd1sPG2lud4YBfkJsNJcK4dKaOmAZtIb2ERuD4CkEUYiP
UQbCWF2muRFn5mVigJ5omZ18dMLKjYXy/Df56UyjpabT2UV6205U9FMgjRvtE+SEvlHV9Mc4eTjX
1SNPlShTOuFU0Z8tThelEzlF1OeZDIL2nUJxa8w7jUObHi2C48YQ4nz6VbyH+fZ/XWNDRbOg/F80
CFjJOy+rG34zv5K65OneiLUrtO9J6SJg5X9kxepbsPHYNanbRWfCN9llpnl/vu8kdH9HuTf23/FD
uMiUpxcAOSe5uUSUVRHR6F7pakI5xvEbCoaZm5utsXp0/Clm4lUam5KfqSL2oRKXNgjpEDvmYeEv
XZNBM7aV1VTUd7Jk5iOs1wvsxsYtMNFXRVbzfb5ZnoCMtqWILeOLn92lMrSauxa3W6INx21+xdPV
61Sy1zQmYL9WLWF0+hLfsMrRDoKVrq2XEDqQgtEWdcKMBfz1+MrHvzmpLkVC4AiXUOIZ1cy9px6D
Mk0bPwiaL8pcGKo3s89y3UgPLzaD92ddWvBmQaKDCMRmvJok7ugSneDfjzZPhKofxSt1jFmBBb78
MeR7BMCscvygL/MjklF0FUv9NecdxQh766qUM12QO/nhhQO800zPkf/BOtk30JuMPghBICYau9gE
VAoVbMpF2kCdyZaDHPwfrFnzNkdjSucpTP/q/5ieKqlMCoQQQB7mirH4Dyd3UhPwJzUtyxyxg2W/
Exguvh079i+dwjAMzmrEFQlJVVet8xXYBgrwrylGTXSSmsa49n8YHovKq/0Lt/9jCsYeBAvhMFdE
gU489lFoFHFEoiG0hj+wjNpW3cn4PShLw0Rtk+vpUkdNhu0xQcJk5OBeE2rg9yuqiBvGfxXlXBqd
bGgjwkVZZJB2wg1OGKHlqOnLFR3WQXVFw/DMpgw+DX/drg7pT1tL53CBffi5pGh0AY9l71gl6IGy
lafPd4MHzZMHtemAvti8631ed5vIubX625+2M1b9wtv6ogapq1TeV3y7oGOo9oodJqrnYRKtMsdV
bvYAZUDftGeM0jz4IjwEJBdtAe2eNXw3TclSV04a4j6ZI/lIDLijKPaAJgcaY0BsTvghQLU6Ybpk
jTwSG9OEVMHTdGp85lh9cCeRRRZslzB3SXJIXYgZdOQi/dxdL/N6K2lIZ3Sl56gvX0ab9xHirDGl
u1fsPVzZFLVah9L802qT0zhFp2FAGwXd4Hjt1zqJkCDeDjvKSSjy4+5ktnqsxoZujdn2K7mzMRny
aydSYttYrNCKBRWdOEbizLJCERg1/8t4XN7r3LwFx328Thv6xvDrVJCg9A2xZTokqUXCDosOC7wD
hnHQoLJSs7cgWBTyTdUpH0MdyPzcN0cSgxPVNqKGUOfPeHAo9KDlI/5SN8nY4tLEBuQGIWysjTEB
xow9S+65hdrpeIxEAyJXNyGsCvJgMnY43ZO5WN8h2ZvoWc9E5j/rxV/dGwzAUZQNbU02AXUnSB0g
El+lFf0Rq5ZF8Bljd6FHxaJ4iMxkYDA3H/ovXIA9Qa3KnE24bKyRnNbebJ74/lU4w1t5ilddPFw8
AX/1wzkXeWpgsshnf5LqH7aG3MoToeqkG4xiQUxzumMTqMm6SMEh7Enyti4MEX8I73ySywOZaJbD
3oB/ybM4ptCDHK1pDLxZYGD/hMjDu8tj1k6Fl4jb+sNfn3P9/amdmzeQ9gTeHT8ivGq5Ebn+6/N2
0dD1GXZMQykLqnXMs+8n9vvigW85u8dOLjY+ZP956EuUVo6R9C4d9fzLHNDypsvQ9Vu7BrIu/fow
TwIJg9EocXCnWK/W4TG1vj7iNYhrLxfe/jebB26/rNl478mKyB5CaIkjwAOV730V9D7TQGNtCM/N
c6RmeQJmJAb5CFKmMFhJxuobrqFTFzLFPRgdIQxBkpgvZTUYhZEZcWrho5E6NmSh7/LGUeDEBGj6
qrwJJ+KAGe0Wd3xK+OZ0meb8dJMM5zPeP6SxT6ZCG40u3lPYtwd7GoGvk4fozqK29AHKIkeg2Hoz
lZ1BNub9dBN90Ci3RIvfVm4wvdNCrRjoSRqdAExr560bJXiN0C35Rhbpzqj8knB1i4NAX3cJ2Zd9
LrfQiP2Ugvzcw4iv8VhH3xye8R/R4PSzeLW44G57Mhf4xs6qKFhMtP+FEO6Ajyzv0/FJdG0/5n4g
i0gNdQ8cpntu+MU1cj2D/ntl0P66VcIb7fa05GzxldOeVLAMPy1+MQxP7wtv/k6nvAchzub2Z6fK
OKONWaWRdTNcgbQ+o5Wr/olY74H5JgEl8jg/m0MB6syh/n6Op992fl8j4qwilvGBNky+xubsZ5Ta
S2C6KYGJ4tIj9LDsSeSR0liB5agg9nj1iGQI//ru3UOXDzZHh33sNEtbkKERouy+qKjvpaBcjGrU
kzI2RrplZdp/qyW0Cb0LN2nqSlS5hzIA5CXpYLrFMJ7JoMsPcb7seBnXPY1DpjnrYY/v0d2zDqDV
0t4bxiVen76n85pzi76v1eWw/MLTJuoN5UZjah8hk1Thez9QDiIANDSTrFFmTvXjXmDRg0x9U48K
glU1BMsv+0Sm/IHGuL/1+iePLey0gYr9+lL3Zgyd7r1hKKSyacKBKtwfL6e1EFtTESJP1gzhpwa+
mlxV/OmC1mbJKf3alF4FE8pWEt0CzQ6MWwQZVY+Wa9lMcqcXMWW6b5ximvbUDw/K08qIkq0Sm/ac
8SS+WWftJSbyUO3uBVb0T38v+Ue13z5pJ9oKhHrMyD5nNQ+D0Fuci7HqXtJc94t0EEaHWFWWx777
rbLkKGE9qoSgMyrvpo1Hbb/qitApPObIe5kiziOEUAQe2JHOIVzxuk4vhIE9cpWT9/5ctof+tyF4
ukxXImu3k0pw2IicZgbpHdGUpRwPbcbm8WYxYzJpIrLKZpXV1Oj/T23R9yROb8aWse3fbe9Tj3+s
VSCkYJbpG5Cx2tb2Q7aH+LRm5LC8s3khNtA2CN/AlvWAvyhZNpJ6BbNxpjmskA+yf5cdet3DuQoQ
NwhtJpRc5LQ2jrpMdMJXfS5khwFAQVgAsPWX5BS4/NCOqjuSul29UrQq0TZ+4oDgEGVpFpAWOXOQ
Vx5PDub8levbxvCW20KVbTHUVL/WX1dn9/VBErIJCu/1/wiIHjBqYO83Muw3KnBlcMze0sYY3pXf
pqgFdPK/FQcMmk+W32sGvCGzkX/R+NZgIjRTCK7sSPwjXkMSp3XJY5U5ic/RqxN4IYtXjjCM/XGL
Z6hIgt2HFsCPFZfytAU8ELnrOg/9Fzs3rVsyN6Yqn9q0CFTaFYMLNGyuMObOjE12q/1qkPwVU4nX
nZl81d5P9OWt6nIWEdneG1Ya2vUT8YyltU9XlwNAAS5RuEtgcwt4jq1dul5l3cKNbiazC/ciw+7c
jtRUUaYY7G0vHIMCbza3R1vn9dci0IfXs+KK8pdRwxqgYw1AXgzssv862C4rTYjdCqHpx23JYoA/
FJy9Nndl0pBGzHj7GgHfl59FfmWOWF/FQaScf6vriTpRwklBOt7AVUipm3kTBiXQ9uRHcuqigNYb
Q+lgRFUxcv+f1nKBGma2Xn3rNkiqzfI/y/AzTzJ/iYcfNF3A+vyaGGqv1GiYeB9G6jGGEgyqlOfN
bOLcMOflf2dwlr/ubFWgqvd/l+8kI9vpOJ8BLI9SQW0kQDd4U8KuvOhVYrFKaGSwJJBqxg42L0jT
vPaNwGSQncPI3t69Vo3uP2bVw38Mo/Vrkui9Z+RzgZZ7sQXEsBARuHMpfRA7jQbW23tncP9CI87P
awX7A5PPJSTazBwj9NYGXbkhfZI7x99IInTKhDr64qhbdU0aLwyfCcek+MZPkgRzra7Sut2YPbUD
RWj7AL9qEpq2KqD7WHR91kD7Gwc6s714NpzKf19k8CPI02HmQhr7ozM/lsvH5kacAhxQhjtb0uc6
15zvuVCy3PYRAu6KeSpf4WCLxyVkca7iPsabjVrnDZ0ypFpEe8EsUm+RUtNbzdAc1FhqmjOI9++Q
518gAaGbimuFDyvYj9mmsYG6cStogW7FuEoTuO3JGuYug2rYWtzm0efn+548Pxo+G5ErmHWbyZ0r
qeJhr410HUn9RULLBi2FOvyw8l/X/z5DTS6/dXJpFKfvtXX2rsegs+LS7XW8SE8/tTQIs2F/yTuu
G21ASVJp3E2krpXWfebQ8CoEKhIfcytXW4A+ncs7sHsQ6vHBj+ZxgjtWG7C9+8JxuRf+aaJzqE8k
lBxX0ttgIoNixsrcfeNh2ckCPdbpm1M6rJi4aSN+ufryljyBFu+oAIvMuOu7aphjTn8+7vxCj7O4
rI35pZhzCuNV58EAVLzXDEPDvqTA4Hv/rOuNsLknXSHKl7ugsNNYUuMnHjNwYLKjBF+G+9jBVeqK
onNBlIlpMSTznENFfoXwt0CvKKCxJC6+MtPy0tiHFqq+E8/kp41RejQ2Fus+3YkBQj+/cjTGCY66
q4P5pRZDzm298vURCZHa9OB8/iizzfuC91EgtQLjqROlWzWETyfCsTL/LUs5V3sxCYSIXhEl+KcN
89PhgmJ926iNASHrQ380oCh6H4PxhUtKrjkLLkSPiyXTcD/yHvhJqMIiP0iStGqmjjmG9LYqD5Rq
5wmHXZjwlPSPuvUL59ktVl7xXEKyCZiMrkR9BiFI6Sx8MagV6nAuPAWyQOyNq5F7duXt9aUtjuUv
iVK2sflMu3AyJr/SrPk4lbVGRIIKnZpvVuTGkD7z9h9bk+u5szLm3gMFH9M89XUhvZQkS98pye2H
bZUg+SF1pZLTIzO/7a3FNzqNzZz2WBxs58f2VgkTC2ytw0vswgE2uuCQUXuZY7h9x1PxCZ6T9Bxx
Br04F1WY/cMPAOPwRjtumTRNQJGnT3g+/KOyhTe6peUaP8+jYtzknV5J55Zm3yDWrkg1Pc3+9TRM
AtgI3BRZdlS3my09k/1S/PmQdBXiJNGa5JOHETRUwnYh43HnnagTFHbhMR9nyVFWAhzCAcSfwfPs
CrT45XkgXTg14OE0adBYkG+JDS9HHJ+NfbSfEjPWgg4yycxQIhzvBiTB9fW76Uqulv77fd55aC6Z
KsyNUdyvqMxZt2YawEUiUS2dU3Bnzyxnzyehc8yk6xGe8BPF306wpZsF4qZvlLaiTyr4vqA0jsKR
1ok7U1s7z68cnusRF+RGwLXdl2mwnZmyJLpkcsaA3xHf0XPRgAdnR65TszaydHZ/sRtq8PoJZTgL
w7DjaQFzc7yAqBrlN8IJ3dPnHMSOgwK63KoTxZAgjDxHwc65NoYxO3EUvP2jgJNw1gHzL/rKpZGp
bgDv+/Aef13C8eBeHAoTdoCMgJc652iN0+mjwyKqcYdZctWWBbtPe5euOL0H5ZMnPlgmDpCROpBu
QaWH7DBF8R2m9Scept+FvJVtIonPs5mffFP6Lu7YQhKoi33zEemUR2d7k6/huaw0N89on47ScNSA
8f+bpsAjnF50D2MiH+bV2anLUjGXEtNswWt1Iny5mrtX/yey3qHcPtYsf6K81g2UHZq3LEsr6MzV
8toIZOniR9eCxpa+K2zNTnoIco82DXl5Tz+ojKTJ9uL8oLbP6DjSt8zoWd0kbHXVYUL7ATmvAOXp
BkrOLqT1MOKJ/JXFy5PZ2VqIQIrThY17RuEm40IA8goI9c+Th/qmaFd1oDTLxOcHpyU41XQkmHDW
0o7Uck0ADfUVGEM8plOOkbgUGFHdxEhvgvH/rIVTSfja/43ahm6g0BzZfuVK2y2NTwmwK0YtwnyN
OYXNJOZ7uYPXMxE9Olp9Qp7ra2uc5uT7TBE2N0icf+ZUuan9fqea9otAEAeaxLN0SnAWVua/vQSj
LRJUHBAcelBxxCz4yQlBbcnMahbqKoVD4P2tmc8QEvSCDQwGxO3T3bZpNBgv3C+xh5hob+P+ifDm
eHV/PVr5+3eiZr/Q6aawYIFw8UIF6YukeF6BLFOrPPYLzfdWbUuN6qFMaOOpbZyj1TNaSfA1TlK/
L2cWXtgbsxX1U5gS3GdCPYe2AO8Rq0uelIejAa6zKGkBj09K13BUqxm7v/X2KzmxcI7MoKwrr7ch
VFy0U4i+TceQstvgQ8HwufEp8Pvy8eyMB8EyRSDzUX+MfQ45LQaNNcrWy8P7wZCV9qbEj57wi4H1
5RV/CwBGbOwUwDXscTXLR+a+6cVWC25LnUNVmyYKvaIbTUFYqXWsGWxnRKfvnM7UlQhO5RtMyxum
K/gIrauEJijuwoZ6+Kpc7CDFj992levr1a1Fs9Xkglj5kECbbVEJzG7RkewlvftOZ5JuhYk4MBa2
Si0/rHq1ViNZGEU4CTtjlEQlpxTP6zjkkQM8q9xy99m5rjU+CVGho/DUzOw/h5K2Yabxuza+IxIM
uxRcAmCqAJEJgvC3I+EXmlSGc/U6vID30n+0d8/C+Wxb2xCldPCveAWqsOBMVTb6tEksqYrFq1vh
guFEUlf5MhSZhRirTEA9rD+JKuuzBAnGOFZiSnyfQgD9lQ2NEn6F/74QRZHuNc038oWxWxkOPVx+
WthFYarzKZlysvBfZmaEn0ZAwupBwLlSKludw9tlCz7JAY7/c2cIV3X6JAhJnERWbfrwREBNPH3s
t8UoYHgHrSfyRzk1fTIlWEeYGPNx4aQQk0DlD3KWO3WGgt5N3egWE86q7UCM/ILT+MHuS4noZatu
CkMBBeKKoeo9y/QHk8ENPP3wK32Nb4Mrev03hSquNIUuLTBnx7fEHf3RsnKrYA9hynEOfe87ZEui
8oM2k2qOf4M4nA/F8/X/EcNKxgCyhXFKTXRJCAcWTQgYeDZOmEc0DeTukIwMGnaSo7j9ivKhR/Sq
G6pSXSp4Aaj75P5fO7HhVXMt7bjn3r3wTSkbgXhfAvbRw6KV/K33FrHh91VmZfMGqtSz2eslFZPq
YHTA4Da3G6CqOJnX7rTdH5uwei/8hXeU0Bd7zve8kQVPVcXynZ647A9YS2/kE1j3A/nOpaII1M0o
5FM7xPOWs/eXeD4W0JDS5Q6wijurMZOEZgq43dZzB8M+nIzqk81OKElX3F8uQpe0G4sOFizCD2hE
Hw5DudUXkBq2iadTua9XEJA7bfGm7c4DPLsKgCV61TERbh7aLoU0RIpkhe/6lD7a2KTkwMRx/9CR
CFUk/HnmL4U9ojBz0Y/czRwQ/GaQ1lB9wL03mIzeFM3ODV8td+u2egyb77JXwv/hW50pNdYa4kXv
s4LeyWVSrSIUxjp49XQAbKgBvrAAxGJpAtqdylf0yPST2+5qDqikYEfTscspgzskSO5ky0Dpm+y9
eKzXTChAX90/4yTnlwnPPWmx1VYkjT93XAeXaXpQKTn8ouTz6dI+nG9QK4P2A4cTdmUT5YuNGB6i
6O5LnRV1aowIBstzoCHL8/WkMjwENwHwpHlA0FXNXnp/J3gwN+JJD6fvMMVrCgkW3GXRZH0kDZf0
K+iQgGvlO+VRIbw8sBsNP/KgxMN91tqyePsc4P3pY2SV7z7VXj8hwLhV4avqcmyrcG7rg1yGN6m7
w93QAdsERjwGRzams6XAjcrJhaQ9Kr4zeNAsJSqhbui2dKGRNDFLM/zm/KyRnvlnYhbFKkMvMrPa
jowopfZS66keLz6AsbI83RtMZi6dhj5uj/sWOH3lLgQrPRhIV20N0UWcwkFBHsY4WXEWPb2b9One
8E95uV7FbZhCtEE8szSXQUo2PRidk53i5kScCcHT1Eto4Nsq9zgVQ2SWYGz9i+vwRVHuJ2RC95mQ
LrlU0p+jyk7bO+li2LSJpV/v/f8ZtNLof+CyD0UVu3BsCIl/CBF6axUSOKsLIfjpMxWmMV6qJ/0m
rRHU0fNH9qduUjmbkCPP6eE5WAt2vTyc6k0brvuWrUtm8xDxvroxOq4YPev4QvtWQ+Cmp2P6L/SC
MtjHr0WzqJ0Z/9FZC5jRBliyRINZjLJip+vKcEuF8QLFcawnt3+2tcY/14MqgOaHaa5xcSW3tm1E
wlQd0Lrbft0XODQKfhmJK4iIIeNQPRD+r+ZCUmL60PSKldquQRGvHI4WhOejiYVfoeF4qLD5mkjp
zhvXXP7umGSBtKK9E8vIQcIwAUwdN6bRcTomOIqnPeNeGC7AOlUsYkcMdJT1qjTKZYyquBcEAPYz
yxJab0kRiFmDrfLOaD1JujpfzyTXwmfSkSSsG/BzYoKwqqxxxBrGeOnJ+hDQvJjFx/ctAq+aMlSQ
cT9newCPxmUY/3TfyLlkzAfmGinVnXO/XnGqtHdSEFopnCSMpz3nD6s/6ppBDhaHckGWeef/qTp1
/QxGc3q1P1/61OesexkfMgdEHqEcx9FQpXeEv2tYJhBtUVH7Ijn6gtztLh2Csn91D7k94J+NGLM4
KkQ3IrcueavHv2LBpao3s5Vy/Xf/vT2zJMihhxS4PyL02LcbugMH3lSwMn0nwaRwZRKr5FJ+ak2b
bqHwRsfKuGa/Xr1Ei9mdicwCBN06g66U/42fL5b2liH0RXLD2V2DgCxxohYU7ZkHKhj7FnTml5od
sWcQbNIJAkjzhWsKePR0l2+/RuQ2wXZQqTAg28QEbNNuTPmMPk+DFyURw6SmkbRtyN3op1u9ald8
HiFuI1LVBwzPJYuDaeJ9s2Sbx4bE/aea7VY+joOeCQUR9EdFLnlkyAGmpOt7NNsJQ7witd4akV1Y
Qbk/XosCjRQS7bb3ScmutQJ8uAVSyUZGQ7LqU/szwee3XHdUnvl2h4hMPFySkFrDBI4s8sdYGbzm
h4YF2GO7IbXvQ/EhhSdd+0Y5PCUfXSHFCzOjFp4nI0XWTdM/nlv6+vGn9pB2HlQ8OTXUF3kz3JKh
IQVxw2dk4zOHVBntDbfSaTfFQaQHWAXE96SKl2jvU/c2Goon+RIOwRm7+R0Nvh37fhtsX8I06Tjo
PdL3d5lSIZTNhmkeV/rOMDMvk63T9m2JoL2XqxjBwurf5+IONYYHY2JWK8orc4xizgrQpycZBMse
EJVErSvSR+xjjHnlEx9u5g4OZlROtQGOCsYQf+jvHljWtE+G2Pi0WsEb32CFfCxF9mPXoKx/y8fj
HhB3AXT1Kzpsj2+uaEbytrbxu/c0/qGrr9xCAvnIdRkBNLdJP24YYICZxxhScxy/T2Ww1eUoDhS6
eHgkA2sBTGNtZWrQPFU0zjBQYBQt1H8/zTMYXVIatEDslKuQ/hTf3xIikZbk5HZIxeihsJhcjrC5
tLqr3wc6fmejRz+wRIYoKtlHlpe6pURQsyWs85daRt4wFSbjO2eCn9yMAL1Mj3Zr0Xv3ZSR+ON9L
A/ugamlYFp4SXOBowPNhR4oa4InOZW83rrkeKrI5JvsBS50tFIaN7fFzkZsInV31xIr7A4l2EqeE
FC4DIExnluZxC2xkqecfcdoYZmUxbyWOXD7epLWjFwuHfGrZ4s6q9hE0hiVqblpIn6OKNHAzvxWe
+0yGcybD1f9UE3GkY/NTtE17nM7JkArIIQmuqdAWEA4O8cfat3gIS9cI9aq8IRrEUI2G6P0iUBsS
QJOaF6LxRgtHRV5B4t7x9PXwnMj+6MT8zxThsGAxNlL1jtHqmPEL2stuCTp2Xxt1F2cSomaTE9TN
asIlc0RM0KvXAa5XLVCCQGirTw+4cNW4PbcQWgPaRTMol5TSop2IcKaWzSIMCzgZ6URfJ3yqn4iN
MJAUDIdSNMGMVhN6HnqoS+W7PSeLI1fdfGDgwL4P2n0YHQPcMU+r8W06bOP/9aW5gNpoxZiEpJq/
Oo6IL9hWbczxXbu1kjbfh09RwA2I3UM1JnV3YewgK9KskmxBSrFTyLhHEE2hgUWW0NdQ3rJnHmI3
l4mxrJeP/7zWvNiA9hzsiwJGiCrsegYoOV8gkszlf2Jwrb+07SIkJnKmvmV5NhLl84b6AZQTD2pH
0dqaYZNzvzG6Il3pmyiYNT+w89U2KADhQQ2wOfYuWW689HHG6ue2QiCGV1ePBOG+UGYMG3RWuqrb
lfns5ux9mnz1UAGM9Ijq/7eVnLZ4DCZ44BxaNlkW8a0qCXTPUdzgPWRekt4osVNSmRCqlonZYnE/
O950UznwUKhDIXvnpgwklT7tQSyrhRlrlkR03EwK4Xb6wn5BX5UdMQOJ2t6Z0RnD+dHNsDNcZSVA
taOTpoJiAmwiRbYVPcrOxSRyPZmSjFxBLJ88OFVGjTaFhFmZyLQiH3FBTHOj8mBcnQr3DDc2injz
IbDFMSdqEeIl5bqY9EPPI+jCeaM/y0h9Zrg2bSfC19J8pNSpHrfwbsC2xXrIeY4uNiA19ZLPN1JU
RGODh7ADafeyC52RcBTMvJPg/ujtsEfSzAt3i+Jj/z/jackdxymjzcEMXvDoJ2gdfGyKZk8Kv8SW
1QF35AO3y3jiLmrRoPkIH9YosrVQDQe+9lWnqYsyWe9v4hdh3Aw2W52t6ndEf4j8Zuynf4GB9z/7
8joz4kr7V5G+6zUEjZ2n5gJeAEUWg8VmecvFBCvb6VshMBCp3oS2OCuGgBQ3mBuThEWxA739LYpj
59Aieq9uaqSA51XSVwfzySMp5XiqtFu1kLe6PgURi/D77tSZkw4rL1wDQ6AZ47Ljf0kNVWVl3MLT
lZHstTvS2lX6w1uuOaKpGIQd9AYjOkdcxG87q98A28uY+se3PRsEpy/3dYp5NYtirvEWgHXS01+m
VpC1V8k2rIYldcjQMImHHS8d9aOVOEZFyNWvAEgRlLCrrDFMQLF2668F52Cw9Bq4mz4BSZ7DHu4v
Ygxw8WgCM3PlKHJBDuaf2FpZBV8P+Uh15PkENPmxQZtQ0XdTdPD1LpYCHeHk5nzK0YWBNvgHRScQ
ijeL4tpDnhOPacgd6+ezHkWB+Ow4eR/rWqeXy4HJ9nMX4x1amnmcCvbR0rypbz3B+svVkbgJozs3
kufKkqGid9Xqe7L3PyG9CIdvkUJW663I7AnryD5tLugHuBLshGgQzS2rCn07l96vz+bE3lD6h+H6
XPx5lC/qD9CWb/KIAmfC93K1FSm12Cwtk/x/edY3d4UjKSW8s8VHP3IH1c3a/chQpcWSdqYAXNVI
DkNpBh4qz8gKpbqHbhQ/M1yapTzWdyRFLoEnMQbgaezBS3XWgdbV7kODJXBM4ojjDhNdmBpPoT0h
Rc/99UjUfGAMTosemPdCAidI8GFg+XrErosW9QdFibuCpI9yjKWVPh+WjuFi/cLTj9GJyelMbH6G
3NI4YIYEmxWYaXe6bVc2MzqhF1L3npULRLI3cg/paIU5RrjVzfRiZz59eBomvHryZSEMIba6UQJd
JJMoelfNdKaXZo9XD834AAo+Ak1OQQIeV+R1ykBiOv0VzrxAnce8youafplwM4u+MUjRoVmkJbRV
Rf1yiG7GcjZzArQ6Y2uLrdPZwImoyXRbUOXhJ+phRk6xlgzIvWhVYG9r0w+Q0Pyx84y9kl+4UVj3
XP4H12wjWDJ33UnwOP9/m5Z3Di+7SS6dyFb34rl3SS86Keh866srrAmcVQFuUCEPR6s04hk3tl43
qykpMOFCjI+zP6x/+eGnImGU1T/V4Ml0W0ylR/j2xtY/Z64MsSfYqHWT7yHxWN5GcoJ65Bg35eBF
32I2JHNaPYul8x1DgSIUwRliTLiKYy+Koa7WlBKjcx3ea25mFTDvsz+yZ+D6JXVZTOOoMfrGjzbg
ZkMTxEDD6oFpHAlrpj2pYSoqhXQm/ayml//GBVJaVOR9ESQFpnYZiLCThBS+M9DkKoghUoTeOEPa
t8jyBg8lLPhOD+hFZ+V/Tb8HyYX/Fk7B/QH2/G7xpjI5sVyafXPIHkUYA8ERKV9QyBEru2xuTTDb
jrABAXxRZSqlzyw6n5DiDO28VYB1GNHtvTNzkpm14G737d4AtLyKYuloJlTcLa6QX1nurjtOG1h9
LEOBu0dCHFO25VZzyhpTwTnAIW6vCgOvS4188IyUnpqD+fNWEQSKVOUkZs1f8q/H3kigA0Ki9OVW
eWKAjvD16aJ496NEXJhmZ96q/O7dkPebl1ouD0SpbRG3DWWjJtJyO+cRfOuJWIYNf7adCfYh6qyn
xjpiaANUwKPsW4n3KFBXmvNqR1pjBUlL9wB8qQ37onzfYRYDMDQQa+/DQmUtcv7wRO1YbFgSFxc9
9TZJBRhI3PHpEgYpZmpsN/yWEXL5pRtEA8wZ1hD6EnQSptYNwAUnkuw1lC1oM7ADsg00gIs/FLL/
UOPKMZrT7mOHPClMih5ebp3fRTu3m3H6qBwTnNhLCnA7MGEqkyC8/gSKAjXs6i+PPbJYsh4Zd0xB
rTCYbjiyEV/hxfXtZJIA2RbGPq2Q9PVMgqYLixUjkpDRiaGIfgBydQHnu/Q356L20OHJkqJuPiwH
esNXZ2YnB4e14qC5YbbMoKHfLZqyeVwvZ3DFxdJMxT3wgng8uX9ScekYQWrJp1hYvKq3CqMSIiSm
o2bjvr3stN5GF4ISvP/dxBRkZ0q8BC2SB4wyPh+/M2zIt3T977xn7qNzZQjKVVrII7HN9jpVxpmO
0ueVGUnsZf6p86/Au9U1bBvWyjRNcFNUhAKgrOAk2BSR2Z3a1yxPuo6FrYMGpcuPS5nQbs9lD6kZ
4AsqHbiulmNhCiyb5U36A/FPsE0a66f0WXBneATOhfUGrb0d5KWQxhcQ7e84IBcZZOKFeIKV58nU
6RvqTTHzxDDQ9GX9WPzZwPQI5lCqspU3hL2NzCcv4W2a0wtSAlSYWzjAweqki09aAlQ07WxWZ4+o
qySrG5v6PLHpYOlDeZQCXLaIHyHlMhsYr+qkP490mxkJEbKDSZVs2bPi5O0Qp4egkkInU7CTLjY3
AkPmvwofvG9wo0JzccQ5e4jEg037Al6l9+SGuKK1H8rvQX449RIvHSevHidq3XGc9vdW3vqtKcD6
wSIkr4Bt75cnTCEc3funycgW3bbJnQIo7JNST9omN+hx885WVfwPYSr8E0O+cRKsgLoyfbI8gqQs
HXAYFcoMXU8wwXacGAlkJMsCHkENeJitIg+wBW74Xdnt0WDGyY31BpYc4mXFQohiYgwTMmeHoZgR
nmB4DJ9tSu0Nlww6sMVEdhoySC4uMR8rI0q3LjL0GLcIXmkLWL78nMfRCDnnjIxITqp1T6fE3RN7
TMTT6+6WAm2t+knkMMtGYOwtERxey0vb5qnF+vx17ZH/3Jpxo06tB8mn4mux0QL+uID5+3w7Hxut
EODe0bnWa4YKY2aJPEe9RghSEQ0r2cK5e0r3kEuIjmYar1VY/imVkyYh53XTM1YSaXTAYKShXqcI
vsn3BXVpGOuINcGtN3QejwQd8u9gror3t6nagvDf8FCXwpgJQ8wdZN9dBV6n+ioRoEopkoCrbpML
VMs97KMqEeoFm9MaQvtI4ozIEqY2ILlkJofmkgm3uqPzCJwTzEUH53VLYy4AYL8DONdAYJAos8nR
3/KWPfyOMBJZ1XbWcypbgCkBHMfbs/45+BRm28cB784VULgur9KSPJR++TnKnJkswBXNoVHcmjJK
egClzMDEyWgpiu/vtWOojfm5wOoMAEiDdWBNN1H9JHRQ/nNVhYcT2zuSStzxoAgzvch0sqiS9qOJ
8J4OQc/x9gjehLk7+/3ST194E/FqQAxGnzemhPtigJSD47JwZPxgrHrbXc6nfKOqT3YAtG5j/AXp
bue+5L6vMAwEHKwVuEqo7rONc95iHx7WmMK6Xng30rf78/+tmsZtelZGPO4dwaU0cX4aemXx7XD3
YNZJWe8NwymUyV57LPga9jubMoi4tM6mJugzM/8Hl9RsV8iX/P5H6rLNrD5Yu4qGT+jNUcHHvd8h
GDyGMMbR0vgs3ROL+xQOizu6bDrrSS2RVV+Kqs6QzVw2EnaEb20W6VS9rMj/d3/R6ntdgWK9rkaA
92EGnp1nVpIXEK98oWHrc995Nko9ksn8O6M3ZqGyAvZv3WjY7MsqCo7FA3W02T7sm/DkgAldYY49
iUiaEqUFxk8mUh42QLs5zNrMi41EDyx0rVReCTr0l54KI05o2J1QYx63Y4DX4INTxFQlgponNWGQ
GqS0PU8fmX4MtYvqQtfxyl22hq11ouB9NE8yebKH+OBjMRmK8XbLjKBi3EBXNqZTI66gC0Vf8gaR
MKnj3eDJxsn0dfS2AH+uyGETVwsl5xI/C5yWNK5ZpwTKIQQEycBgpKknT11J1QnNv4rfrY5aLVJY
eYqYs1YnAJYdBBWvNb5bxJkrpExyStAW0JujYD4sa95DGhjTWoa69rzYbAMplF0NdZso8aZAPtAy
bcrRUuKnf9OFJC/Q4w8CkhPvQIgSu/twlva6WME4FiRT2FTr1g2MSV5gI4+BwNMho7yFgt/WMN0c
lR0p2cmUXfKzDh797AnRUIiQEfNQp++uikGkTPLIqgi2ojUZIWC27jG1MHbCXoqz+NmwF1QtqWpS
itndk8TVeYK9QywGFOQ+LtyeMXVfi+Cuf7jFqIe3+qyavlFDcNCAdvI7zTcBvIKK8oZNCqHhtceC
lqgJsABqhsz10uN8lROUHGq2YKEUHfFLt/3uB+iKlMPPj4PMaXfdtpUos1LQS4gpVLrjJ60NrjFa
mv+H7rX/jNcHZRr73MfA18LhIFzi6gHFHfsoErGsaP0WHiPTh/+t1nEeWXav4/RpmlCSJzgg6+yi
l7qBxCZB3QFWQ3Fk8U4Kn5q1m6TVMg+ZhcYbo+ZnJIeWWiMZq5UbFMQD9y+PPhzgNpAT3LHpFXA3
70ipZr0HXV7fe3Cih7UWuWUcjSmCULUFUTnO1MH2K+FsdU0xqYjf0SMTGoYFNQ+IcwDBbl3x/rSk
24GeEhvJ472+iqksssTmYvI3ZPg6+10tzL20gz7GLZCtwdOOfdRi0o0bjMms9pn/rxNWyrN15KWM
rWinU7nlPocw31eC3d+VR0XEOmUusIiwC14CwmBN77inQJGdyW3PREcfGLdqn/Qv0f6Ifb7trNgf
fOtdqJWX71vgseBBkcXyKwpOIk85xJ6nJ+VWAbcw9pF0TBA1e4eOWuS6corH9yz7FglAnwTi4h3u
FIaF0zIIzXrnJgtY7P4cpnwLFGj1Vbjex7hyxSH8AVvL/p29Vz80F3CwYuYPKdY6eEvY76P6Bhlx
vghHk0ddp1mV3fOygsoGO+i+M6bouQZGp87pseMxP9iOkY1yzkBKtiSgIPSWcAimT6jR2L1cuDej
kBp8oWvkArVB0AKQzhX/lF39WY8D6DrYPm3BXUZrxNlk+CY5oiTQ2/09BTC+5fMB6qmabvVWnj7G
coIp7YVGN6zvuzBp/DKuWTCjB4OSNlo14wJCTg9wl5BSSDoymTq42DofcEgHuAGKL3ohIi39M7tZ
GUC+ggGukkH/t9fySrpz9IOUPjQi7t3w4Ibu/hLz2vJQt6sz7H/apzB9tpXJk7Fm3rddq0+nIAbe
/Owe5NLv5GSUwaDEuj69h8iVzZH3J0No3xH6sXoRWiDKi3YZ2AtIRucPoZw+tF1T9boE3JKyj93p
V9ex64E2WnVhIf4ExVQgeAP2ENIARhYaJHfTboZxNf58/XygZFPwjfJb77QzWeq6QkIWFEpi6MO9
AFec9h+LxdSu6+sWpX/jcNxnr1YgcPQAdlwILnY28agMp/dQGuZOnvLtGTCkzWwUc2rpUOLHT9Rc
vw4tJrYaO9aDVBeh4VrkVSGe2g2ZQE9gpmQ5gjHjB9WrDuNaYIunZxFQ6fBHiE74xiwchFYWFphP
jXXcVX6Pu6nNp7P2NsmEFoyk8i6EbOPPVxLAd3mep2h8PFYapvOHhz2BsZQ6TzYZ3Kh0BLgSBDhD
uLOxNbMN4Hrqbl/G6esXxg2nTg550+9yIjhIcZfmbb9Ey2GMJvb/Rz0fs4v5ivc23FltcDkyDMUW
WuCpEiSkDho2/gSxsMPkaduuN7KTdn6wFAlz7LWN0mmGBsXIc2dIbVb/gqsPeAb+1ddKwPg8+qpt
dz/5syBbRCrhvoKR9O98GPmwTcIqFvGxm/SsC/dlLmKjquXnnqnlyweGjXSBGttZs/IEmJHuhgdm
lBrC9KXuuD4v2FBT8PBqSzC4tpME4n5yLkyyKcMBnKUETkUB6XeXLF7R/kT25lqQYXo3h5jr45rT
UUiYlZmJCSdpWjh8tYisr3OCeAtNkl7uCOPx87Gj6KiHnbWUexE68BQ/YrnodzM7olZAt7zlHsg9
5yncXgMPs6B3i+WDKsNCsoxc5rIDnQ+wXXy7wMYVmnTUDcfBu9YjMdVpPtB4/ee8zjfumxRYgugs
lRX98DHfnfsgh6Yf33GyHlDnrn/JyrwIXpIwaHqTDlvInx59vkmYPlkxGnfFkducMqg3bgGJW9xr
qG4s9kF8IljKKQHckcX+lAqairCDq8qzz1ckrZ7ZBdK/djF4omgm/CtXW8vb6SDZtM1pQ1FI7aGN
EVKaOazNCG6GsuiqoKzHLT/8U88tKdDuMlJGsdler19JSs5gd8RbmZas+9pWgE3NmU3Ddc2L5CGI
syXu0Vm1knczG0cjNkN6F1Ta/RmHI1fIGUKNkxSt4tGa8T28RTtkqWh8F5gaUesZCFqSPw/aql64
T+FQwk1m2OdsUl3Js4GTBKdeyETeLFC03NQPaObxJk6AAGMKLghk3nPLERiJg99ligFS4RtbKljc
DKviXvZdrWOr5HXbF6rAWDYNZR2LeO/eaFsoR/SbnOL8vP1IxngbhRlqdEAFAKjv1UALXkP2uBiS
XgU0xz2ymqbp8Lu2nO6mIcketfhutTgmFiZH24F0/JabGPTye9WU8La9CXMKTphf3mPs4iOXDo4w
kuLSCm63xEbURX2DEKDYKe6VBwRe/qIojHMRmfrXGHVBugwb6RskAzsnOuJlgfVv6wF2SHRwtd26
+2g2h2jBD8aCPLXwp9Ig0nZMhug/mseMNN4hRBwSLCk+Fv/CdWT9tzw1nnn/3FJ8uZf0CQb0AJfG
zJ7J9DbgplCOMpgWy8xHE71MQEpx15uQnwKO+ydU3CaVj55f6Y161TC9ERzzW9WJiLE4sINed2Vq
O+XQw0l+mS3TOaSs+D2QoIxqzwc/Eq1EP2N3ipwpYmNsrnfpxqymGXqBMbMYAJ/aS04HNasMLpdJ
oOfFHF26RQ2zaNGk/GKg3VAzhTWchmffNlCEPo01J9VEor1Cb0yPNPnt9tLUVXYmpFu76g0004D5
eMK1rxd8VQYvDL9onuaX6Laxz5WwSm4yGN/lNwfZbiI7H45CGWjUF/j4ot7gDOi5X1PZNG4hCGAG
c3NfhkkZ1sblgTmlDsNYr75AnMtAvLLVmDds5U0mXsm/ljR5RRzoQCeBkOYcRWWfFT1sR/Q/5GsC
ExtdhWH8e/oVex93JmKwKGMy5nyuXaz3Q/sEaQa/aNK5gI5Ic/pTauEm/RsgA1ESwG2plAByO4KI
HLiq13eT+ljoDHRBgmu4EmfBmOxOydrFJyrxEMUWD1c/YpzOynyOKreHeS0jG5GH5zNgdAvj5/CM
RG6LD2I3s41RAs1CdT2HrQCadaHwdF4c5hf8qWUPrCgXKmUnPMmc4v/eFcdNuvBm7FWUfj+qtMnK
rpjsf0K3E0s+Bb2hNyRIlnmHusbQIRgrCMQ5Dvm9iFumhib2xzwcbFIvOsOfB/CJ9bd+OzZDSB4G
AnMMlQV9a51Y/feLONFJNmthNfrTAHFJip4kEGXZt/6BACSHft76Mc8K0VT1gtgO/DgDFEfpyFwR
psgbipY4yHNVK1M9w8hzSHLyhkHdnAv+/5FcnfkcTkGffMRq2f9jmq1519bQWFXmCWy+/ys5A+hz
wt2bTAFG+kaX/YYixk1cnsTKiZ0bm5kenYYKxTJh+untqROmajf6/kvMvDC30FgRfL7hu/ZtcFc7
cDX4oSIcMFvE2U27kk519PWNagJtsjT+bfvQCzDIcAzperQDPFfg/IJq4nnpOtcYQU78RgTLg6Or
Hnqf8GJPwkN4tWKNEB0c8fzhnm8xJg8nTyDLTff3ay4jM1IaBgjVF4xWupUt+lcOa+Z8Xho3AtIo
OaIy1kOfbFpn59HXsdbek7MzyO5Mg5KICmGtQtgfXuV0KPjp+aQ7RNb7AU1kiAZWEuExgD0DF/QY
lovbaCSWdKioiJLcE4Z3s5dSFOCAQ1C3N0T+T7wI3Ix1XJ3sn3iuE8bBm0/Zlz7F4438PUAOzUEh
kByDxZC+uTwcaZ6TQAOgjJ2SLUfDAj7Yv6LcKz/3Br6Eq3uRlp82++BLFK3LpyeiA7wJxibpAlUy
J3ei1PC/C+Ygi27/dBzLxQV8mSmUng5Ih4EOCmiG3KQ99ws7l5w6CfvotwPL2goDm/fEVlTW1E1x
ZxIlEjJzQQo17ANxaMygdWOoHweI3Ijb6JD5RmL1bC+BMy7N+4CJEnZiK2YokojEb/nXicEv6JsC
z4hYjv/ESTcI+Zbd/c4dYdPChxf41jnCmwmgPeufgliSNkqGmBvZ8J3a9zahujOmCCW7ytpvjpLk
bz0degfxBaIcjPAYQJ39EcJanEIROoEVb1ESoSYd8IF4JzHKUowiKxNIn2FwOOUfSRgZSgBH6pNH
HNMGKExyd/hevaJkHdjYkAP2iCYsp7LAAvXzV4YGdq+bV2hnTeNVWTpSO2ekxmIPXn/85c+pon4p
/VZpwbjantK3JnKGA7+o5YZZPplkwyaiGOh3g1/EienL5WBr9lz/iUz0CGgT82TCHrSGS/IQmTAN
nR86dEFM7q8Jf4tPTZjjw4WFlFxyqJ8LuEgqLioOVMbyxBY5/79dtDdjn6a9KcBq1NYBeplW0bqs
H6mV1T8Y4v8b2paFMNuv/2uX/SD8wffifTjtN2XzzYnKcBMprz3/OCi+CR192+HdaaDzQIxdIYJM
EykcGuMvWMV4ns0CCe9L24c5DFnAziiRiEHCpGWMHbQru0C2iKCvuLR/Ifk2u1tI61Yyn7eTjdZB
+OB5o4RuKK88gSTZjerNss1CMG/ptYO32LyUZOAmNYPELj5Yhz8K0SZwD6jLLzeOIyiQV8gPKke5
kISuCQs5U341yly48BCQnqzWwy/q5fwQZ0oo46pVCN4se8DeCHm7EPSdDNaBLCunDskkVJ4qIwFr
Xvt+O3WvcTiW05QfV86aqNoIlYN7x3broQ+hvx7QsKSB0nlKjKrh/JqagiOCzW41wkoX4ZdsjoWU
J5gDUabfdpnhmd6AdSWhiDgHeuZcTe/HX9ZjqhX+2oUIlH0eU8vkc2wlT7m7XuR6BShFjJc945Fl
zAZTIzbsWiRMj0tUHgvG4bUyXhBsRuKwuiCo8YjGOguYng4gyF30uJ0u/23WphOCSQS0/t522v4y
Zef64HEbKV9jyY+UdeiJBnJhNjSMRomHguNHpgWQMkyfYrdjiGTduERDvkssf+z2SeyO/Stg+aFs
34awujn9qhQ2iILGbyBRTqJWC0SZSU84ub/9SMyIXU3r/AE8mJm2hOzqn18BT5yxUgTD4WgCwPZV
a35/S8sZpoChr0IdsrqA2wSDZqQZqttZ6pHMFi4N/gaQBkQDTRs4FAxTxJzP1TZm3DIXkvZsJ2Lg
D2YFQthcz2N+oRrr0WAJxwzB8c+F3gKjGU1SIfbXI2O678PLlFcp4GvNlc4o7f0WjfCsmINS9h31
7J1QbvMFm0xgc6zxd2eLMHBnoOqKDNdEZZZTOHa1tzgrussxtj/xRoR5wrVV+iFmn8f7/+MbElLn
0VWqiwvaAF+fj65ZG+8dAMsy/egKXet/a6qgWhI3Iq+OqtiG9VLetxRBeUrV2jRdru2b9zyxcAIa
vJ2E/q5j1nrsSk33VOl0M9Qbki59oVqvHm1AOPWVRrpiy7fBFzMsVDQzR9tEFqRAtJf7+XhIr837
jA7kSPggPOvdgSVqWQqCCWtJguT/YuEvleOHTNPnc6mg70jybyzephPE0/IclwsumsN2ZWO1r/uo
qZToFNNCoCXug6Rlso6IpBC4xdTWFGxtx+zRiWUjnuTK1322c+YkJ1AbRWFiBrQ5OQLbE537Uai3
dScUoJ9/A2BeuO86DL/VU3T4+OSS0K0RmdURh40Pbr8NIJjvU5xIhkpGbDnoMsJ50Fvs2VsELTFe
bXKCmYLzFI8D6rR8YmVYezTcVRlhzHz5GJP6XDRjaDGAgq8sbtYz94k7Q5Ce76N5R5cs0Fh3UeoA
S3Wf9Ah0E6lOfLHhnAaYkylQiGBneU9UmklDQezM4ztw4u0XReuSYdvB+w7EbRnJHSwM/l1jVu+j
BiZBZKMYEe6WRnGdFiKQH1MXobUHNANRj18CBDjrvJz/CC1jg4dhYDwxrmWFIIC7v8pfr7rMbSii
Knugyq1BWqtf85MfXq3Yff2BKNiFAmbeDxfdi4Vligwawg+4FFei0F5wYQYJBJu6hk2YcT2MsQ7/
3D6Rw+bS+LTA6Fye9isnCHWoH6O/2PVCIzG5QMH/ynPSohGloS3hgAjLwOQ/BvJJ/j3tyd3IUICy
LbpdnKNXqqPw+pCMC+LNr9ux9UUyw40tfX2uZN1/E4ytKi9EZ/m4Y/t30yy3wvqA5rg/X2k7IXLZ
wCwNS6KscM0Im1VJy5ZMi/VMBI1E+QJj/fxgiqPKjaJBdk67BWINRA087TrVRwTQsqGa1LpAxBlu
tGlVp5gNiofeMsB3irPh0GFt/N/B1qgfcHWEQl0vGR8ACRMrjlHjYajnQ/GPI0VuHDs0ejTwllDQ
DrD28nmk8iIEI3gyanBVEy/Der0zvbRxQAn46lsi9tRDvepPY4HKrZAZTFZith+N8L/zTchT4t5b
YqSYZJer1UdywcXf5Vq56j3t9mpljkXac4/pBQfkw/U6Xxt2tSCCcwueIeeixyz+SmDoX5qe/Qdk
7gITqc30QAxc+zM1uxBkt+j5fQHjsB/QWnAgLg5byG5TQg6ucxLP2O+wp9LnPLF9fQe6UbkbA4VL
OctzvMeH97cN8ZytkWSHkh8Y0IsU57641A02EYS1yOzsX5kZ2zoW2YE0F2dh0CLxGmIjXL8uEEyV
a44Yq0yS0/vDQd9FZCN+i7uxrKYF2jjEA+gO+L+UrDZvXAai3NE1cW3A/1VB7p+5nV7xvEIvAvB/
xSrCwb8M/0rlZERwdv1HaeJwOtPBt2by5Q9mwjVVpDBpcMt0tLu9ABFd0lYinqmmRBC5DCv5/SBp
dsEgF4rErOlHBM6FLXpnma81SkoKQG67wkrg3XZJ36SmAam/w3f90YIcNCrNn7gy5imly5DUfNCv
hrTrjFhjSHMD7wBveQtOtYaard8euh3CydkFVjn52aJWTv/mC9A72PwncPswmYVQSozsNyDb/2QW
QmhTG6XEYyBnfFQPbCsdzfr0sa31vCDnfUOVpvLyd1d4thTGQJ+x1wZpWc0hcmtT3Y6Bh/oFOO+Y
9cGkiWMby/4zcUHGzYjD3cMjLyduB33SWerNbXJAYw806X3Sj6ImcPDvgvwZrafcevDYxRmMcWTH
aYEgggkvziDmfYsPxGR5/688tB6IFutSYnT9ixvX800rg/D8yYwvVGKPccbQST151saxpO0S+CUE
0RyGCGe97ejJVkGEs6IIa7dZbyJoL33BOC51fNX9u6JiYY0nDzzpduLCIecag4ffK+G75n2c6uJY
pLn8XEDo6LSrv6gsi2bmIGdmbRyYaEmqyZ+ByERkWHTh2suVAEKlGavTZviUkG0lphe1zasFH/8L
KGHJiDgkNuqpUTXDhykTBmTnE4zGNR0kiNcpgAm9PpVRSx/DrtabF315X0a2egN5/G6GqX2ZScGS
jMXusw5km2Q9dpI3IVbRX0znd0qGh5Y8TxpFpufPbWYEuPDnRNbZa4An9ZO/P1hGjPDr1fAlfe5z
DyK0zJBm3TfJcigDzpJM6kqEewl6KKS/K23YBwm6fWdhz5bJ/hofS0CzA550zeeuMiE2O+vIAhjI
p5dITEcMAXY6H/+Z8jttU6LpvdIxJZoNGG5bW7pO4jBsZmfAg+z7NUY5O11XenV/+wClWu5X8/fG
evlULbJtNzVxdoacn1+f5zLmvwQzwOAvezjxaSeZQpvXkiaQLMntrX4aH0wIUkKRIoBbHnQE8+Cz
yK4Lw022glhx1/UuMROKJp5x7L81SQtDZf8xeZbpchQ6B4o6v73GjUlGPE5lHa4PKnWKuOb5n3/N
m+t+Q1BGZhgzMQeIG0sWlfMujQr2jVV0gFz19HWY0bTHpmNAXpZIyLWFh8MmuLMEqqCq36fyQnzR
1FBItwJa6crNfBuh0Pn79ZzZQfDFIC38Mx173EtaayS/zvxYYSmOoub5GI2LC8/o/a0PxU9co5Ny
FnL2uozpHptkQw1peaxOzV+vQ4lRTw9Pq7pI9FryflmF6ORRhmK4b0bzU4deAjXJaz+ud8g72s5r
xlTm5lu0WlZhzxTbwgfdq05Fk3+fyQ+AcXBV0bV1yZUs0EN2j4pRUEhHxo+AuMY7EhDAFnvZA1on
bcbtBvWcCd/GDjVQhAGGVVl9kjcM8vTQnk5nAe4+Xzl11xbOum1CUkDtmoImeMDCblY+DQxy1fqx
AMM+PUGwqR1NnodRX9aNj5u3Z9wc5NkryYYX9yASYAJ1LOcnPpuyjOUiedIbcvFeYokS12loyEd4
Ee5+wyF3eczJVk/6/BVMgFZrVxwVO04j7mYbZrfPPX15ig88LcvErzEttEJG13NesBF+BYz5rqGf
q1hwuzR61M3Eq849Kt0EC1Rcynh07VdBNiFdINaj6wdV5hDa87o2qn+VQTwM2N9z0F9FBpm+DdrL
mvvmI+8jrWqcafx3j9Xnp6yd68HXWLpIvwnUdg3WesQjFICc0m6b0HEQFXctmHfQqMSvOyh4Y6UU
DCHboZagYEtQpg5/dfJOznzSE+A/6HD+R4P3VmLcYJZ7YdLVmuPCgv1q6+/r2Wi1pFh84SQ/+lr4
ooyuIZYvBzQeA8UL161N08rvp0RqUuwMBL8SExqcSCXbuPqmgTcOKolQ/9BUZoDNwNkLHXh32fIk
3JKXUcKuh8IhEXypXLnWmIuqCduRLl+5x5YHXIVy9V9dqPQhbLF+x43ie0y239JNLR4JfnMXM10z
7ENX0A3Id4UNjG0FQE+JfeibCZUs/i6NGyTcqhEJuWsMaTHaU4Xug/EBKUXe17g421byjqywaPnI
W9VJJYnGpmP7zoGKYzr5/00kPbB7Zh7S3qlXbYW9A8edFpW8rLNAn2GEN1N698aCnXSE1ngCRP4G
/4HHqYGMiJknEhTeDYs87B83pmI8bPaR0rSPcU0o3bOMnTp4CDNejb5VscwC2PQM1h1NuCXY9eg4
t66Xb+qUg0h+YWsVArETyl7TGiqiYRXr3qN4If3QGCp3ugup2cf748Y8KAC8KWsmb2e1gT7aOgTq
0X6r0m7sMstKe3SyJMbhVKxvYqPEYzcxKXFRjvcOVoHSK/oRn6SXQl8I9VrT2rWd/EVBEiEw85+v
XLkQuBeHpWcZTkmT6ZYOoyVAdI9JUUS6I3ybkcO84UuDsCcTd/i7IAN36QKQfuG0NN38o1wDPT9j
QAGk9T5P4SDok7JS489ZOFHWglOHZ7xHNNzvFqbD+RD0BjKuCQJOu/Gl27qnd/r0yPSDi+rKmqfT
thftXpcrfFHIWpk27FRKh+LGH+mFCrN/lhRw3LePEiptzcGkXS2J768UE3HciHUek2XLJ+EjMIWK
TOdQ2VSC89zTqBRDzN0UXhRFOO0Eo5uZXgOKSq9dUkUxxVkY2I9g2WurodJrMHGSvR46jsxDpCK8
6d8tpaDtNPO736P/+zo3zGGvaamwnZVnzzYfkxrHAy4Tk13cF9lGWKSzsRwrwhbrLZOBXOuqotPz
FZWKgxTFiYcmzjnvtZtFufElq1A37vDQ8yaYUDK3cjNAGuud7XC98oJm9g4jV1iPzQ/DruEHYF04
oIMoxcD0t0BnRnu31BO/uzMLja2C35hdA/i2s5o8ftWZW5O/rZP9kkQgkqxZ+29M8nSDLuPmfs29
Y6eV38lb+M9AKnYwqYYusNoL0PXhAXXUvC7J+LLUgPnkW4ynTTHBvUOpLZ+qiVdh7HtAsEAnh9ZW
c9+6Cl2waPfzJyYa4sccqIcHGH8YQJU8Ot6nhl8E1v2fUr2PF5LawdWLforUF62cu/chmePS47az
89iPY1VlS7ZLN2Bp2fWWasZN1PoyslimmkAvn0150Zk8J3I+qQbL1vld3Xo3e6vto0a5fJrabHxy
4Y0DpNWuKdqkTr7oVvyQltXnRR2/UuzwvMQQt6eK5Uue9DvKO6LfrfQzPkKIWooWfPLdYtD0MvaE
DDRRPuPphsBAH48hJt3JtCcSky4S8gB/mYhcnEAMrPH/IKLXfoiRMOYCm+rs+ebtIvsf/810muhV
+11xVq+eY3i3QStIVYMax1MYjjRoQ23/XFOv5xnESRwo5+F8/6BlJuqR4tQyK8JIJu16qQ0w5jOj
fNfXyLS31ueVg/1cKVJzW106F8nJwKaWKMcIE9O5WfC6M3xPogmki89M5n9OrJADeUpX75MllZRS
DRJKdCsxRlhzs77OjXS3ioRBMoPN+4aCe/clZojk9bNoFZGifUL2AS3dFn5Ke6Iio3ctSRICwZQC
5L5hVFE7NKoah+qFKFg68+wCqIwM/aysBRdGasrPQrydyIfCHVhXAI3ImC8FBEmd1SQ/im3tThTt
WLZqwcgtFQdPMkJvkNyhPUUoaM6qUEpSfKjB7VQweIDb9+koAaGsJLsgkyK+NfcRCbFJOS8lO5HZ
AwsqPVz5c7rQncn58ZYWd+AZELXKJB+IN8ejl827np5DbFktnsIDlJBlnuq/N9M8bGxRtjuGakvY
ELl8vlBWwjgV6izpvMJVpZrOo0FpWhxdV+3pUAuPRUYUrc/bHR83oTsnQ6vh2+Hvu3DnlCbVx65l
AClhIxXtG/LrFfAHUe7X7IJyQ8g0FSYww5+h6Qq8Q3/ukXrkEVenKFJaQ6kg1W3H7zSg/ONNTneI
W0BXc2JV2NZPZGRdkOv9QHItdQaFbqCY/SzoE+sq33+qTCGeHcAN+ib40Ck2XJ1BP//lLKL7xIvV
2nRYn4xk+7TWulnvqJSIdphvJvNeUOe3YW8BrnrSCvPRSlFbOevZF54Th4W9slmvBxXzb3duqyG5
coJty4lS3ArCzhaoxdJuE0Uh0Gd/4txkAzQjUeQKuO1GtsUY5BB5NmVulo8al+coIy90Fadir1Qr
zvMdptsiMivAUI6Zpv9SHp+vBKXEy7omxurDNBIcz5Ddk0FWD0pu2cX6pIm1Mr6CAqlDDvjEVag6
E2bSJLbRqEcHr13R447WsKLPphggjLh1K/oMaWa6EYge6p0PFKb8J1xsEBv0Ykrc1obR+16kC4Hm
aqd8oJw15kpfvNau+iQjmrrAvOrP2K0CslgsSxoVfcTQofOPJZCSiDfuWGfS9qU26ZO2iiArQbw0
nVXT4pQjw6JlqviLYAhM76k9H+sszLVP22ishCdvQ5yxYbMZHV9w9r6P1CH7rVBRh8AnLldQ4C+r
J8H61a19NL21JMk67EyM7L2ylgCMaoXSowDJ0ZNqNZjZtNFJzpIHwTyCAaBjvgjBtOV3WkyCuDVA
TrsnR6xNRbT8qNSzeJuF/8AipqZQtuLRO6ztAHpdETAy4q7FZL6j5LjbWAxlFFYFC9L3r2Co9jrE
HUpuBWaW9hzr6WH5jtLvuZg/Bt51q2t5z5FNCjvqv5yCPkM0N4zMDK5nV8ltMj8qiITGNWT7AloI
nkWheNl1bCnQBcXDO0dEpSTTSofn4EdSvpFpvZanjVmQP9UvIjw4BelgpFPwqIkCDUE3T4k8OZhS
McCyLsz52VN/OYcP99BWHrAXwmMbaTHsczJiVLI3BF5e+aSUQyt1uKxT2fCBktb2eiXav0LoQ03e
ZqFakJoG22U2QfXaltIbKpSazX7oW1yAKXpT6XKImMFGVgE80k6btthl1POMRr41Nbg4z6pMfORU
0yugAzR+W7QIlFO6V7OfC+LqbfOgVrmRM5roKfBU+o8S4b1+aGRNeIYK1l/wUyd6t69ycPQUu6dL
Kmzn+R1t7C+B0suSepE3lUJc9SJSxCuUIbNKhOHdLSAj7ozSk9mkQfkSN985KpQRIaCGuQicvWuR
xKtnVsQnC4OiVdAEA8d+4+GukzSLa12u7yUn2l16miT3P2TvNqmWn6EQwT/xV+tk96lV3mK10/qe
dLOhp0e6BbqvXimvSYf9pU4fH6etSpIxfZruNXiLHSpx3fSCY8SnilsACwKS4ij1lyWUZIx+dfxp
dNnExXc2boIup48pMYuRMV7bJwSRB5LuuM9ctVfXWecRgELAbO3i4ec4iBI56cSSNUkG9zJ6R8P5
oDEwS3PBYJMVMxbEPKPfC/tJHiudKBuE6EiVjV8oZACIR3CccfZSxN/8gNMoM7o21IbpfqBW3Hmh
keFylvbS3I0Z/wBhtfYuLDvYVLLxlPr+q3fA1m1b95Uvxz9X6LXOx7RQRTuPyg8WdOTfZNMzEWcF
nSF49Z0RlUJYsL0ld7gwNmft+zI8eEs3umPYnhHalCFVyn3by5X/NGfOY+CGicUoQwHlNkZq8vVs
d5ixoPhK08pxpTE3g7fVIfrL21o8X4+vKpXzVdBxEoN3SuxPOhQDFlXZF3K1GSB6JdR9JFdZJJC3
nF5g5mEO5zy3JEgf7JL80kPXg8i5gxLMSMLG5K6wO+ZQgwcU2IOWhTL1pu5sx8e3dWcI6OkSsvTI
RiO8Le5CL7hq0f6fEBEmoSep3/UMXPw5PglajtlCU7PpSxobiKawmhUKDW9Bo6SIzds5H4sRiKoy
3QCWdtHkZncZqvC3tYCFpeSfspF0W2LgBINzw1J4X6p2ineUN1I+TYdUkyjrtJuhNXhiu+hPWmmQ
NWS1FVI1h7pX4dm/THIQhbKdh2aMEY0kaIOUAGYC5/3qyXrtSK1NRW/RHId9z5iitfvE4bZ1i3bz
dCmzOtu9UM2NTQj+p3WxKgwptT5WHytUow3c+YuR+A1lRma6W5EYGH1HZoUAjLh+DAjrVdho3nXt
xHO18RHt3ilQQiS4yA4SCRsZkiGnTlDxabKNLpkIpf2iYezWnXvwy8vPheVaHUmz6vVMRd859IeV
7GN0c4l+YI2DrVXw18JoDT0JZlC+eO/JswrSH6fiaEBOjB9wRfn9b0eM8Gcg10b2Kpo6pB2F3Pxs
em+hwT1qjeaDQfUAv4+j8SqiRgshgk95jehJZEaJlgnwva7xqveBLOwxxR6OHvwlacOeKLmqmbRC
OdJDPRt47ArY6la1GjE9fG/utiM1AVjhlOWqya2PDBuIpGucv1Uh8K4FQlW56ZML+j1c33/Fr2hn
6Ae3vZRXKCk7923iVRI1dBnx5PHy4HwOXszNPN5gR44v1BpeNpZkSsQp1uItWusz1LcLBjq2pjuw
g5DxLr+3SEEtqodhD7xVLgAW/ZdKg0HGABAhSxHFVtOgWIq7wmWFQIYlwydjXFmCLll1hVv5K2dg
0ubJTjx40q1ax3zZDORv90Md4OJbI9yTJfgifSy7sp4OG7cN7flyyj55w88ITXQpUlwNfoSmxMSs
7eQYzUF7kD2sPIZDI+e2+l+OHGYQYh3mwP1cz+SwjMD7iwAlR3nlM3Twyg3GDIq87hG0Qssss1El
kv49593vr8P9sRcACraPnCbMBgHYKFHbWsnfVC9/7ZIYhQycmmgwP2JOxA2QzElplf6t7A7pGWQm
9kdkPApxt13O29ANpCUU57USBIlAhX1oFlMfFD97yIwdgm7DzhiQdFKWbSa+EyAziS5oCfNnAZZw
mTJiMJu3AKj8qLyCRgrXqWCZFtZjtRAshswm1CFqMpbbZv5KsXwV8KxTvSOKc5wFsYEuDID6qRpY
Nlvwn5GI9dKls/zFdPD8GqS3CYW+/92kYq2unyitXj32Q9rm5ye7H61J/fnqXlw36PCQOTh5vm2S
wmKPADtD/dKsrLOEVoOPaM2j2IRg7gSQ0+VFSrJlMZSTeL+A9cE0HyVcNB72FHiIxPCyDJUW0XVd
dQXf5//tW4kfkvoEfIEie53RwHn/CFKtlzeelifran9mn31R37HW2xARAD51Rvw0MfnDi6qmki3B
gSu2cyNjbTQ1QrxBRzS6uY3t5HeMaxCMVGMvryJaAboXTtkmz2DLYICtLoehQ1Ec1fhhrISqssdI
woYpVUq/nOAdxCHjdFU2PcTxKPmW4Rpk/7dxh34cv5eUTmMQ5F2hPY9BT3c1tr9Y0sSRgDWBUAv+
QvewRpk9cF8grko18lWnKl7ZFVaDJFq45DPzUjvdLh2jZFX55w5N6FXCsqflZir7f5TU5zKDVnpR
Qhk5T4+Y3QLSEjz+EdyDEAMFZpGj4pWdb1paLryE8YuKU/wehjgu4tnt41pQsEZHV7MPiUx2Yvp9
btKjFvPJRKNrqOPYmvJi3aQw0xU5mYpqNGvedNOhCd3mUsv5DdRKpzihBFtbBW9Q1RGKOOtpb/l2
euQ4eV7WkftGrRboFdBjKTBj1iR1dzwxHvejWFzXGasBvP4l0q7cwVurCTzXx2iw8Cg1m5+APgPe
xHTXp3onRjylqnLbsRYHZtdN3mH1fgozAFj+SUYWD58jd2XA4geBlQjcMSATUegHPsku21XaZpeD
7DyOb9diyOM7aZTfH+xkv7lEJt5FxJuw2M+cmReZRzR3Ujm6hLXQmL1ljw4jVrf69FTry2ES2UR/
RvToEa1P20GnsI/j/uMTBZOBsSqg7nCastX5W9gFYoWa1txRY7/Xk45kCs5MdiG8blZTGJeWY1u5
wLeORb7yjvezuOLjw5aa6qBNoITHWQdr6mC+CS/Sc23k3ezqTb6rJPeRvBHmfsWEAUOgYdjDNwCV
u6pdtFm/TYmPsu8gKKyVQwveDfRUgnwnhKIcO6NrqCDPeXMOCNSZD4ct0C0laP668POt4QAq+0mi
sPAbedWnLJw/y7eU6kcw/PBkGQj8Au0pZdMVjNKcIw/uy9+NpSJ4BIlkP92kEa1+ZCcNLOrJcCES
TOFKHmwFvsdN/Yvp/c3K6GelsOuNXrtdbuMR9fnEB4bK0Zv885OZRGyLk7p1YONkE3t0VCGIN8dJ
rSMjZ9Obft2Z9uZAoXdH9+jJd8zeoPbJpXZWRZG+LhtkZnCfM7d4DBXRa0j+uh4BHlmSo128zZiO
SsA1VrpFPiquN/z+wWrZ74+0wgZ0cfZDr2hkZXvvMl8hDqf42wd+P28TE74lO5J2id8jFfhG2zdM
Un3D5Eotqumr1P727qqVv+2nO/KPNbf1T2V/0i6M6N4PrLa0cL//Vf/uNuD5CCcE/pXjo8GD+h6G
/ZFhrduCjQxNXnfx+FFSM/I23Z3+PbwnRmiP5iOm1fns4dgXEEjBJCLnYhi2DMlHVdd8//yblZ6M
9ZCoUNL0+Spibl4qv3gLkKougllwm7OV32o63Chw0JbmJmxen0JUTvDYrcLcpAjXaumK7NpCJv66
5EqVoGzj2gTyaCUMHiLV8U8R8pqKjp4hX8Cxb7vJFE3ePJfmbza6lDL99TPgAc/EkAIPGGVIz/EJ
QCTTG0qSbikDLAk58Vwt4nkiz7mcu76V3Ze6iZrs4yMbYgHh0BZ8D7f3iWLmRqlbp4a+Sfss4znq
zkMcQOo6sT6+vlsMM66QptfF6jwP99aqgqUWWp3iG6T0yvwdHn5ckCrEvRNpxOTRkY4XsOc6wtno
5EMHa6JMHGvECrkyP1Wc90nCA+L/Tb/wGZplxCKGu9hmpL9P7FjROA91e3Zh/ynrb0EZRw1QUcx9
8TFMKXZJxssyDPyWRJFQwXUpg8zpdX0/Ou1FmVc7u+ZpuqkrKLFn9R4bwVy0yaMUGRIQx9oqwtjI
35RukwKb37+2h11KRs3uR4sLw6YW4FQ6BDsQVl2+yBwkTkVq6BvRuNTtjg3ao9PPJoAtNhuS1jMM
8RNoNrFmQUeF1Q27qob2iXWJJWEC51f+p4c8YbM5DZ0OlSZIJZo/WpT80ElHHNrWcj5UvJH3+PCG
+kDMf11YQJIR+73UM4v03xDJ6odcVIzV2YMPciIyqGvAtasjh1R4zgQ4WjoxvIBpntAZCd2qrEP7
m0VXBFBgPj4C4dBYT3sWIyVi/rgCgVELDpNaf5/ZaU3hd+HJRYOOvxFlZYeVfRw40JRF37WLhrM7
Ga/48jB+3YN6W0AAmy0Tf8d07bxc59ua09TGICQ8Z+fUKmt83uDHjtbtR1eK0JZrnd6yiznHuqJB
C+6nq/lwnLEeaRpeE0ZnqEvLA6BItnL5yp6QeYijETga/NS4FEcdj0iLwN4Pnur3Jm5WLGUxq3rJ
j6IlQ5Z9494RijkyScnXzWw1IDMZlBsCBGs4J9j8pjqajV72ZjuEsUA76eKwIEnN9WuZjyRTMqns
ZYNPfiORGlvjMtz55YI7tKUuq1RpC2Uv/1Wz+ZTMdz18eS0fuePtALBk9AvNFRkM3py86PH0MRj4
uZZrxCzA9sP02hANVFsOoNM9gLCiU6nW7AJ8OWPKofsWBoZKeG5ehqYbAa7hNZutGLC/jN0d2cpi
Nw1vJuw0fPH2TPRWKyk2UJCGJ5zerM8ue0NPh+djjom3mZP2+EKEzH+GImJ2m/s2fsVfhPxX1Rqa
pSC7N4YRK4ypy8kW6INIAEp9oMF7pCiEhN0FNtwENTXX/JapWoEXZ/n134GljMIZ4B6fzHnpqtKs
L9QLyFc+2NTFTnjbiwH2qkOSELfaS4lSUZzr+aLg0tdFjX7f6miplfL6rgn9ov0yCmLnZvsyuylg
CSEIk8BkH1gQ8XeG9VtlXpxEhsOsO6WQj1PSDxhrRi/N0w2GUpdqwOc4VXwjQ3WMVqWrHpS64M+K
RxGQVOivY1/I6VmWqjJoTRkokSlAXZmSUeebV8w4CSz3cuU8vlXZQR6ny6YDK1L+OcXQeY1kPu8+
trUDv9Vh3d9a1vrpny3RLTSfkeC4FY6Sf27eRvHDKIYiAeV6z2MHWlcrNmTrPsx1pzdv/yhzGljx
2CJteo580zZVEyfapB1K/pKdOZMgrSaZc0Xz++dQ2lnsR5qdnsYEDj+jGI4Hp9bNThZ2njpIYoFO
9jDucfi5sGZ8iSx7rtFv0zmBujIRaY/ePZcv0grOmqADaCeDtxjyz/HrvmwXdnM74tZWCLWgtlQ/
7r+gZDwtjOIDm2kMmQqfthj+bavgjE6VmMP5Q2pUU1KK4WhHdV8Z60gwdRhtA2DRQwzcD9Jw3yQZ
AAEDtFzAqJQ8wdVBTQ0zq/ZxnsyqINLs0+y1HvRjdVQfcGSQJlILrNtQPTX+k+WPPdOnW2A9+fZt
+BAg7nUNePoCi91oIyBG7PDS+R72wlMn8jZBefk9fjac/A9NWp782H+OFrJa5ljDYZvNlU6K2Uqg
FYG+W1hU+BtulTl3UDo770Qc0AcC4CX9pDZF77Y3PtAmFEHAvLO3+RhTvjkUw+WqDFBNUdkJObq/
dTGQqMwsoJXMNrbfo8T51HV6j8YbwegGx29PoFAR6lEZrmv6ot0mh58YcRatx11k0VB8rxjPM4Wn
F2AbLAK/bfxXG1/AntXGiG8tHg9oQiZQzP0+i7n3TqrUIhh2IbG++lxclkcBmdBqELBfMbdfroYF
K6oNSl4iH9ZDjTMQaFXIKV1bj8n0e5Kmy7ApcDvOsyAXjBKEUG+uCYhn7Xl6gfNFp0xIQIDCOxAh
0R5NCdUYHxgtD3eG+HwCpkKGhNlmf+tMltd+vTi5FQKKYyLUbfy3H82y2YBYWY14rya//05B94Hl
zl57uCSe6GoRL0usumq/bO7V6zNmHC2vD93bYfsIY9eFtmbR1H9xtFxzSvexpdWh18GQ8zkt4kLh
uJQ1bNyv9z6xxstn+/65X5fwaxvXrQke/kP84D1jx7wFDsBbwE1qJApyDkcOAh0DnO2l0oqsnmD5
6igXzwnD6l7gZGq9+IL9YOAclSjVweMEduPhq1I6xj+JfE6pKv26b5UMKgwpiV+VMOTWIUDgLicB
sDLjHU1LIX6PxnkEq9iCnDq2N+46cQ/ApK/d8Tnb8BgyPPFqODp9lyofm+W6LjXeMvmIuSLpoDDr
EIIpQvJMUQQ8dTZ6HDmH0iJ7Ho1edXQwvvjF+f+oiyd0Sq4UipivzDMG5JZlOXToLKNOGF9Dq2SF
xboY16B3ARaaE4abiR6HndfYmRtHGWRZjMiEsdM599+Mxsbgqzc7nhj7SlKwazc/ohpjE+ozaT15
/B5JAEzbm2E0ToPfwWMfcGDaYygZ+uZIUiuL3MykcrT6Zs0T/rzzWCLctx13kgHHdP/ZrXma+omS
1iciB5sTVUUuYAfPLNHyAbYEx8trFj8Ap5s1pFkT64DzzFN6ZXww2cLBlaHrIb7e38p5ZZyUPXyO
rK85Vss7EFl76si7jmdRjGge/2snxa6vc7RMoCXZk+G4YgZ4zsq8aejNu0dxxaofpLC68wmcfvKQ
LLbID3NOFx3+tVX9M128M92zh3FixtTqBnvxDvp2nh1VuUuBWmJ4mP2TRYK3FH7CSCa6S74L28F0
2a2BNE/ki9XzOdGkxbZmcz00fUyFe6hNdrkeiixPb0NQK+F1Sn/eUc4DyJn1jCWYMFfrBg2u6vKa
yl4PsWw0XPwgR/2NWFojXwiEt00/BckkJm9i3Unu/1QvGg+sDL77WOBTAW4JQhRMMi7W4aVFM42N
uN2XYKET/Z+YgH7hOYIAOhfLX6XU7bF06aJ6leStpNmGxDXOVzlVtah+NcTrWUIyrUy5r3jrZEvz
/AgrWdG1+1gKy3vMJOO0I9Ti5bY1CkS0tRIiRouYYwl4M/hGIp30pe8L/dOKhm1EXyp406iVcfqU
afG+xZU1ZAZuLTvtkPj+/QHNQGv+IYBNNr5rRlVxwSULKZAA7OlsEwGUCXK8ZJgw92DEIMrPGM75
oZd9hF+VNyha7bzb69uZXjgPwoppgRlehZ2CIUVn3axONy7hvt80zK2KAhvPg5gfsMfkBK17vLpD
CRcX2Uh8LTpuMjX0moWmXKVa7BEITyitWJEuJDJzYvCRKaWcDG/mDniI6IFRZsAdNoK7zVyByk4e
SHWt5AJvoNW3nGprbHZq3Eo6LdU2UBfuoDIdPeGLQkFJSG/1pgwBkuC5FMEplNhscenC6oNtk92H
GBMxIQ6hDEuzSwHRIhHIWQ3Z7BOpTn/nC+n2oAufxDh423tF6ZW6/NHGGFYwrM1PnB5MWAjfhcmB
WAgPZWaCO3UYuL+fvmOVQY+mkHBDpZ7SraZ8nsMU4OOcypQBFHsRXBi9QSqa0h/QJUBp+Sn9npRX
ey//qMi3yQremfTqK18PMbRcIyF6/r/FVJDsdWJz0k1lyWxzOV7tiem3PPAvVLu1IPF4YJCQa1IU
2aJpJeKL7eRuTldSq1LRCvZm59I3FmP9lyeu1cLlzzN7DAV+wsqa7F/Rlsx+pecpNQcJcWwt1WHo
isnK2zRhxXCUUaHScKVzinE03AmYrOSklDjdLjwIsB0xPM875FdibvYd3fUwSkFe2JsEMCO2omaU
m59QksQdbot6I2SCHxcxrN+ob13LqGBNkEHx63/8Sz2eqV9yO2aTfPpDmxJdvblsjhqYorigm1xz
W2Z+n+eWnEWjsk3Gxt40yGAlfPaEFr0q/VIARJcZq+2Uvim3kbowHAYBHxZeoeCNVKXWsjpLy0IU
IBfeKV9v1zFTflQsYdArjwhReDuPqcpn+tZcctqHe0Si+isSYK9fWzrs4UxDSrhNkyecNR7ZLvv5
9EAUK8YH62vh6TsIb3vv+Ic+mspGLA3xVjJxm8UABQ+y+8tsMtTD1fqFEIqZpLjx3BgC9cmk72un
S9zOkqKm2OMIFd70grZHhjDcAajJWTt8FVMzowXEl7MZWNB4TjGlejpbWchZZVdz1PDyCBPmjsMn
WfNdoOiMCadDRL0DPKNAr2Zk+/D8IlVQeeLkBXXgSSEXz3SF11EMUONAZsuqNr6i5Iog9KLhsxEm
fuAFNi1XNKoKe8dHV1S2wtj3NUQ9xA87Db4OppwYTSFHNrIfcL1BfQE6CG9JWq8TenpRLmg1WlUt
Vyen+KECKLxGA3Wh+Tb7166rb5aXBCYK9+qHDQXV1+af3nDvzA9Q9/uaetQYJ90GT4Za2v2hG0Gd
WZQVxGY4j24nTAaC75wFm2RAmKSPmZcdTjKvMjmnBVWXlFX7ZEELlDnnM7KT1MIJd2EA0jTXunJl
R6cQ/wv442VAZxORID7SL8VDCiX/o6frJhVTCYTZoSgHfuATgO7BOFPkuqTv655NiUmSeySGm4+E
890Hpovx4ClAVxit1WzvYeNRdU/YBePqPZDfi2nwl9QYmKUBKSvYeemftcYZs+Y/n5zu8LuyYok+
Ch3+Ys4cV007tbOlBbIhB/d/c3nSMWwnpf/XbGUbdCgGKu5KJTogfVJJJpN3yVMqQ411303NULD7
oDKrAJybrEnWHPNYuskYRkpcgygwxsQ9f8eKCQoYf37KP9GvVc9zUCYvLlhFW5n6MGKK9pL+pnfw
ry6jyI6R7XOarYxlJZiQCisbInHrbzFurujMpYijCDVmTmRFiFEbhXByBDcs4xD6AxyYlVBQus5M
sULIeFfwSQ1XIPzogDYKSE19TcD1QW8dWneV2CjTiFLmkkbirV3gMq5IzKsPZCItj/bs/ZUrDq31
amuYjyjBVLivWWABH701v+32hGKNCbDn2yr1Ixc+Cm556WnYsBZDeSuAbfo1jo1PWW3s9ThdeVxQ
HkqqgPrGUqhw8gQwSKmzY0s+wTgujZu2M7y2pTBQY8x2cggUair5UThZXuZF6lx4/s2s6CsFwY5u
8vBk/cvHiH+iatdYTuoTu+02sdhRNxnABZWnF4USkMyjdC0M5gWcduodNqh/l25u6789/4FT+PA4
5/oTOsTNscfE3Z6DesZAfYOL302P+AKfidE9K1KzXbhK5o9vYC0vh9jh7tV2ImSFW4v0c9NIsEzn
La3wFSvIad4U9X6BdrW3nAfEIqWARARHDkQGvuv2l6v9XnVyA6muylnVAazHBOdu9aKRe+E6Dpgf
m32SYLoJOMH9FriARunVZyTXinvBU3/cqUi7xr6/CF4tvo1HY+lRSXaU23HBQOyKUV9XuhyMMYWK
bfpSlCegxYRxywZkWNCjXH6EtZEY8v9htXIGIpKmknSyFT4MxUZtgEgQIFvbwnDbrg718NThIPdm
QVxR1/XxKkj/jTPkF3G/Ukwjekzo+WhERnOKjTOXAG2G4DrkNawACMVN7ndhUCfQhLQ2ln3dUwhK
BqxlHE1KOaaLGKo7wQB2TEWOtpTi2SIhOT/lo5OfVO7nnsYRGFQ0/Ws6SdonPEAvlamcuiti1smf
QdE5buGg3NVGfxrdydCc/IujuI1jShY003MqeHfy9HJ1ies06L+Wl1TbMvqmOVjRmFBvUK3z8SbK
Wmpk9THLdqNxOiTAYhTd0t6ZVYCd8fPruL8VVj/KhNhhnf32zL+cgwoRbeaV6JQ0QWxY0M/cVW4V
+v/nmMotmd0qaOvQRlhLeG71Dj64dI5+N0vAF9750rn2Tq1BzUa+L98VZbKH/QRAOaOBqE20NaxJ
HZu8OLlH9hzKcG2s/WZgGGbgT2CtivL35fcfEhyKV1OchSuMBhHM3gCH3Xd1I8N2VLNEZD45hlj6
LfcASvh7Zko7aaJVnKEZgT4C6fcfjCaVzdPmjvcWUwdRiaudyVyha7mqmic2q4a7sxkbvfUtBXBi
q0hM6V0yNk6CCIvbaPv0z4v4oOzSRDHOmbdr24RIYtjfkeDEV+/XGmDA2O8DSNgAk7uyCTB9wDF5
QmOg/XbUK/zM3yXzMwDiY+IXK6gMpBDc7w5tt2ZD9tCoaksHwsxBSdc6M09eZR050905EyMt5mJp
HmTOy3ePZZFBs0Kz1Aq8Ozvrg3ooTJYUi/VV7MAJEN0KDJ0iE9uA0JCuGRvz++jHovdSZyB4Z+oA
aBmTEJCadNdcGyyS76m6bSAFNIZt9AirHWqXX+d57PVqcj6ycfSo5pjARynrW7JLJUtG8qlJY6SS
TNZeHw+aNA4KmNfbazNsg65awiT7tF6USntp2Ud40sA2RuveuvRm1EOTrZGrO8eRc5FrWoVIctFY
xRQTn9iwAVtrMvQKDhmsBBqUSHjuS0oxfy8kmf/0xUcucSTOepWDvKRtv8FqN+p2VStUZO3KTQ3Z
zjRSdXS9aO4jiVx7Pc03rBeKGS42jzox5Az2zO5d2WsZ7ArS/AfuuEFcDEbKTcSe8mrY4m79C7pt
NlgnLHvJxyMw1ObAV8QSjKy9faZfNQrb+NSgL6TWBC6u5lyjEacEYxxDWlmKCuzIzskEIeUXGPpB
qARqHgHeXFkZYyNZ3m2wxKIqw/EdpSQ3EX63VmPXMHt0FRAQThcokFhpSte6pFcvQ5QRTLiVlgGd
JpMHbVKJH6OIgx0HddRWl4ZG3Z+a195UIDMSfn0GPD5wEjdr4NR3GlPcC0rYYBhv4mWKHlb4HTXg
x0u//f8zTwa3TiJzBUPPZxhwmhJ2Am3qUA0NDwJGwbuX2cy7H04CdxJdw6ym6/z2GGy77POhsNlZ
//iozt5rKyIguO9LqzpLQZtL7r3fVVtqJq0m1glWbcRnpFtoCnsQdeQFXaKAVa0L/nBRTNFdM2OR
5lcmO5lVQwD81NI9xhQb9xRBIdV5aBcPBx0g261/euc9pzQuPTE4xvsan6xe1xHwtx0Op+BWefV0
O3btS8gJX23KCRmID2QQ0DZj1dJB2dOEgppYQkKONO4XXDZ/J0pW7prkGo2zMJg1FDMjc0oVPY9s
d9iYSjDRqkWpMJARZQVW5MC6wfzTRq56Y2bGtHd6PkkiikP8Me5AeyFu8uqBgFJn0tewO4b+xndf
kr5Rj4yCxUIgJDUc0IbdJiwdaRBXknijRHkPKASA65WWv+RnHjcuy2ZCLEqLVaavBNk4A2kgWDSP
Cs7NSsGzK7sXH1ggsrsRxoFzkI9kdhvVxf81uLshh+Z35I3EjgiWAA/wKWcIpA7fUjKFDcL7ieSC
/wbRZLR1Kq7Y6VHInJ1Ry/b9l5jM44wMJrOdav/o/qw0JCUAiDGFdsllRZnle/KFPtaryiS8aTbY
pkGkoSf3K8UoTI2cKFpIyfcjCYDu9R5z4xtW++zDCx0WPX01DuPoLqjoUopI+1R+6ZwYL+zrYqL2
kOCq7yAeWcsmVVMclmAkuqXIUhhj03KNO2eo5m2mWWASPntby4o+rWnyQ4veVZdYRWntLkIAyG6K
XXzjWz0Y8XnLBMHoHY9ZsJJHuGukNR1w1VIJmCI1GAFMEtKi7/vBt79HROQsFk/C9qQNJHFN8RpG
k8XNwyFFGjsQp9+4jtsb3U/QTPUCyhAZOtOnmu3g3t7nIzux0w17w+5rO+TQLYn9BZGlKfKReM+q
EuuH2obqU8ceajLL9en5paSwoCm9+JjvvWAsr/8ocs2IWHRDrcgrWqhdTHpTDhIEOujH9WBYppbW
6LdyJLRVkFgAhnHD5pWSAoErCzLIEbl7iSfnd6sr6zQvbRnyyXgrROSySj9h7Np8Mk2O3Ymo9ktw
ZNpHHGezQE6/Z5EyX8n7Zcf56V6+ecLSOhfmXwkSkO04v3kPRYvY8c8zzspH7WtuwOX4eHIgSO6B
is9Uj8+UN2M9MTqE8Qx1oynsRGSB2zh0Q09VMkLXkjzUE+ft/O+XLeqyiJ7i+7Et0E/WR+pl8ABH
7k3hVH5gf+jG/qgxtBVMJTlGymXjjwdKbYj+DvL9Bxa9c4MUoK8NSIH6YtzytDNqtCvGOAacLvhW
dkS7EZZpC4Ejgg16J1uUOXX/kG2KklSbIaDJxqnifFLUAOV4xryooF1b2cSf11SolXGiSAaSeXWZ
fce3cnBEd0KSi8rWIpES0K2IxIFlxRbUwK8B03RBObEQjbYdtzxFzLVgFaSmQHyjeSz471+Sc5S7
dG4pJ7RFenyaj9F86Vg1h6QyW64WHQUAWeJ3MRJb4v7jZPUqbDRz0FQdVwzHWo9KXwfkdSobrbYq
ZnGXMwDSvpJuEJ3y8GPbhTRljYxfw+U6YziujrMlJKFONH99A3GDxyCl/MUT45iAK6gxuo5/iQqN
zcYAATANvqVMmurlLTUoLjeWzMv1TDrJ9qlAmbY6TI9dEhoIfyqYxTXITYmDztveBPfwMxSFQhBO
NsjV8N1MpOvTFokg33/Fs6f8Aev/E+MttRMbPFCaRdT/Y8Y5laa6/gB38lc3rhr6m8LTcokfHrBZ
jd62wQbYrTCxSagElKGyZVe3Lk7+9MimV4LsFV1gjcXUt00n93YUTLXfQleOY9mlIPXwzt+hIFwv
u4ARrE/vbXtufB2RFWSyYF+lfnGfHCqae+4ZHrnqnLnlqWLpLxkWF/ePanbFW1nFC7qNTUuSq3tw
oD6YKQ2eyiaKHo0r7QdKBTePJoWUAoH14kqHIgbiRADJL6W8lW5BZGN6yBWUErzCRh4xH55O4uFm
yVY/uuiw82vGv4NBXhfuFhEgNd/0kd4KxJhhCFVdUFPBmbyKPpaguHY1wUAGcc7vtidJgvOEA1Gp
sXizR6cDMpzy82xfbmdbp49Qf+z/ilKvsf2RA0M3dly6WW0EF3W1Cgap1/WCcsA1E2jjCJc/O5SQ
vZxIZylMP1+SV/hTHWBednZaCpw7fdX0jaZhnHRR46E0wIoolMAh7Qyy3EF3Oz5T9hiHbOueEXvB
WVXbUjrbpExE3fYq5nejrtrHoYg9MAJ2Ql0UrppgHbyINxqm+xR1tyZOnJu+L0yxw4z7lA/jyW2A
pMHudPmPKiXcl0m49CrMu8QHwPwam8h4BNPxDx4oTfbz5TUDVzxRlzvpwuRG8ugyDJjgfCQDi5uW
kRjBD2XMHB+ixBsGqC9zRm3kbrnRWOi9RwyZTSSeFVzpNMwKhT/eUcZYYjAo4MtYkiUpMZEYagOZ
CRlpIQDjKOfup4J8QHAU/d4OOPqHTqCAOgPSGuOkl0z8p0mC9c0Xa2pUYqtA5sQHNVUtt4T+Wa4k
/MXu+a8gx/oOv+A+9ywDE/oZpriHmeoCy1puT/HKKYxnlUAl96GiyNkW8fR2DgWfUsT+hqUaY4jk
1Zi9paimFcvtsr3eaCUVHakXeIOTatouyjBxydeHTBFWx9hUiOAV42XqbG5+6EFSIXSMTuN0jKwm
XL64mzNrbDM15/6tBURd5JZshSYsMbm6gTNVUl+1bdrFfqzZbwYqoNa8BOYbnp4MYvxQd6Wu3Fco
2+9C20Yb+HQedfiFy/CQctoJxTg77Rhme9kk+JFXC0XcAgIdv8VOBuBFBdzPRp8nyG5d/dEuKN1I
bFi6oCSTYa6M2yBfsqmzvP2QBAtHWKjNkFzLuE/PqRlBPMHvpZ5Rk2rPrL5gebRS1etzBrRtqv1o
CMU4CKDvKGrv15U3yMxp4koUja2GCDrVaBipCNTJyWkaAIZ9J626Y2A7XZXVkdueWyehPjCraokg
XWiiUQaMfR/Qrb8T3nNfXfoMFkeYIOBQZ9v5dCbN5yBFj5Pxrg61VYHyUd0aj1l/+x6PjhCuaqIU
Kqd7oR54JuoIoIi4QD+xbSJTGpc+ynHlricIHxACAa1RIJQqNA8A3UPcmASoGl/SX/m+FTlF/r+H
21yqdAIAK9Sx/71TFWiWfpIHw6V9wqEJdo9g6+L50sC7mFcD4+CQmZYPRUP/zp2pnVQ3vqoS6JYW
1mceFMoso+i7BqvH/4gc/W3LGYgXI2eM7DrZwFM5VghOiA0Imm+lAG41vm17fZpyApG9v9yIaWCD
A7ikpI6Dgxu5a02PHsFtu8l1jldNGzfF4q8RBdtZjJ72OJCt7LK1lDxnz5pRB4cPOGsaZ9rgyN/8
chq5FqWAz3aZFhbGJCdU8k8CcHaNqHQro7I2K/PnAMDXKZaOSQRPGo4sRnjGlvnn5sXCkz5pn9Uh
HrXGSWRA/hlzbtegnTa7trrwvizjCd0AVnD5YJbbTm4HVOZO3068y7qSHwiFqhwAphiTpAEEHjwA
zEakNxfSUFnmkCApwijKwwfV3j9az4cSeB/NoLDRUiPVSgo7yGjvpIDbOIjGIggrcXLfImvhSPB+
Ik18Fa41SN+ht/d1My0rkEo79b2pC76M68hNRuNmw5X0rmHyHzy1Vr6epRwAdqoyChPSYKarPIDn
hXJBx5qCFjNjg5S7hb+I3QVotaslNh8+1JY8QAdwe+0mKHM1cxgnW74mO9VzhSic0z6L2/CwnylV
4wnl9ho5eXswDnnQ1oz0OLsdlqveCmVmlSp8GGGtFmzodp82b2Pb1vBptzMgfLsyDAsYcx1EaHrn
oiXmPmxYWLcj5coqnYfLUXB+yPXvWkJW/67erizXo0n98AyWAjHKMn9nfSjKxfM7TmgO0KpvzTKI
Uo1Bm5a6uySqjhWkQJlmkjYdGFEuyUWf8ViYUNFtk+a2lIUE1nzov2O8E9UANNoQqh8ct8V1Ec0r
u72byayzXBhLgogBaUD6tk01TdAm5nmzS2NLwW/CIagIZAQkc1WOV338ebQZiet7nqyCpjpI82QA
+y027HUzjRYvrE8Eda5SBp9TFjxXonXSo1zQwxcyQZk5S715qHZdpaEMpDGviTJKvNwfQVG0FseW
eWWcPCTim0k2APBn5VF8gyHwyIyi+n0A2+Ldngo7kzlFr0BcmbcHIOSiu8ynv8X8XpJEeOOP9Trv
TKDUNkNyqAgm0o2/01CHFzR7H3quFFdoQL+iREefVwn6QmNO3mrVSvDQNwqqufTg/HT3Ak7OQm1y
3/OuMYtetKDhr08IEAi0QK5Gx/QshqklQUQr3/KIHKWt7kNFCbcTm3pRLwqkoQ0rb9ohKLHxrMUv
Jz4edMlrF30GR1zjtb5GZulq08GtkoRJIVUsBP0UH9XbYjKfzSCroZHqo19s7xv3eJLeA24c5JqU
Nn1SiGfnxn6OWNcoxSqLy2esnV8cMSh+e19hq0ORQAQvSnytZgGI7k9LJl+JQC9srxycrjV/cAg6
zi1egn6mf/xIwnvZKJ78QsZoPEro5/M3f3dTu5fBsTXXnOzOGU+TOa8Jwsjd5JlbiD+wuvi8YcV0
z6YHT1mOAEmc4wfcVE28SSGW1H0o9JstRFmaowNkUYMgwe1DXGkmo6p8D94B78yjL8dKleauOLcw
PWEV3mI6eWW+WfE6C2O3Pz3saovvvyMP6ZMLVmmcl+3p56y4P6P+W4dUatxZS2HAO7XBXjxMDOWW
08FfEedSK2UaORi2+Cb++XmfJRUte5R41WL0ksXBwzXRkLuNsbirKZGLv1fn4oDiS2XZIlnDORb5
0mtrJpFKKahJYsoUNJmpaOiCrr8kOQ3fXBg91eo4/gZyVSQMUYOr+gExqsiQm4bV9QKJACs9IDv7
XyopAz64Hj440kI7/SSLCEZ7GnanPwwmz8UsGloadSZl4fZK2hpyH42k55yWK16AEZNjb+Ty1DzL
NmJlvfTA9Ikxs4z51HzMHogdZ9Teyi+D7zm+7mN6+c23u0sS9/dmR4Y0nHGJsdLrYCZpy0Mynq83
vgcZIJMipyl/EqoFkm7DKhaH63UldxUkjBXkC+XftkbfgJQV9bOP4MfSFFCzC92NIWoe68K4CR8T
o+vVpP5qxn+HxeqNHhuLaoj8bJQbh6Z98N5LfOVYsXEedqCzNn3iI0FDMu6ux1to+kY/2fCOwG6L
2w78Va8Vl4xgNlIxOKk3O26hVzLeoxezg2E1Mge5wBG4t2Kg3DChJ3OfJiDdF8fb2RtN2ciTf4hH
p42sO+db6FI0PpVDTJ/8goZWXIF5e7J8G21YNZ18B8BYwZCzgFjmrxtB5Dqr5gDUB6ZjE756LuaT
DQFhR77v+AILgYTz2+EFaLp8HI3MWgR3wqznI2x1+uFxMo/puf5+KJ/eHpr47K6ilEufkJxwNSOw
i5hApORi+28zx8Vn6jUUIevBDzujowHRAF6hfBaFLYubWwcBUspd2JLQpiEozFdSoDHFyNcMjcsl
CT8/2mE8A84fIcdSOr1+EYcE9H+yoRSdT42MXdVkY01v+JWMj2G/uJCCDbf0KnmrJ2F3tyrEkB7X
E1i3TNRCPhaXHbdrGWHlDiRW9AKVJuVZ9ryS5u8FMD6AeUe6W49PlooQUyQZCXyxbj9/+4rhkJVs
sJ3nHzgtKMMV1ewD38qizwY08hZXO9xU3/jlCjfnGKgJEg9SntrF1OJr1wYGre1KayVJ7MdWQbQq
ggzfINEnIYY1rcKgxCeopbVWQyPV1I8MlmMCsBw06KsVCyAX5bGTrvzd9sYXGYiW+RppdAv78bFE
hnw/zWjFGecOTKc6ZYh7PLGYnpism0niDcsSC/aPx0QiL9vwXIbAbLyDALSbiEm4l28j5dP/ucke
8QnvFrM4VxWC6cha8yqVfFqyvdSjiXcoLD5k/swDwzF6yNWw2CxJw2mPCn6P9z7rt0URq/AoV93b
N5B7oedah4ktJ3sgNwGjmghHLscMcgCxUseQJBwzGu8InqJ6u0PbFAsRsnoOWsPTfG/INNVsQB/p
1GGNlaMh8n14ZImq7GBtSVGSDSce/efVeW147SHdDI2fULTkOepU0O2+Go3wCIsHwIrFSGv6Q+Wt
O3W737HUQkuQvNNDA7uMjyO8iY9CQNYRUx6zVUH6gkRusOUFrrUNR3iNQcci9+ZM8jvNqy19miQW
JqlGw8OIYXEDabiyoz7c6a+stoV37ex8SaUFXbRgbH6gxYDmd39GeMUipLTR8v/dSmRPA33DrX1W
Dp0V3bSFu51ws9RAZDnZ/I+ymtDCFgRLRUzuLt9xe3WZ+6i0IZsZVO9UMncSqC8OOK/tRIsItERQ
GBhTnwb1WS/ZX8+iLL3w5BGBzDg5n1/Q4QT9jl7OJW6b7hs1A3pYsMnWXMTA8TobsHLUZgA/bGtS
AGBwvwAbbWjlorNUwlbpXAoie1CxO6Lp5eYPxD8u84zvgKaybD4nYB4YlBISyNzfN3Rkbz16B6ND
jeuA5koU8oYoX0uxhYcRcV1RcKurfUbxn+cPqTR+slJA4j7L1Ur/b8jvfS+urBH/PFWkWCqrDZzL
5UUCKFAiBK3nJf0BvFtCPLzsSnFIXD6OEFkcmhl8uc9g6KWgGsOjD40fJT6TTWkgE6ZB4uRowSOZ
/VBhJ2i8fX66tgVPT5SuiG4070IYqAXMEJijaHYtJMdKoypCOB+blBm917O6rsnSi5G8RvTdPPWO
JovvviFOXDRiExSW6x1+tEnXJICspYeZWTgXvq4/rXkHzYP0tnyvscX43vIBsQpQNRA+XWQ6eh3l
6d+72XC4fEDuKWCr8azLFqooGAmPZQn8BwEvhCWXJm3vFHNrFBOCLa2ZtaQT3BaKj6DymnGRrQnv
QLqs+47iLnBEY9P4Tb2ecQuoacQckd8bhHZmfvPHsYBQ/+GF4qLHxGKww7VDi0s58CdcBTHnOgWT
X6rw/+gyu5BJLcsK0FhKfM9S54muUcHyqrmWKp84yTxkrbqIB04zcGd3in30SYGRNH/JlCMrFH8B
Vi3HSLvimobMgYK20v+zfpDfKHALNRN2mHjS22oKrcdHajZr/G7c296SPzW3p7sWm9YM/QcOZaoo
Z5K57RL90LNXsZC7xZ9o3fk5bm35XNJ7+8bIOgHxkJuSfJudSPySSq6zQlEt9x/sdkXTCu4Idx7I
ohmoCOBfp/vsAPaYvph2UdIIa/XOhi8EB3pTAN6TN6EKgl3+aBurgfRciuPqtpOWwvFA7SemxqFJ
s9EniAqVWC10oko0biafevCPralaIqLAZ2tDWeBEcGygGvlaPjbvGAoH10F50YivdxACK/3iXYtT
9R9CYCKHh4HRmSKSf/5J7fNB2YVpvW+PgfbtLLBTVQbIUm31PptULcVbmpoeOqKjA4ThEDyi9Cyp
3uUaEv3/DfivtWJzBDFqnm2Upp2+2ku461uiBY+soaWQ7Ya4HUq9DOMQOalHwvSJUoFtgMt4UgUS
5UqX7KtrjAyobslvA4WyGgysE0MANzltb9b9kOvH4/BtXviT4Q5x+ku8C9UmSIcnfQzjMxHX7eMi
ESBbXP/uRVxMUIZZRRNcjwKzEPuWjA0A9PBvwCim79q6sJCoKXOaxDFtc+9SYI21a9Uzz2+u2Wft
F9V4Cw5tkCKOf3VkWjwOqB76+vfJXJ+ydBNXeve2lrqO5FObD1Qrhr4wTUwWUd0jyHsM1x5q9vhV
03e6y7pdQNfAztbqwIrUXtb1JEOEqWg7p5d0tv8pg6B/dfG9hr2PgWG3uxUrBrLeB1e25kJaJ3jZ
D0P2uS4FWxH5Ec7JvyiRg3Om3CYqt4L4MqRrjxGu3U2JRFK78pUlO4uvz3pbWi4JRHqIMVIVFeiN
X3aSwBSnNiZn3nVR5x2bUIpSs/sXsTX++rZ0lrd+kpi16r+FSlgy5Rkaf7/VAVPuTa+PxQftiYVB
r7p/rWcMWJx+On6yZ56vr9A2WSOk4BezGK7UTGHDfPg/OvE4s/SGZg4CBW/tK3qnCNrsDYnK92qy
KvFSa5rCYqicw5+okA8tgJuUDI7NTZpf4Sy3PCC8/zbGBxwlld/kmoIOsCPRrk7lUXB3V8D3xDF3
0AUZE7Tre1Dv6+EgTwLWztPRrBU1oCo2jXU3fthqCQv+pHFDOlVMxr0xNQZmlaD1BpFz6sRTu9WI
Fk4ZuMVkA/j1iGXQLRcJCLN4q/elRE89jJ+2RcxKMuXiPmSoIWMzkSEOF2SmITRgaGAJamZd3iDn
lrMxocL9kFDLxotVvR/4khbqfZ7KXbIZ/CeZxCw+YR2iIds28TNrZREBMRwti0/zEhGxYZUPckKK
XbS9ih4A2SBKSClCL7yI0W2JhsdrfbrBHahoUiQ5e75PTQmU3vpLqYRSeRE8NFSl06+CbXDbZVo/
rMLC92dH4K84RHeZkExJNGCyguypbGljM1uKtR7qfR25Y4e7nq4ElpBEz73oyNGgzOXHxF5ctwOe
xWeuvO0td3hBr3zVk1ixnedRiStC5RWJwqJRgG3GiL7/kE4dJ+MtLVZ8jBEzQ7KaeN8oanAoTIiH
frbBjry8RxlHlu7QeGN5qh1MVKSR/OB2fiJEmnYO5ecBn8WwecxVsEzC0LqqWelW2Im7PUPp3IdU
jzQWGBGUGg9g731Ux4+ZqVH/4OC3sPKfzOIrVqZo08rBk+JaX+QQ2yhKHZZk4asXWq7EuQxI5TQI
w6JqOhvil/eqnlDA1XTLkdN0VcMi6wkjnue4UlYAS6P/T5zk6XHigQQd/uZir2NmIogDq2dzz+xh
tor4UeBAC8F/F+sh0L1e422Edc7NQyxC9rlvj6IK6wfck49M7JEYeOz6O7bclPJCYsLRMrA/XHwW
KYoBIxl5jfER+eZmjJnxr30LzO2pEA7PAcG+337lLFbJmg4Ogp+5nwWDhmdq/eWoEuZFVge4SiUc
/NrJ1+bQs3s5cWd0VawAxQgVUcuvF+BqnHl55h1lOHqjOceqEWJKpz2dfLf1OUBEt6ws22h6xzJt
UlfpbfCFO061kcYLSSnDrl/OhI6pbvgVMzE6kFMVYSctSVwonM/XqNp2Y5n6lrjis4jVXOkakz7e
7Nao1xsrEh66nlCWfaaH6Hz4uuH2tN/U9i8A9I/X/85Yu3pwKWyApdQGhbME2F+Bd55H/I/pIDwj
CqFzovO58ZUeFbtkEzWKavEJ6ZO/QJjynt2m6ThrHLFNUOls3ZdD2v0SzOycTXwMHwqPRk7Ss1qK
8G6bG1djfQIj8btN6IknGmYIM7Zi1uE0dr5ltty12eUOuSgB9vVzq+sym/pTyFepD0KxaPU7+puS
LGaKkZ3EEKTKlETwQXXiOEGZQx9oJvcPdjmP6hqXGnmxw6u4Vfki5II+g/nTKtA/6xUST2hCKJJc
1dwZ7ZtweWnjNqVLRsXsubTVWn6Fzo+K36WDLakIedGwBRLeP7B4DF5VHszJcLKRFqkzbw12mu/g
cl0G91GdkbPw4/FBxh/6VS3HYXgEJp5RHuNAWqXXitZUAOkhRYyjpibKcHnvVs0icUF8jnoQpo5j
WLjsWQznllnSKKPNYxAUP1mlYCOifiLBFqpN3BA6jK0/UeyJ/otzI1EbJ5BDwP/4WRuE/zYlvDmJ
EZ4TAPrRgVWHe+6gR5mfxg6I3uU8t0Hpszzi022INcA3KP+FTecLP2q8cHHQMAucCWcsMyCxycLe
CaBNQgFGR11hbtPYxG7tZqwmLsTQtnDypVjLV6S6Q4Z8T7eAzSOCTpIKiVrngiQWjD/YwtfqVf14
kQ8jw9/1T7eYUxmWn8C7t2lumstVJKmNDgSO62WnVbJQkmV2wktcU4kvNHTQ18C8b7WtUAtcmgl4
FwfH0Sh6/A1Z0m9A6bZGWI0/A9bZ49MF1gc5nUqxMJ4T27n/pPYFA6sdLWIq87S3jnjGP/wclPZT
jB7D41MUz7KfczOWPEs/XwXUSXGL6WzsR1n2NA/xa595q8QfA28bELihBwPPqIyNrp1yhQuLzCUe
fFdMc0fZYwXkZyfAOq1QwCT2+6SlSwx4KBUNuKBrPJuXMcgsMDTip66vdWedtGo4P4gTQ2kFpFm9
IhNgVxocC1OIi7SSzQpa5YTd1OF2yYIRRBoC+AsSNsX50nwtpt6QsdxLE9SP8z5uNUVrNdHMLEEa
YmIJnwffDYS5pv9xgPEOpiYZ3qQSb+V7pJnM4Vl6aXMcRNrK49pS6s5tV1opVMJpeHom9W8L3DwZ
B22ty+Oyk6ZQbrDOMtgYoEOrW58FqjBFhJ4KnGyknEGX+mUC43vahQoDK1jhAzWVNHkjiqRO2fwF
CMFBHUeBGGgfEVZ05Q1vGzZBG3xgbM2gunMHKaeNMphlGVKGDhyBpl8nHbgqslIyuhNqlfA5tOsG
jZXckcChfUJwn25U+OGypFI85z+d2nLXwRctFCk8tysUed0BiuXy46BwMwB/GbLy/p3g0tIlDJ1Q
ccUnMH2kHK4HV4iJeMCYIIeKDWQ9rtEPGQg6iBGEIp9aVrqciX01krPQJLChUpJwEH1+ZnVgQ1Fe
Y92YMVtdJtAEgrnallOYxIo2IMw1jse7Ym229DrEMhwgIRZ8HCmvBaqTQGNfqOs00hm9HUUlASwQ
bhHTXxeZJC20KRHvPHZ6oDjQ6rJSYJSD52e6q9qCfwDW5QYxYm4PHimPx31wQKwaf1N0MHq4cJEG
vpqSKaxnH2rcfgsBVk7qaIa/x2co0WC61St4ydefAI/wvWRgBMkrb0F2p30IUYDkPZO4BZEF7oIN
hdKHfPeNNCcYwZDOUhxeJpi/VAAj0Ry5O0KrPcMorwtzeJawC34MEDo6FWovMKKdM65P2Hvq03Q9
q/z77wnXFBdRywJTX1B34CLgGfoSp1iG66+EBpKQ6MKw1yEWx9DnL1axfxC1W8+nEgB1/4HH1CLg
Q5LYDNr1uMa5ceFqCgvxK1aUMXqcnuJsyTfZoXVk0QmgviTwqVIJvW3rMi/q+/3tKwKOf62Faltw
6FUTmp+zzRdZb73HnaAHDhzY5gmS7xnC/ds/qAIGD16+sDfYpw89i7Vdun7jKTlTQo8xfDF/iqV9
vDceuF27LvUDvyZPusrc4gIvaiAUfjOOVZFUqe4gOAJ8Uev2Qzh2eYtnAb/T3jTekHaIpdfxZP7c
YG2hzgBTISjoBS5IzOzFm1rnUZ+RUiSGWcBWSrWiy8SYQwQHb8JDQG3zSGaHJ00BCaMrqXrsXohP
lz1LQOgvzXfUaaKjtwozxachqZAz2MyEw4Kit3j1I2dAGYJGYHQTW3h7JEletmtUZHGk+32G3JKK
MQb23jb3UhnPrb4wlup3cNPlZTYq3+ptnzAsIXfhLpPPS/V58s/LpwOq7OXBgkZ9m5jj4Jqhuc51
0iIcWQq9smJklHh/fg5srt03qFl+WAVSMmpU2g/3KEHlmXGXTiREyrCyc9NgKgq+1KB+kXciH+cZ
ZdQu5j7uHVx07AeQQJACOR3w+7kTSjV+iUKSfP6f+Gz2qcaYZAW7s/yAn2LQEEUxMYdky133tCg7
YHuGfu5dwpWlYBavC/A/Ez1AvD5HycEsZO/kVj+F7VBRhMHHhb5eDaky4ZXB0GnB/VaIojyR2FOm
B91kNcjCluVTTkMDtEnwObQpAfkGv84lkZZvVZOV+qJJrYmfCDwCM/htPsgILQ9ohNlavwc7C/yA
w9frWEBMcDMDzYfSyjDmxq6jMrlwHyt9L2TMQh6pGteoToYP97ACdgQi386kjAN5Fl7whHiOAKcA
fEQYbnzVViQ93gaRahZ12HghBps7T2qbNROE+tV0aNiV+UDjq2RPMBi1BWkVHOtGClRvRD4c0iKd
kwW/hAFbEsuqmNDRegdvxILUWnqaDuZPz1cYg/SJpJBECa6izKP230QWyqfP0UowbdxSpISnpfhx
2J6I9BZAasazhCTsr+PnQ//EsGQ92PFKQXCuYSG9+rylhYYP/G45FuLsRnwMwbdi1UWGtQQwEDaH
zgtAWaICxg8DCYtzUOUYLpQlr1WrlmWjL6L6RsyJQ2K9QDRa9zg5xjY+PphYqSPZDtijnhxukzgx
vYI+JPGGzAwalzE+/ctRiNfJRmi4ZpzAS4ol9z+msBoaMcJJoAM6nwxk+Nbfj3X/wCwQ7dhYLtTv
XQJJb9t9Vc4ghfiXNirMr90Sp/RiHdZr+3Vmun605ATttLhYfe1R1QhGCieFLdZaBKsGLxh+6aGf
MQ6prXuh5r7HV45vwRR0xP5ri8+/pDjla6wHY05xIdWWwMA2UcbHWXG7HVb3gDksHop6p9jqUvld
Fh7f1+WJFZbP6vpfYbhv9wHjHVLt6uSyym4280NTGhP9BOHjD3LttdrJtNv8JXnk+4TbB976JKK0
I+a0fvfzV4QMuakeYH57NwSh4fEReEaeqYWKalQPLWt2fzVn1vA07Qi02hTuyzdShvMFWHZk3+sW
rsNPLxdSxGbf/Yk9yw2rvtrqoqJbr7Ij1YN9rxcSOIpo4hMy2j6v7qRedGGylJMtpeato7QqYjLM
lQNCSRuKq6G1/tJgf73EhKnOzlaso6Ljf5w+jorBUlSUbQSGprrPdFGqcxwTzgEanLztfYsDk+tZ
8c2y/rpxNtXOJsmtOXgWYqWUdlwj1YliUVjpMlgehWIQtox6U6zjZXRWviQ3nMtX7uKE7ba3VWdP
WEw69ksN/jBmQIV52Kx+f0ga1bL6tkrWrCONPuwORuzBb6n8HSwivnRV0b3dEzARJNamLn/Kz7U2
WmyifQYWD5L2jUOBLrOGehxV9gCdeGyF/csh+fp4AmQK8bVAVYwR7au/AEU+Eu1H8kWDiqI3TE1j
5J+qb5ewSN/wTmqYcbg45Uzvq1N3Ty7QaxBT/G/vC1evkIjLJKNeKhBRDeJvoguCWYwOpyiWtY9J
D4JwwxxAf6/Id3tQ9t12uCSaf/+n2l6Hd0RNgFaCkjaTgC09A3tXMgKf6wmSrS44C43RZFEvLIZu
fqtpEoInbqinNaL5SNECFZhDMiW8tMbc3aL3hcMhD1m/Wa/lHvseHjl/LnfDru9/MprytCQrI9Y8
cTtKQO86+uoxsGnxAgqwqo4m65a1e8psLFJDXXJ7OzM66tn/IbWnTn4MgvM7QT+Xfg/4muOP0CV3
InOhhq7wPmawzGeOGDaKzdQa8JPLyJXKiBQzVLI80hVJ+U6C9xLMVEpRZ1IoNCyT5QZKyx3V8TFH
zofxM1D5tKxfJwvn6+luIs24MFXlB6HxgsjzAmqz1YDTUr7rddcB35uSQ9uRm13i/BPhHcRyWcXD
XVBGhbqp1G9YWEgr4+6CoabSy3cD7KraQEDuKohwn5pUsxI6nJPG0prY0nIT3BEPw6EXdZO9PzTM
uyvJLasTXqe7NaMeRwBPjM00r/8HKsAfFgf5Pmjqqs57Gr8FcusKzn2LvobOUsyEcDb/KVvzddWO
TdqcrBgCpgK5HwlhHFMzpdMgWXRLBEXfNRsNWFPsr7VF6ek3FfBxIRF4VIdduBIuXYgKLW+UFNmb
ED4ccuTR26+7HSDls4WhIsSMOOBSQlerzPEQ7EDa0Fp8Zfhsa825n+CGPfu/T9Rwat89EXm1WNQx
D3AFZZDi9OADUZEYaU1jvwQuzuiS4uRVWunjzNvEzFzhSeePz+CUdHPa2XPmDDRvAf+p85WnswBP
xbgNltfGjWkqWPUO8z2V1wgXtE2gnSTi45xUVYllYdoAHnZh1IJFAafolMaK9iguN+Vq7pDSJj11
Su9eA8G/W9JuH7ckH3bSogaASHZTR8p0xGvGsmv9f7M3a0dgoax890Vijyso5X3Uw381QW7wIVre
zBSm5qjhVIzOPOuSjZzmjUzzzEw03Uankkk+vQrPlegdEXGmsuLyEW+MgakQjv/X+ktZ5cXyDk4D
JjYwcyyFKRQGj2zZfFzBOi/oljdPyRlOsHqK6vuvlFYLEc4sO+9j7nvwC/8XZeg4GajIxsiV1BvY
ChtFofapMbzQFWnLyM3YLEIGFkfyFNQd46CbiMGI/2zr7mMFvXyXvUf3SQ0ZouhzIsisMhQaEPoI
OZ8vjJnkKPy09Lc3rJe2AXgSo+TjIjzMKbFUaju2NEVjP20YVegtY+23YhETfpN2zWJkH6MsyIH0
G8NtGfslGUtLr3inKWf4mm3a6fRvqmSpA4n3JBDmM6Hdzy0wEQyW9q+0C3PcSweeUS6tXJVQxXBD
WlAEsZeNC+mqo6sfI7+lzNP1xAGGmDlSrvo9h9LFfwj1Z+7FlcMbCQYFbIwzAAvRjt1vwaSh1P0q
uOqYPLFXcuDNCO0I450s2U6z5kan33v6j2yc2Z9+OSQX+GDoQJnN3fpQ/BTh2E/tL6NiQZ2jyR0k
S9vtaYrMW1sDKKNbmxE9ORLa84LVJwLVm6r4MEivpiicdwf/f6g54JGodqmxQJ0AfFegBSu9hwKu
P5fMaTBag3pFdGtrj7PMTn4wCxo0uEbGACaqfEvFsBwItBUrnZNgpP6eYG24iOvOgjSSEmG28om3
j51odHNuG52aVSQaNvVmP9IXFXQyghSWhM8ewdqvixhKGq9NyYtdWXxOC1x2FwaMb3LFQLVS9Q7+
T/VPRnBDoazdh+0A1h3b9SWNDw14FZiX0ixxM7IHytJ/+ZDTB8aSkD8GmxaIkXcX6IQLEQbZy3Pd
fI5jLLHZj9HbfW04xT+N0NrrtRlBNG2ZozFPsQAzbhkvgtRb1XtuazdhzZ7XxHQlm8BCDS8iH3Lq
9T0HgI8LIIlxZ9MowF0SWG2eDkmGPDe/vvoZDkxonZnyR2kjKXlk0A8g83fxv9YBP1N9sXmxky4/
J594bTXXsQSwkGd7oz5rk3bKat9fAUuz3nxcRX4RqnGQRMxVgaaJL0pnwqLL2vFx/Nt/F9lD0jwG
6Fw1BYguSOl3pYpOkVyJ+2sMqeicvgLVR+MB7u3XEo2E+LDF56geVhaN2GJU2ia8TEZ3nWo6NMfY
sRg6aEs+h2D2TAFivQVVnTeBFXZ1vmagaaExjkJBADoNCi7Seg6Lz/xkc+ijgBxGkhI0FYBoTNtt
yYrBeNAYUPdHXCcCoIyU6XuwIhLz9zyO3xGCHwUx02rV2EZOCQmOCbRRay26GoFBXACkSAd+UT++
QcDEhmZbnxORfhsEkNcwep+8ktkxa4u4OIMDeEQy7si0X77gKs2Mes/3nVf4nGyydEX3Hos6iiHc
jIkXLCxJTPdIKY8ZPjj1vQAN9E3sv86588RKdrH6aYuCT4CfbmiAAhokyQwE7iKg9bYehT+gxgxw
op+XmIFWBWfoKb3TLTijKP8T4i2ZOpHEkeXdgdrv+OhZq5gKHuPqBW6xn8fGtFkdAyMcs0DFLYEO
GBs/3aVTjzyePx9VnJy9GB/iyEWrGensC0HqP1GvkPDerxHDDA6WE8OjsIlu7S1qs5iKttUqF230
QBKaZqMKzm16hOTR+Bxtxu+uChpk11NgrexCNKEfWtvQcYLWEZGx8w4qxPIKJ9AzI4cwybirJz9e
pMMbO/P0gKNU28hIrZz7xTWkas3X6W+L9U4yD58tWbGPNTzJmW9s1MhGiLuXhSsHOlybl+ZnGY8s
TtC1jRudDlFR8S/FGDvS/cluVh18449FwgyF93Tnb0T8cVjWUMZStrfBWF3lSV3/Z+BQGlu0dr1h
3tocMX0leVeo071ZpK3Xem37wHwSOM7l8U8fileEA88FoAJqLaupfHqpKntoR2xalkUqEypaVn1a
rdilKVOKh2uPn+EJ+PRyaMJJGzu6MRDNE/ZuMImgIPKo/YUWg/L06gU5Unn/4tGlxdKBfKXgqAs3
wpKPuzF0zlJ1IjQF1T5UKSVq3w4vFwfTJ6/jq7w0JVLCqxCfUFR9BA9DMGKWcD4B0Ofkgy8GbKTr
KwXnHpI44JMy2314qZ1fvaZYM+Spka3GQde0PxnYryqJGytC4KI/1ZRrcXcEMATNQw7PveeMszEf
bTPtlLfjoB7BlQn5odRy5bBJk11j46qJM3BqjudR1/l8VLj+TpRvhtcQr0GOEf693ks/9loQnsLR
n2x35m1yGzc3fyuXscEVz3hC9Bic9Gw/ycCMpL9Z7CcVGFKbdmuxXUu6rOvgzphqd3sqi1vWHnm3
ybqeb8RfIiM/pTJUrHTKUlf2A3liPfDYdwulFagVDDyC1k/IAYBdi8IZ5yz6UDCqCePay4DLT9Ug
Qhhho5W3NSWgwBaPFgqK6FbcFBp2solHpRfe/RqyNogr7ABwGv3sZ/TdgHmxzCfibPHlyURsPAhi
amSvr/3pg2ju3UDtuCCiQz8YWnWWvdf809EGQ/ZzQVJfNeTy2mQFBwLNdAEAS+Ri9EWPdBPllyum
csXTJfPRLukgimwENoaux5ZZMMpZArruf7If25LUJp7T49/txWcuAfXHfIwOqhp3IyH+DW72ypK0
UqP2CDiQdetW2EZXOPQwQLjipO9Uf4/U6gPcEXeHrRe5Hp1vBz/AMsbU+QK5ft+ST7CwX4pA5y53
Sb2GailVhZjCI6au6fhZdP81QjIR6KE8ujs5knQL1Ix7znyRpgXPk80vSiDV8ug2mmN3dSVBIsFc
He4U1glVRJ5W/DkguRwCq++4YsTqUO0b/R0PGG0H2P/kcHQXZjRl1bLYMqRJicLwTtrZPce+aB9g
0hh7ZtNWfnXXZaCIkuwk5yDomHiNBCoOJD4ox2svEfVadQec8Qf4A6w4SsyCywLuWFf4JYfaeMJD
RHz0IizEwnm9pO6iTlE+RyH21qi9Naum32OAuHQZdspxwbctIIw4BMo1CyOO3WZIkbmyvdL+0oTC
CcTwwHPKGOlPFgOWSkTmpbpPIobLFR0UY6UK0b1QCmUSWtAM/l55SfJLOyM+YZNyvJ9mVJIWGASJ
HzTToKIghopS5ToxiIjrrLJ65h2WWQhB4tYwwNTotMtYmTHoFGz24hOU9uwiktM8yz1BFwm2m1AN
DFfVSCviFvd/3T5VBciZC1dfXFfIszb5qxf5HQooRPv3MJ9jhLsWfSrklndaagAGr8UCNMexwl1q
y2Y+sFznCvaBglphy+UEHTKeZNlveWG3kMRYDME2UJUln2lr7bAkACxS5Ccoz2yONlGn+Y2z4Rzz
9zMFreAXF0VS6r8c26zLouv8Hr7SKeF8tRBsTIQH5FUWkOmC5Fc/yp+Ti46UZ1yHsTNKcJJrArXy
Y8AKOJj0D7gB7NSVnkD2rXchYEq7IuxCwjwBWNWEUiLF1PXtM4SAt2t0s0v92gEypbQaXoH5hwgi
XrWhQ2LATRB81XyAeMxwk/MIlEDvpZeMr/9OxMvsEIHrCC/bKbH6nJCmvTWUYrJvkpSOgwLcLgH8
jWjD+hpHRJTkA7MSEB9Sj87M90BrThP1FB0m1QP2Tu2ghpxXmHPBCd357Gq9fopxjDKn+/7hUWBG
daUyyJhriBfeB1YEZQ8nIzQc+erJjd69DIGTAqUUwtjP99VP8FL0LEl9KlqgCicWZ4xwXK9ffuXr
WGtA/OtTNY0ej0JnwAc/3bjacdb8WU9OmtMNRYUP0xcr6tw/FcDT34kTc6KnfuPCj4f1vZf0Kv67
83FpIMpX6vy/2o83BJqc+GD3j682e7CoCOqiN+4yfnXZW6IFIzfmajSFpt/Y44DqJr3vB8vDmSRe
yR2yS+83sisxjiL+FO6XHSsQmSfIAldHYeYA6qJLvf1Uvm9SNGOvMOTcwxB86VfpPQf4UbqMXYOH
OO1ODsh2qc7IanZ2y/k/ipkG0vzP+EOrWpRl7oea4roqmzInUgax3skCYtwVuQh+0NISncyn4MWD
DSbFzCV8W0QEvk0H1DeM46udZHHodsFoO78FLIdKvptGA5YX3Y5+arMRgVPoIOnek4vSdskraW1a
VjmHZ0k9LKKymbUZ75Mr1P+uMJPX8cuw/S9aUzZH8ToNeW1S4kQkKD9iOlTMrheYqRGp1Oqshi/H
nbQhVUR2SuGB1gcbVF5BYKpsegRAzqGV/8Ee1EtwGSx27yNZ9bO/rW6P4njJXvr6hZ3A9k0QVcDo
fBsccZtqrqkKsfBs7ijgmq7ATpFbjgDJT5XjNffQC3sCi2jVazDKmE6ZmPOjTeYuBsGdcoiVyons
autFOeHqJ91W9TEMmj93+VDiWkNBXNTmJYhC5boUYtQNJOeir/kX/XhcE+cFY5uF9ll33V40Adsw
wdblY4l9s7WtyTrN8raU3TU8qdiZ2yVfOM125eOjSUor4gqzP+VSQhgoGnfnEhEoKxahiOBomiUf
cdoIDTlwzguG7JW9ytyAZiBaF5fIw6K0uThPmoWoWvWq8seoAoftuiw0J7/XV1+OIoBteRE360Fo
lroWyupVIh74TwcoSzCly4NWx1SkrHE2cjEUkiFOb09k8WT8bKY3HDMUCA759GSMR/GIPsJ00gbd
m2IchUmqEA7I0jIl9sv12kWz49dlrHPoSe4SA7HVVzEI/X8ZLXElXchY2vsyD90Eeenn2XGbkXMW
f+97XHqbx4p8wM+bBRxguvK9Gi3VDBxl59Y+lGKW0j9FZpu3kp42gDJLcMO5jb5zCA70FPItmcau
Ua2KLuu2RKOK10J4IE1W9UKZOX5IE2W55e2LhQepys8VF9q97X60y3VjAQqcLn+/aTArdSxtitwL
RLh8Hf8IX4yGe8eSm5JB4bLiIKuHTkB0t5GQ9N8C0hpfSsIspVuQGYmHMGxG2CGLVYMbozM909kz
0rmDM6f+PgGAhlqUAjIpR9zhvthlHxylozcHDxzcfPaiRlA+/xp/TtyDwHgY6fWFAagVApll0sai
0sh5aywXkgr9O4hMBmZ1xdFa5yxMH4JoMNv4+vXyz2QoHBiGGZsIGt8bweDrkRxoeyGhp13Lncbx
SxIfZuH2eakD5xJu+Ao9gcbUcA3LZKne6UQD1TkiLI4YSbNMLBKqIphEgVDbzc0cW/CFS00XtPEi
MY/2iyzXva2VRW67zJv5euRwKjmytrMoJ6LSINx0PaUIXvTLCo4jgXTs/a+uIPwjgj/vNpmWcUm+
bX02Tv54OBH+cT1iqru4cRksMqjYVoUY+IVEebGzTNG9VBoVgCii22Z6d8VR9I4eZynhZOw1Wte/
ZHZUahhcNrDAkkDZt7wG45JcdyKnOMLyFOBMVWuf8HHgla84E1Wqo8/lzQXDuWIVyudo8QIfU80q
ETJ8JhcBhm3ssA5ruShY2NRsyWTDok9NmrZB4oLOhuOmEaZX9/VkSF7yVbEsNKbtH6A8TlF4PhHp
2OgyCJNti+mlqN8et/5qruOtk+5y3cFF52gpmRQSXYkUP1koTY7rt+itFmtaFb0Ch/zIdei+BRQJ
G+2nqHvul0KarBX/MjCXS5EbIl3xm9qe7zHNkbeCEgVcLlJoPuEtJciLHGxrkPbpnvKZR0Uj74bG
dnuKQA63jg456T6oKnphPlxklTxlT2wBH6n22TkqOoZ+wjzfdkqvNigWMqL/fp+G50CK7GADR/s6
TdWhkRrbSbmFO6Jqw9zb/y3aXOI0GZTFaJ7Dswxl81JjabiKgR4DCEIWR5FwK1boEotZAVBOWnyn
FBIrjX4Qr+1bX8JNA3llJL8gLDPi0k2yb6ulHBT7x0zD3CyZkFK3u/NrNIP5l6ferQ3rMelu53na
TgsU9fpOJYga6oZqfzZSNFTSFPN+3R+wFvO0sDcsacbnh+iX8PrSw8TYqv4nqF96CF58OqR6F5tB
2ECnXK35u2ivLfxa2xBpKtWM7cW6LRUV8Zrote6c+s5BHvJTvrc7H5yURYcjaJnB+vCZ450gc5hi
otB0G76MhLQ9iCXkAzFVI02Gug0/ibO99CUQe/yxcLrhGohuRD9qXoFpztCZnaP+xUAWQHjYj3in
ImQ3SJ7hNYmLeOlkmXx4AgFQgi1jRurSrssg5IrsMHXVrkXf9RnwePgtmQucuhABADkH+zWENH7E
m8W6ZAeYWFt1jQy4cIKT0ghlczXDdEVrk4PV/MPM3uz3nA1mwsuoYg+LeCSBC8WTYLnppREwzEUt
IOBCx9rJ1RheqjSfmTWhDPfA7XqwX0LUl81kEtGBY8DQMZ7GOZnZd1gqZvrBFUoTU9FX2uSSx+ld
zXF51UTgsTy6JoZloLwdnI3wX+krMhlkBNDXl7mq4UhsbMngFOh1claIF2+YRXv8DOT5mYZ+CVAp
SLG/lBm9TaHjw7bVbJ4S1SP8SC6hqO2d5/YP/E1TddUTrkTPDicWnfSLMYs+0O4nqUeGIzJVTfa/
gvHXzTpKSadaTw4IX6xqz8OzUgUa04PUbrF7QDuY9be/p2FUdKJOWpspFyPgZrHfay0Yvmtwrd12
PoFHPF1gAf479jZsz+sAtV5LEVVoMC12uBi1qSXUSbQ2xYDmdOhhd+EZ8f1s3zgK7Krn6jA8+Wmu
aiQWqMUnm1ziYZYEN/rRwgrjcjfko2l1O71TdRP5jwtR6tV4Cn4XmqpzKjdMXMKHcY6dyQuV4Iht
oQjoUsla8xlw1eEMJWLFqihff+yxpP9nuZ3hfO9L+QVOL00qX0mqxVpvxqJzZ98O43R368rb2pm0
P5rQafVBYzqqa4d6r/Ll15/droR8z3vS0d6HR6Q6cAxMhz/ZnvBqU62WZC+5MEGi/rUKkXM3WcXo
uuF7RsDcMDTdRFrR6F2yRqRxN7UgAqsSpWpRDwMSwopRmb4DkfTkhatjeIY+T+BVp+UmX8N3LqKF
qIDWAUazLJbxn7vqgFzST3Pf3KbXgOa/Dc9h69VyU5xInNU56k7xRS0dPLbBFw0OsKIWEs2pihbt
3a+fhk/pSnUf4p/tTfs8ygTM0uhQpgYciGt92lk54ArcDU8OJVBCnGf5wFA8cdulobFyOTD7dCQc
Fzu0wDrjxtjsgnb4WZ3svnv6KUn1Pomk3AUCtLaPBMLW7t/WfFQgh8d9qnRzNoTvJbD4XivkRHZ8
Lkt7/ymDr4QIQRIsLTug3ZuLvITdCWUuV+YjjhU1xz6bGCp24JQ70o0ldCunMAkrk4QgLNjyr6B0
vdBewPzlr5+wMsERa84BrYh6BSXsJ8BARa64bYVsbQ/O5jM6CivsV6+nnVA5XvA4NRcdCCFRPAH5
Xy+dYSc2nlRefG2zJAczs8uXb2T8JtYWpB6wF2lqt2mnvgS+mfhUcGru2ksy1By4Q1tghb0+NwUK
XF+kdrTaL1Ka12Gv+8eSzzIusKZG3yT6TmLgWbfTO+0yFy5zQKcEH20caXQwIXk6en6fn8aC9XD/
NLKPMPezx9pzC6lp2uohLULzzq/v4emxbdfEFXFvbaA55WPHTKrPlUPPxbcnj2DOTz9AssY8vUFj
2sWvIFZC6/7+369DYRO9/0LnhIKi7hMaZ5x6tDIVFpKWF9N42LDYXPDckMks1jMZHYc883nnaKl4
D/1llj8hEDLN3ODSXT9Z8AMaD/P8M3UUXl+32k5+t8i4GwrUOCQBOhsz7ArDUJWAUoVr1z1bsmDJ
czswiyVpOW/kq6vXPJH33IY53+y3fiIrNZiqaKILEHbTY6y4RJnLNarmkzYhBZK290vtlRcNjqOK
fm7hG/LJS74e2lktm8D2xWwTdMdowV5AaGxb2AXlIfm2/jVAtlsW01mlDxQP9xjOJq+9gPfZlrNa
nYh0gZv1wGoiyVkYrYb7HFXUREGrJmQT4YAZlMYmXeUsSAN17aLJyNl/8s39Nc89eTSICPd0qw+c
5TcVkEsaiULMMoLx0rcqj3paL4G9peZr/+j4NhHflQGlJaEwd5eaKnjUMIojfiooBRaHg7VAa8Ps
Ea6P3n3CQvHPJ4QOkLAdkqvcYDdaGqyHpR+f8csX1xUSgNvvVE8O8z3bYcR20TF4xkFSFfz3wXVr
WsdgeLSW2vH8Y0ebRNcAAF8LNtVlSRr5dxVNMggvbJWdgroJsHzq1181zt60grHUQJtrESAa4XsN
M5BDvppAbIDkOTamdfgGF8iakfj0o7T4WWgDOdKJ5gbJ7T20/jGyXDHzODEiZBVquosiW0cTgiOg
A2gXSNTfC6ZUklIf0h5jHH146fejzzm8kgILkTURcjR475yP/uJjTLtfQ+nLSOs3vikm6wqvB3IG
GTnjREEC/nxqZBxUymvv+BnqOhrW61ggQp8NaEL/q/P9FZ2mdl6HGx0k50hEOj0XyViIA/tmaYFU
Yos7KE3iBSNmCHaR9Se3fmLCoN6p18RLd1ZJ2E0EE2vWLPN0tpRdNxa6gso8fU7VkTD+F7KJAddN
bJ/2j9jxrqZqFzUKfr1UppOlkFyXkS9RmW9S2GiFtt0Z4IkciM2nbSGOA/8JFfvwnzbKPJOp0o/i
5zjVpwRhn+T2iF9sqWCc6XNE8hP4KSzZGwWwmgHYZECZazx4kraXxWDbMqEekGJzLaqzT7cY/5T/
+oLnpo6xnMIT7yZasbHP2EszNJKgSJ2iX+V3+PrgrJeq3wv1L50girN3Bdlf98VZvbKQ1SC+Pwhs
3srR+XUtCKjVHUMVkLVekklcQoviCX7IVhD9u0H9W2YmxBahAIxG5ZHM56GX+pRHEBjmJAAFVx1T
4eThKNqEVsVt80Pzm8iCx4tUSm/XTYoNHYonY2MFI9AtVGQmRjnh1Asi96H5hipo3249gKFPLnoT
RZR2Yi4hxuxpB040t4oMFTitOpFhBOcZCiVcGihiCgrbH9D22oQq7YbLSS9SUm8PcI6NWztCpz5O
wadPBy8KGs9PA71RgPU34EqE9ljIPsfFJBdHYz2x0mcWI6z3U8ov1tDyLeJIonKILS2cBIuVe0a/
3Xdh96kcDz+KOhykr8jHzt3T1shFHny3GnYJR8TGRJ1SdA6I9+v2RKowfz3aYVs8PRCOpsDIBIbI
wZLH7ZKeTb4XBduZghySAuHvAgF+kx2iOguqVmMqmAim81hsPBeztlwCIXGp71Xedf76HTfWEjIO
SrZIvDSgUxekjAl4zrV0nTN/9HYtvSIjkXoffj+hDU8sKfhPtAwGri+7YfrlN6ycbN1RCI1xmvEi
jSW2e2rDQI0Ku45T3M9BjNV+1+zv6dfOYxvRXxr0RObLxL3YdG9FY+9Pl62SLgx6IdOq6kmo6cCJ
ytIyzNgwjdJ0mfETHXBRwUVJiUmeHZLru2oYJ2bdqRPHT5hrMcWwNFvLsZY8klaot9EFr7lIG42d
cF4RYcs+3foF9HoKmAKVpV5uSraFPKQrUiipe5tZxOhMH6RX4I0N8flaCMJWJmSMDYzcduAiEivI
QkCTOHf0sWbxavZsat+GmVs2RzScIijJyOliG0MRC+ZRJHhVW415Q1rbnUSh7N0usQ7zCEz1aaVs
km1egiOuv7pmwgDYiFHHrlKVAcEKqG3llbn9w/+ivkmLv9zQ2Zle5+kEGRyyv1x8ujhtU4mivBRI
gKvWcH5ETT8FK7Df3bPSxD4ZLmkoD6XXRyucoZZdRbG1492YBhyFAgOD7mSlI7oDccmlXMaBYqDm
t5q4Wr+fjGEwmfVjVm8cQ4DKsk3Su9nVe7G/Lna7HPXy0gUL39m5VXF9hGSQwTNG369zp9DYvq2s
DBoI6oA4ITKJOWv/fvc5O2xPi5m++pR+z6I8zFzWVIi52bSGpTL8zxnO7wvlx0YRTn9EIJPgrRdu
8zDA/SKxUGCVyNP7SMRHYrcZsyJ3QKDp+iSDWM9Ish92IZPZ17BaHdhotAjquY100afbHdgRmDm4
1j1rIdz5aggpXfAtz8C5mI906+6bECQs5KQZ6Jhh6sEYN2E/k+LIiN59MZoHMJw+AeDdj2TlHp+6
5RcP7BiAetzEe97ZYLWCprkBLClO42YTqkV1jlBUhZZDzH3/dGUNM9S+J4X12Y4pFp5fm0NDlVG/
EAHmZfaaWhhuDHDNv37qe0ZL7L2mfleLdlpmemIm1d+TwNiSp2QBSrePGevbmpHXnJBDMKASjuyB
gZJpq0kjD5zYtx2eIQiSiTfOEYW4M4uQf/VoNo4GUawLogEtUxj7rDgYbILxFTOJRqnrwvK6EKSO
Z8dHhpKi7xu0QWZ4dE6c+OM+Z5auyEj6qkmexncqrv4xJDFKWy7cBiyc/c+RKWwoqNcpAeAyGxgp
NH224HznMcE3F14vE63MNRJsmPQ00vpDrjRIeVg+RJOEd0dQX4aVB0tHqjGOemR+5LAGFUderh9H
+/GQJEHuFMKO7Mkmvxbkvi0Fq4xyLFAKLIze8EkD4WJHTn5DOFS+sPbTmNxiZJ1kkMzImPRHy5uz
tqv0xZi4ozL0vQVsDnb1+aPXmpCVI2akhfE4X1OagHk0bkhHf3a6BdemQym3wBxRT34m2fzeQuQI
8WUh1K7wMJCWbWmBpfTLzPHW4LUzhcleDTLeyXLPUjSWgdCKKCxnagOymL/cQ5uN1WWmpm35c1Ku
JMIxwe+NeWL/3IXDZ3f9S/nIYNROOc+5mLY8exER5gSqZJgNLKa8vbatDqjNc3ss1NZFX1L/M6aS
D9vE4y6APV+ZsfCjImTN4FuPU6ol7oyIBehQpiyYlpsvw7KZWg3mR60D/z+FD7G6poxaLsMkAbFa
90AlgI37rR3mPcVeb2twDyFUVlh122TdR19lMSiDp2R8ueqFyLh61JErlGugOtTwLcgeF7KKysNu
FowK237tnTyRIeVf9jOcVVByqzbs0EcJ+9DJzfq1kNRTibLr8vmVT1AJbPM+8lTD3Q6Mbr2fT72f
7PB9Mkptjqd3Q6w+ms+uZIBBA9eceiOhTsR3D+XkXpILUx0X+sqTjpA9cvyYS5jfCyn2e3C9hV7S
MGO2hVnV0dJjZ6IIJ6a1VjhZblUuQfALkVSsbi9scyX8H957jMkninUOL8cVk/ROauuGftTsrfdY
egW1U/Nzoh2gZ6xqhBXBE/4XVQevP06sT3cK/QLcXZTixYQKEGKdg6YdhWXR0QzJvdfXcxkxNFNx
gQ528f8ioxFqLEWCXirAsOpMOFyHGhvyK//glK4kAKXOPNiKW38KIqAYGbXXFlsxtuLWDmC6Kcxc
ZSCi6cs/HirHb4lFf9iZ5tP4vSNwUF2b1+aQsSwcZ0qzwFBxUxnWo005g0II1KetOQ8g+ksppQSA
YTQwdIZlQwEAVuKrrK98qmt/Mq7ZOTwR27dzb3+Uuu42m2ReYgGEsNOd93r0HH/IHgYAP1fEio2Y
Q/x5aJlS39syAjlA510dNVqy4zcTe4rdOhXZJvCajfuVcpGsKYpLBILJsob9X4xL+bz8ChkwH0lV
qTvxS2WM1N2sfKUAoEUesZRkZQ5bqFnZl3x1rvyGb6cJ35SZXEF3BdRVtKalIpxAt603gh3h6sgG
psCuwY3ZdWWN50GQ9tbNKYGL10o3Zif89mmkiPCHc2PzwqoTxIzrHs6E9xmH6dPTOZ69D3gkzlYL
rUD5D/wfVQguBQdIsQqGlQpPgxgkFKAerE9hGtKlEZ4sAWfawwM4HUmuV0JYzO3JhSoKhMPdeDkx
rL8vn5u5uomQh/rZvyiT0GtmgxNm2am1hkGbQzAIvxwFarBYl/uVIsiJ7H4nJPOSEa/hjiweZznn
GDCRfO5GCT+qS7Wu36P9ZhR46bxCgaMGl1CNiK13gnVud1I8WwwlgZbF7sK+UC/9LzGXrc3Yfy0C
XEydeME87T+Yd5yeMnEmEaOEXENBqg3b6TLiLOl4DAtw/B4rmKrqsDvfOV9NpOonZO4l7MXedda9
fw6BiqrLBB3KziPU5wde0Lp9Uc9cwcFVwbQUak3g7xwlacugXQZeaaPDU+mPYvAqQFOTqBDh/XV4
5GvCVtswJJV3SA8souH7OZoXOlN20gJ5KuQPCa/RPTW+zey5FJKjdQ8cE7ZS2TW3Bqhucx4chIo7
iVF5rCP9sTKafHFRCDq0VsChOC101yQlvfZxghrxPOltQbL557Ld0s0ZDYG7ImXnooXAUg1Oj8GS
xAbb39YZaCPkx31D+GCEip+2P+slSFH7eNcxyr1cqH2VSA60jOVhoT6ApXvANevrev1orTXFGipr
T9h/gqfoUQwcnXa2BpRX9KCg67ff0oIpqCBnYKr+AxIw3rC4+7JvP+8Ixz8cgAMWP5Nyvr76zXIX
2bKJVQtPY4wrepoNzt2hX+vJkI4yrczSWjYd4jxOS8r8cRGgvT8QHURr41g55Y6GK1+aLEFS6vMr
tJvgLF9wQKdHbnplicHOkcMUhbk+/zmwjd/6q1xDhFS77a+LwJqpRZmjK26EbFYApJl0OTdh7CdK
Rt6y5ex0lpAxu6duXO/P9s4J/S4Uei6R/XsZMdnSqRcjKiINFvbPvS8LwaX6+zJ+6WPg5uSdUyWe
o1jT8blwMVUuil2TUXJSAwHAv++USl7vGuNzCfRkw0t9iLimm3zB/faXFPElfdZWL/n9BQFPHZuS
jLWUv/6rgBhfBDPqwT2s5nQM5TaoFFF6v5ISt/YIQv47qHRSskC9mr+867xPaAtTqzol0/Bkdl+S
QE9sACcjbpR/0VRE0QjObzRl7pMv42DCNYuDVZBxKKNDiIygPz+MnOXOq5hbT2s2Fefzmvc2qCfj
nyw17SDGwqv52YYeyVydZ5iwWMD66er/xJv0SMXzmz5g5nbWqOMk2J4sq6x4nN4IwA5VIsHyeNT/
F3jFUUJKyBrUNrb6CHDxfJTPYh0eNBX4FJTHHkqICH/CRbEkBgBcgaxFD+zVi8RPNisGOSP7olCd
FLIAkQ+4XYqBKltwbUphdGXNFBSgA3a21GzN4GOG3cdckpahSgtfgLJmYiVxkPbwOxIT8kee9tXo
o1Lv8F/AHGaPS63Pb4S1I+V6SLM8ju4r9Wy5wCvR4ZmVcXyzc7PK7NYtf906ByXC4VTOxk0PPv7t
y4rxhipBw4e99UUJ96P9EHtH5jNQUAkh27DzhSmSQDN4pXa0mipOkAlfeY6CfiAJyaZUKui9cmwt
/CHAJKoyGdclL6QLoeQEef5AtmFFvF/KLVuiW0SROv7vo6pWZ5uY7yjFW3DS4oBgPwfMMJstTj4Z
vyUQeuZX8nLlyBLmD82H6TPn/6BgIMPi36/lJp21yYzoFjy+wZgMrbOM2RRmgM6nAcCvrZ3MO/cS
wgr4rf9L0HtO06ICzhXDFP9omg7eafQVe+EgL8cXctj1aTwMh5gSMnkI8Tzo6lJtSGTOE6+nFWos
4aXW8m41gCll60NAJqR/hWZCVyxRS+/ARKGflm2hJ85zm+CjTUmwmHB2cSMBZ0MzWeXv+OxyTkv5
i9ksibdPCU7MQ5WaAIROW1QAXhJFjbYSHe91S9a3AKD2PrHxVdE+xt4YIKBWFj/Z6mU1o7T6vXOZ
R7X4fY2/JJKnHxK2k/lWwK+aEOEUvsi/BVDac24x2wQLw3KqLtB7kmnXt8+EuhNO5EsVrG4A6d94
NYsIeEGE7zXArWJgaaxCVAmJ8ES2yMFkn0lTvae5KVUewh518GLfX+YtRZN0cOVft2bBgd0n1NeF
SJEzoe5Neg+0N6Ph4sO9fvI0W4Wjwe0qOTN/CmX7Y3M5pV/KTVM4N1b4/HEvvSWPQe/NYyfUtuG0
IaDCzJkh2I4b1GKfMD0cbdt1CiRdW+Q7h6OMWt7sHn6HDqCRpkfwytYhcM6P+tmtWILxPe/rYBpZ
M4yCJVipoTcsc/pXUgbPptoTSPr0tsM/CK1nPNUm+atKIuJkGQAyyYEfmZ5P0dna3OYkRQU/vPAO
S1uytI+eqwRW6j67WhD+RjW3cWC2dKBXBCu37nr33WHtirDdZ+2hOgFzpovxXx8z8bG0801x5eZF
xZ+Tg7gXbDI+VzO3kJz7Gz9PMxGaY+4j44PN6Yk0r0hK0rcz9OUNTnWw6whIYf73QtwDV4qGlQXP
DU+bfJvIdoOiLmfuvtCXHunHKX08p8qKXajyqrSk6fj8rAF5MisRxOav/YyXGczRfNHs2YWsdnH+
86grX0pSxY+/7ZfIpxWsoD6aitFZFbPAF0RHBPempnrTRboKXNoa1fLqsVBogqs/bR/19JSI5dM2
/+GULMatIvKWd1NonBtNHyM81SWgF8FTprTCoa9wGYqVPA7EJ6GJzdIPZ1e/S5JWgoQzSEONvarb
PaLB4GHe8oa7yTagLERP1rOZEJ757eUnNiajTlmKcp90P3Ru0HlpUY/cdNntasqMlmV5jORMscK+
L8g2dgFIGQH1P7WySXHDOClszWmmIh1XLAiKaijN83dpdpVQ64gJe6IOVZQbR9iHFb3q88sO2vtj
aLQsyQCtxXyec/SOd44yZGrlOShtjKfNEMlYcXNe5RtVUpCpP4R1ff5ADPYFq8JXmxl38KZDmQlx
31mASUTbzhgpBPQAvU3poxeWXjqcLp3OXwfCT0x8daczawy+uoY+C/979TR/g6nH+c0mfRKa3aL2
1hWJxgZpdOerR8ZYUOEvqCuYy8HrZMcreBbJ/z3pMuEHOXo+r0CqRckXuZr4b/XoD9vWK2TYuz0b
40nmTBdjgXIz7OaNxbcA9h9GvvCbZp7hFqha5a+L+mofVRpi7CcSkrmFIRs6CfBGELDJW3fdr6ii
UGOF6BvFCwMPtlFPNO1HaZXiUqvjAZZjkIE+3HJPFMSS8F3WvVWzJfEOlOeX1NRWK8ccy3pCbhtE
ype9eLhUDAXOqIfqaqxG7janBiHYdYad+EoOzG0diNt7eD/0hAbNYDLw5rej4g39SfF8o/2wQv3E
eDK8w2Q8TO5i+GKQKUfucVMQKQu9IlqvtOAVZwJ4DtXoax4bJaIbJmxFvP9aCypNzSGhZvNnKthx
8yYOSRoaqttWeIAEF4Q7qgpdJhgsrEyuz555I/6hsZWkSl6gMOh6dz49C/ubq1sPhQslfCUMcbSF
WeClqXTuQK5F2CfQJ9jmsglUhc/CUEB3ENIWiegLbEYPHgztl16KbQjSsU53ufIz9vXJL0H/WaBp
4UXd+MPYK7UIiLCIwBnwvY6OovxDnVkRU7P7Rpj9f2BVVqgIoHWxZE8Uvb2AVbM2IwVbQBtEMqOq
v9xO4TFdEq650Wh7ifrS4nIt2a1RpPWw7qyRiYJ35p/XGa7EId1xpDqLATnTdlGmJubAhxLDnQAm
8Ph6cALD+6cM694vMgpgrtGhsYASkqt6p3R/z61f5fpmRyJPLkcY7lMqiLV/RZBTcxUGi8/x3oK4
leKNf6EIIULdWcVpkGWE1X9XggtgsIw3tY59fsUlwt0Ai5IIChaLjb/+UA8JmS8NpwA0jpfIY01W
hcZgAaxxZlYi+AQ7yoOgQKdc/Gfw4IQZdKDTQ5lGZOo2l0aT5q9nZotrffdFBWgUYVinnoHZ6mAM
fGSwWpbUNkf1RuS6piGqbujqqdGaEc+ScCLh2JPvDQvAO6gmmxkfhS0IyJ82vEUKtutuLmnZVFft
owlQ2frmq7tDoYT4eQiAvD4YXpR6EzFceVezJNIea0KIueciRwsKeERveyqHbE2xqnTn67xD0iFj
SX1nWBAutNeYPYZvvs9VaNYfbnX++z/F6WUgBwIWJZHMV38QkymWDWBibyRFGoUnStziHTkjkY3U
0PydzUjXKxmNRvh9qkIyCfOAhR0FgOHRRXcy0puAPb2CoSfnEyjJIrdx9MZgd8KYD3f/R+Jc3qYB
MQWKsrlmBoxb1oWbtf/1bWVT814Jlx+fNxEA3Tq193j/p+NBv4SrEZmiTUokPIL2EBzx3O3QdNGj
4CQmURpZeCvMhcGOVmC2oi3jnd7DQwbs+9TACNeBvsPPpJFJNK9b2kg7cdCULw8/H2GoLcivgrsH
FIG7qYtgqIHMnXWe+RBq7bl/20P8Ex820YZbzCphQ4tl1YU8KfpjUi0/NwZu0y/V4jTGlYEKl8Pd
46EDbVCnwdixb9LzJYGSorIFwNH4XMqO8gQae5WpBRQP4+5hzTBpgdMPeDU+I7yM7wzV+TSe8/n6
SznNLrc1En1es6XeO+JxRa2FrA0i3uhre6uGVh5MF/ZhRZNoItQybVMj2obazuhuhr6TdUMHXyO6
8Su2PoF2IQXIKUztLJ0OZcAGmAqM1cQJXFf2lvZc6WmUNC9oT7PW6oieOSKI1depMycW3mFAMfYc
N1TzRKL3KcoAmW2iO6opzZqzjPEvVWj9rJWIIEx9JKGwYgQWd2xtD2kQuSUbsCnDnTkqER/+gp+G
FhnmjG/s00tAZqVt5n5rXKHCDo8v2NEkX5UjbiL8/SdJLrqSFyJyHXpFo7szPjEcDjCLQfbD9mn8
2UPvIO7s8hYS16mlDhCjGZ+RGtwgT2remKGwrcWacoi5n3+CuYD/p2plQ4Lo7QRHTihraKw0ILZm
4/iWolaTK1TkA9Y5bjT6H3WBiojvflQwbrGVqBvxr86dAaDTOrP3KypU7wdVZRSE2/srHDjJyVo0
L/IIJBJyws0KU2z4xURWdViKCpUvK7OSlNVfnhjOWezfN3i+mkDAoyKChJC9TcTA/WC5IANu/CKz
Vx/12VlBw9Xqwip2iXAxi0VJzEdCIzEb7QO/sXgixH++GzO6Bdlq+IzsOuJT/eQcf4+GbY7HxzAD
b1q+lUcYL0MUDQaCSzHr1Hi58pgOu06J8yJ+qTr3AiaLzIEU1hzUdU8pZyuBaz6V9a+ABQKOvp23
wmh6FC0Lg5wYX5sMLM9PKp3aHnhjVfWHpfduoejeQNblXF3XwWnKRPdSz9duarxK+GK6ybC7uMVT
EfGlVDFkfaQdCld2KsjlMhzsdmG6Yj9o752Lg3XA8F0ZMgSK+bOVDoCTtNioIrCzP9Kfd7s6Frsx
e9SOKTOlLIY6Yt8yAP74aqGiufqDWrMbM7eMTYKNAcTgVLRWmbb9TSPb3xslgo5OkbQe8i0KNfMi
qoEB8fgZ2gn2ylN6T3VokN3aYQxYi388cksxrHYTcWE+ZMnxo5zR84blmtZMUwCbLdhBCcga8pqK
Ff4e/sn85AAq6AEwVcWQq6MVnwU3oHnDdIqNI7VYweZScZM7R9OVO4exp/uzNqQYSMLjfeMq8Aoe
PmxPKDn5H1AzMEePvEtaeAAd5Az4QxdPg94ypDu012BjF+S+I4qpL/nsqXzbw8g8iAM5S16eNQ53
SJh1c3DnSMVnv3IzbzbGQALXhDM227IUItrkXfmIjIGh+83GscyPWd//Ad9DlMhxsCv2zpXLCly1
Vz2bEnu6nKIHzhD/5iiQXPEvtdHJ/sBI8nM63ySHnDZfuDUEbFVwRpQYxra3a6IM76Qt8J9dWRDe
X3dA1Ls3Mc/neEs1xZqjDQQbKYogHu7dbjh/qaEKZwiafvlqMMXeECFQdl6OG59iGNL5ur1I0DpK
RzgYBt4ux2WHtQ72mN6v5J514yo0ETqIX/P6UR89rMXW8KxLoCZ02sfT16FWeZiVODCsT6ifzreY
kqE3SQgvcHocDjtXK+h+7af4lGipFoYL+IFbeWLienizCu94obZrIMXqcGY0JCslu2FdW1uRp3GH
GpJvhyFZtyJ0AR/c9QRr6/LSVLeHbhAtLTLJeUaJ0YgWriA6L3jUyWBYkHaBv98gm5qrFO/WJNLb
2wmAAC1z8WeiopI3VOH7DycNjh5wwnb8mUKAWStjEQs+bpS4es0JUeKTwrccbQ9ZjvyKh9JKIEzg
LZDWDb7ywc9srK5yqzUYzT3A+Eod0FkDqGdCrTKXViVxYtiY2j9EAF8kRGx0ImIe6KwiCPv8Kf92
BTXdRgmUNBMhGKQHt0/XX4fu3E1QjzR09DQ8+xH20FHFHjQ2GgsUqXX5mRU8UwLKT9TQUOLck22h
3qgLT+vgKg+gcgdYPjQlImQkkXzsXsEH3zAAb/QczLMtMUQFg/z3QDB84UUu7K11SVu1wUfb/abk
gQ5cqE58iToR1PEio8puRtOqiFURoXDiwxnbCGKXhj8LI6YiDgSQzMJIYUMlkQ4HJB0d3gvNBY9y
TR3mTn0zucNLFoXiujR5dev91pcOUfEjTt9m2W2cyk6orhZzvR1PSLZYrtN3z9r+h1l3Ndgdi1j1
4zRNPa6c7D5IWxtaof+eposPhPiG0q1Q9+vNmvzwzLF33ochcZCaMjw3EYon+lui4yTtziYDxhfq
dnZxa+z0xyugyD+PqsdKnDQc84R5sBRY/EeVRGVzVEHd+IzqR4kbDN7uGUKHfablk62gppW+8Hc1
cvoOp4NoPiZt7huygn3xfqmXopOwng8vhuKaRavrNG4girFR1a9VenMV8zKlgKiQ6wZIjzcIvDqz
Meym5GKJWr/46lI0EAHZU2Epw99XOkuQTIUpExgS3V3a5UmTLwFK+2gP3oOxff8edSDHUOZ/nGXE
5rGzzD8IN0XhDeKEUQGxE6ZCttvHjF44PxHaRQMKcDdx3uN8lU1UdwhfSdD4e5LYEi0XAT6C7JIM
AXc9c17xX+CQQJ2dtF9ElBCGkP6ChFzx7oxkKoezf6FvWf5+9717cAfnRUQ3cbwyfiMlH+3nEvIP
qwzRmXqMRFi5ynpkQg1c61xx6N/gr5lraYl32UGCDmjuj1FC+TyYzNY1PzH4WOGAc7n9lZ+HtVn7
omlvpyx4DpQ3AdEt7F6j+/SQLwpWbtLPUZrr2eo1j7bMuFJYyIlwjLWd5lmU+FY4TG07JAK9a2V/
eCjp4r3XfSXsyIy67/WbbsKLqkrBZYRccnOBuv4QLLdHSC9arXsvljH58EDQVf1gPpUV+OEfkz2S
eb1374LYpP4GreVyoySVfte25lhEtLa0GSlijAyaL69g3mpmTjaIfA/0JERym2O82CGmt4j/NflW
45VOeUZCiWQzZ2nQvRflgcFQ65PKjHwSo6KgI/ER+BFFXSZoXiRu/hmqWSxdc5+ysRqMo2VSxvJ7
HLUoUSzH3/IBP18GfPe18cisgKjnfx1I/nM3D5GVVAJ5iHnt3X6KbEBorFBJRlswqN90QmJ/EDm8
p/So8apWKFElkCOMXrND/ik1HFi5soBnyVBE5ozmpm/mCkmlxduOPBU8gnMaCG+nqKGpTZ+LHRvc
xZ3HrdvYL06Yq4KMpIwZguQlkc71V+YDrPW6yh8hSSbGuHfIefaSngsKnyt5KQQQQVXzNxaPmYs0
JpP+JA3nsveIBgrwx+ww8hQFENZshiYHQblo3v3v/aichnq20Uc97IQgg9CB8OIGjAfppbJM6gja
Sitep6F54D4xwzwqM6OAmfCZ5zzTQaNOJCCczjTMhd/TYjXpjWT5g/gUiznBglwGXwbM246NddOE
8HM4BmJHlMpjI//1wzYNUABD0dd3Z1DnmKXEVTgtQaKJPSCmMSNEyBbPYC5vuWfnZxlBTPjWVlqa
Bivygnydq4yzu7TfyKeavm1xoAkCld9I0PRiqJmx4yWWYUNUYVoBejOQSIz0uJ8bQzUYGytgxafl
fhFNnH0fuqqGf8LWtVZpu2TIuwf+6oInvVee0cdr7TYZBPM71ptJoqHEnnRB5D7LazjA6oiydgUL
W2YhgjI9jHXuBS0JMKOCpXPmi2KZ7UpXoaMzHjYSG0WYiq3dae+oI3C5JhxwO8Uc83jMlbT2sN7C
uA3fIh6YF5ZvgFCrZhosOY4aOheIOOR5NTsi3cPgCxDm2EK4ElIqtzfdtb3Wtfsf72yrkusduBLZ
IZJ+mpD6bF2u0vUo6FiqkpJI0pIFMmFdG4Js4gyj0iTyABJbtWXXkFOVepAo/IEqQMfCpSxgPe29
Jpf4l1e27rGyUOrQCKRA0UPFGdD4lnUyTIakHSoK8iFfZuoC4SsCFgK4g6SGR9lMJ/WMm/cosx+L
YqNaMH9ECRfwGcLh2yXb5z0FFG1e/aRk9acB/EUxwEScT9wIdn5h+oj5XQAP5mTyojVWiA/Ny9YQ
SwUGULRZjv/e9Ld4ycePi57NDKnMNDPyZMvkQK+v7YdVEVwICMrEQ5q9Vdmj8TNh+J5bPOu/JFLE
OUzyTkIoQebVJl4kC8eWFjg2++F8fpSx9g0NELM5qx6PMPGtiHPq+JVxwenQUo0S5AtCUVc2hix6
9DLiUX1sIB3gpF6cy/9+BfirMrK++WQ3vPQbmdC8nK2DQEQznnLbwB8Rlwq8DIkrGv5hfbXJIlzi
EvlWIdXfuD5UrDKag0cXweqcaj2TCmT7+bBzS5UY4SYfaz7HG8u2RdxUt6FAVy9frHHlBkE+Hktn
HMkIxaOQ8WyBgdauXwFnlKtUdN4vge+nKURJkBV8zB2+GIrZgRG/H/OsBeZpcaC/lrjDVnu8UrBW
+pIKkuszxDYdbRTvLbsgoiBPVAC9jfo+roxnlopYKuUismTjPmc1H2PVusIy7UM7XI5ym2onSLC3
JBWa8nSbr3M6HxZrY4qlPJacXlFdTreWxmjYk44qHbrTp/ft/tBUj0MvEXu7QHvHzlzxpKYePuiy
1ynYIyVypXyfO2gE3YMix6ryqwgItGkq9vInUPdcIVygAEYbBDUTmWH8codFjwMF+0hktDe/cJyh
xdhwBu7zKjbqjyu8FLlM/gLne3qlp6VZsU26KRz5IJXkvToE7kSu9mBp1ztSpe3YOob+qQowXOLx
/ectH3qIOGexRkGv9uxbTzmpQQMMEbNN8ILx409MG/jjU6lHtz+E7zOh1EC2vu8cye4bQydwTtRF
N7S3mNQs83K4fKtwce3IJOYrIG0jsARKe/DgHymjtRl7mtQww4HHQKCOxWgR+8/KKNO/UiRG5q0p
UrXpJBb7hxMSSrWfgl5fDrXuA5VtL0o5ZQoHW8L0vI6xTwohO4D4yKsOEq+WAePKDwCsDbBA7utA
sFr60NuD4qxlWPEWjIu0fMc3hRpaIcaDWLqitZi7uPS7EtLiJ2kCKXUBiZ9RThaLAw6TCN6Wvb/E
F3lj22+6QRH3fazYLR0vdjubSaPZExGwvTbcPJOSjBpx9v/16mYOjWOoa3f5o/gPNGYsKJK60nhL
X1Cbdna97qXxXUHk7SSYgN6gyLYixnm0YHhYoilktN0q/Kpf/EKryHGpbBj39ZVpdgwm5kTjDfmB
+mVGxcNXsdy/oPVQpS2KGjmeC2+TgJnGusQv4ozOdw1+3MjXz4B6N6zRDaIlscMYaFDRj/gjWJkX
HpoXSAaBg4xL4dvJ3iAc7r5w446cCqbF9SzRF4i53PQ4Xs5MD+Ik+2qN0AnDHQHQfIqktMDeUx2E
JwKuAkzIYW8mVB33iiE5BbhTjDZNCkP66t2nJ0YLpCj74JvYn55n5IgMZvIraR/vI8r7ERvTX4Ks
0GhSUzkB9RLaSMKRh/xXlEn3THiLz2gjFJi7mU4QU/Ix6stRMLqJlSlBO1mxSysDP6z7dEZNx7ID
c2w9rRjmc4ByWuMxmgVGkm6O+2LpqYApgccUpf0xJT8uXKauhFqpYGsGPiFawIS1f4tDHjgGaS8U
QDhXzOY8eoMCZPRpVOaGEPMdWYqxNmvt9i7PNJE5B04Ti56sV+cuWUiN+O0b7i3bJ0vPf0uAkIfz
6BYJ82wEY1kwNbxsFZ49AwClJaripFfQHpaU9BG1Nx5LKx8CGbTTo1Lu7w7T7Rnn/evZO7/zsX2p
VFKBxSLkzFNwMRRddmUoZDxwh1ZkYJkYNY8mGtJRxw7B6TXG+m9L9meSVfqezC18OAkaBgMTY+Tp
cBRs84Y5u4eWF/tqT0zlDUIV/AZGx9Sup1vTqRcbKPRlYtMB4QrCuSA5htpFmaTs+3bUX9xqs2ce
KsI4jQxuNmiVX9jf6m+kr3Aje+NcFTrKNodVSY7afqj3yl5pCj6kRG4v3inBZJx2IBTGYkbKTOFC
LAMRx6BoiRZGPnN3kKf+DeV6iYZCrTSk/EYjxGRbXSjH2sWYzhVFfmqnShhpO7pLyR3HKcuWZLzL
khpAmEI9wbNzCIwndw4C1R0DDxnG5UDoyFZ7dHHt2k6FXkWFarQHqsa7tS/NlI4Uk0V/qxa5z+sN
vXCidSOcwSCa4WYDC5Jp6a7HCfbZ/MupZ9sccrD6PBv1p28txoF7Bg8VzuuPsTpU5k0ZI7P9/Itw
7mwghCeVo3IU7XetXSuOc0rX3/9gZ3rn847yGcuKvAIilBJ5B7uwpBhni6zFbFSPlXfouT263wA2
SMRlqYnXfQmJFLWBhTjTzhijyBSP6NEFjfUQzyC2BfNjgDSgysSOXZjw0aDOcF4WTzSRboFnVxx3
z3twWlVAC9P9xXvpOA4ZLQ/L/tUwm+VTQHRrPYVlLcc+77zO9BE3wy68kAU2pTQX7qQMvsieXdff
H/K3HUFTzG4zGflhn/P6mc/8PALtnjI0xlJ4iS6xRd59oJLlJGYoUHpPq+LLe2UPeF4FIvvHrnG/
PhK2xVXN+TjaqEZV00heIvCVfezoneBfyNHb87lzSJr/70P54ljFMsfCyqqa1jPGmkiv60kG1pIR
Gk4S+661ShmxWP1VstDfX/+a5f/LYzkHA2cqJarVQHiqGJJWP3Sk9p32fcHj6z5PHC4jxRlsPrUr
sbqn0wIv9LFi7kUWaQvRr8ndjeaeeGLTYZrGRL5T1mtr6rzj6ZjrPeSRRoJjucmHhrbvlQ7WlPXO
gJAnrJIQ2+g+RRmabtiEq5RHtxyIu5pii4OyNnXui8bs1+E0DbffXoEdpKWEey522SHqWTH+WuiV
CdE2Hs+hWfVrVKreZhUen421kd8MT0oKB6SzwtsdVhNmoKb1pw7IH5WquDh4W/63tk8SgGipg0sG
ifZRmLZgYwb3wKlGfCjd379BBC5cnhTdOq8QKsIjGcEpwg5jB/iK3KIVi9BqBItrTkPX/Ggtb3G/
ByCjh/j/ErJ7086qgiNuUoF1szI8RCnTB548OUP2QVyoLkqWfddZBTJ1hoA/S6pU7R8rPHy8uELJ
Y6lNmpBFL+JNHIPVj937kEBHywEIYBuhk/8LA8GzRSQgKHBsxXmcRcsgmtJHmUlp3n9MUQD3eFRn
Z3h1R8nT/mB2//64T6X+h9492SEgxIOiyNB4xqLaR2G32CNd2L4JmIKLthkd3Kp9t9lbMO2pCGT/
I3QzNdKvd1bEnmheTCiqolMOyLXt6zZxQ0zTJIAS2lPM6IPXAF1FWdlvjkLlGs2fZu/twwbqg4Mv
u7MTv/wM8YsF9PGoboa/oqXi05UJ6vTWCYM94ijENDF0EZbsCDieJ+d4DBOSjmaV8Ua2b+j4704b
7D9A3QkPeiB24wM9BwWN9Pe2sB6LxtZWBGrPN2uMuS7m2KhANlqmIv9PIIS1Yot+NkXQrTsfxoBg
Ei195OBLNnLL2j4eNVhp09wREVl/yXGn1LFYO2kbVCmL6VXZ67fYRdZYCuW6duxIJsDp13/kK3yl
PKmGvPQuY4wwJ8eO7RQXl2oSLxp8Q9BT8A60jYd+Y/mx20ndQcrMvESBUW3vuduNAsfBHno97W+p
afj8N0EZg5ZwPPKzt2BD7pHGlu/UAg81k1ndIaSm4cGvgR8IkofAv7+LbpOWDTzmZ0Wrt9jmgQ7d
AUTLKtQ0moRlh9R1mIJDQaYgpDQ6ZMOVxH+Z8uwDM2Q9y3TQHJulTWoc0FtLfSrgQwFkQmSNyGU5
XwKbEk/CNUgD/VV9fXHH2scYyHvZiIn+BBpTEWNLtBCEY+Hkh46abRmJhyl1k8gJTJrpeAgpCyGi
/v+mfabNei2NxuerJy26HIP95BJsqoaF0DQ+nCwgIjGRHEIQ3uI0GGi+Iuf9csxrbLHWjWigESCy
DsjdN092dtnJE6+pa6xxqIP8PHQP7OvTDVtxg5LLhs65cfEevxHZuDFW003nGmd1AMOwM9/JGdwZ
bw7YtyETj7MWCFMbH51mwQ7bWR3W5DhXDDrrcsqp6d/MMVSdvOvvd3YS8JeKXGW7tAdDcFRSdOBv
xnzsWJneh1jMiXd7zm1svsQfML+BjSqA9WlaTT4OiNKBI6VFb7depqeMnuSDI6zaRXFX2BABkZOD
oqmh2RBv7za6tMwhzGaLUaa6uXsEuPK9tWlcPC4WdMTkIBgUPtQ6PBH/AXJ+MGqsq2ag6oRo6bG/
OOe+cM+u3DirKmYgrXMF0cbYxnX2IXMk/gKX0ITUEcJSBUmwGVCW2A2tVOf/r3VMOJFm/xxLv0Mt
86ap47UB9Lnp1zpUiTa5EwR1tsuFLhaAUyeb4K5Wy6Gd8pzV0OYpNn+X3+O0U5ti1uz8zv8LUtXJ
xVT2Is2gmb+9zcyNHUHtxvWPCjWMiV1yOs6oi4cNmA3Gg5TBTRQFUqnN6YxZG6/SYlQSmPo90OrZ
3mS9xrHLPd9yzkhRc/+ugVrlmRe2MSYcD4fOAgjrc/IVSe4agvbGVtcJcpNMmqYkZQLg3eZDdzKt
S3mVUzAXB5N/FWrSQdVBhEm3tCbjibAzOQe4G+lKHCpjpNgol1wOZ0KijotH1ZLi9l0ZD6stCPHa
aq9AdoDrYi9FbnGP7rZK5OUK9F8kC3t5baiEgizArTJL+LZ58Mre35HJbwgLiyYPRpp2+lcHiJVH
a1plPzmitSNrT6PJEXx6sW2m1YKLADUPkaJFA4q9ceWpz+JHAZAK8EiKZf812xL2+P/chPEtVb/R
Ai9DaLoSjw7Tb/sSXBbX3O5ME4CIB6pulvfE5+B87GXTr1Tsqf1VqZU6RMWlb4WYdO3v5y2L0PDF
bi8Di66nut2QxyRH6NtmXRORkBBEF/yOGVnis9OJ5cavHocw190RJBL3mxlGFK2qMOPnE6Mjc5u+
kKT1Phu7/7Z1z5Ie4JYVqw/NeIBSS1QBzZkCx6kpTXJx78gDuG3OGBL1gcmBRdc7FGw4WaGam1BJ
QGpknO9PEAVH1rksG1NAwpsExf79d+6/+aInDuJvAyPFyYtc5DV8/ooPPRPVjNgw/Ei6KKnpNfxt
CNUC4R2raskgE8YM1tmaDmD8G9ZW90GrjX0HDSH5pTIKeAyV8V+vHtUcs1vwEopXNNpFk+lVrVQR
tAsZyLspg1/8p9t1tPBZf4kP2vi8xyBYres3Dy+303sdLXlc5UVpgop4l5vx0offFCdxndZJuod7
qTVNsy5u8JD3O2GS81+A1xahkqdkxrF6ZLys+/zCiu4JFC5G2DV6ThqTxxeRZ7l/B7XJ2v2YuImL
A78V2UxWkgWF7SNKM/fJsmkcBajFBq/2RLYmTeRm5YraYdxqE4kcoKtDZdvUjYd085tyc/d+lcp+
jbGs3K8xIEiVoYQFJOPZIep7d5siUXbnh5XCfBc3wzh+IezrvYucAdr+2kN51FaXom2PLBz9vS/C
BaCF0d6PmXaFItq9dgheNaEufy7lNeD5d3ZOTmvMChr2MMrMCELXerYVOsCI53CW7CcfFbYQAGFz
Ni1fflxP0sj+x7m8WXJexPjNugUuyBeL2w7kJwRjgA21aEsRNQfLhQrUPLclHEVL7MRNiM/6qVwM
tB+cLssnUk1CrYc2kSg861eqZVAMkEtNS6evi0jNa+g/vDFcaf8bMMQzgv8vtY2YUqqEYJ6jut3O
JocX2I4CYJOPWSYgf71BBaw8ghgTIpQn/BLICrcNfTt5aU6rRY7AxitEGcYoDmXzqBDg2vfBDWjV
/xTWSLoEiEXbaUGbnm9DCcEgwLFnrq+2I/kEo6uv2RqbRUXUI6IjLJj/t/lSMTntfgUrwGh4uuVb
6C73bNF6xhQ6f5vgmxwCkscIo7ZDJVuS3kNsYOv7wwc1miDkDi1ANIpwU4a8WHVCuYJD1mlJhxM3
HCSXyDMUEY1K8+DURF8Gvgc818O9TKv46xce3HBNO+yDL5Wk5Xb1I4lnggBYEw0l/+RvxlxedR17
QG7pJb1IP4Jq9/Q+oq99QmE4isalqJv64Vtcqy+FM0OZMPw//jcFPRAHmS+OUVcyH/lo8tSnGrGx
TAmkgJjteVmvTl7xQy+5CcK2QU7NqjA90D83vC1ty1YHSgNyIIhdVwy3hbKDc2pwc0iEwBFtw8A9
nzsmOVjDESXIrY2zSaPLWHK0SZa1k5+vvAqrTNKlNnlmF7hZaLakSKhFW2eaCALd42zZBgQ3us0o
/3oSjoreDU+fsWwvaUAZn5k2b1ef22VH7lel2dFSgmU2DvbGbpffaXtOZMxqGEmkqfnz/kyT2y7N
nZb5J1AOeaTQtfm+cLq9ep0kBM3A2IbNBu0sjakdwOSZt388HskGXxwM+6DB5r4y69sEmtT+ygSi
IyK0UOSD0CWLbQNRZ2DZaxVo4trKsBe9AALl6H17NU1JEGUw5mD9lisP2/Xa1g4tKSt1xOUFPcdK
saOjwtVRpWElTe6PNrcAUk6f7fLFbGgiF8paUCIKIOw5yxP0YrJ9A+EmeiCzY66BrvOsx/ZotIF/
MmCUwYxdKLQQGgyEEHaRztZjs/sEWy0T6hSryS9PJU5kg08N0XvvpkL4EUjRJeDp4aU3dL6RS+JD
sxT7R1feiscy7ew98XVsOkdwh4wTpU4A8hCDgnhttuNlEeFSURd3XYvVjWp/2gB+Pccr7XfPegPG
7lunQ4lhqaG6eREPU8QLnr3Ait7kWQm5oJkwmSde+gA4a1DSs2jnEGsWQcBVmftOjPRTOxGB2D/1
E5VY2jJj/XpsUtA4p8jPQzuAOIzhku7iEfvFFjxyriSFn4NQuOESqGTrorhx5g2WPNmV2BuxxXiT
djTdZQAkysIVQc8KAPbsoPy4hgfKdYXcpgDGG4izzMFArMKBKPPYIlFz3cGUOlzgmnxFWtk14kzo
Q1kq6lXXIwe6cf+D2CUEOhI4GHiWXA4rn8nehpcLFCUtTa+R14fcBUiC6lmakkHEmQ8eohpgXU8u
P4WPAICb7MVj8Lr3iEZ6Z3y7kipNjcasdB8Pj7V5+FLPrrgUNmYsFzuUFhzo7331ZGRwVkpOxHX3
tyRNyYY+YyyblcCHoW8W4tx7RAVZr+f3x83F2DZqKsvJOdl5NoOMTjXsekKTjoUeCOhinJDfeDbh
VkQEsX+jbwsE5VqWidqgxXiL7lUMhyzyqeoxEM5/UlcrvNvcuNe5Hv0vXpJtyg1MvgT73i234dwE
wjErcj9qhfjAqWmz73lpWdjxWe0FFbJhlfm9QmJlkq/mOKReA1LbY7Gm15KAhHjkwaiiU56LOljZ
nYJvQmmqinQ0ZbnKK6EOGImiKD6gyP7L4op4wTdDA/vmQvZhnf1XgbJdih+m2FHjZ54TxoYC40xk
P0/yphceoGwLbWkCxhqxsr4Cfu99I++EtNWEjdXeEQa8e/eb9r9oSQQ7KbtnqXiGBSKptOqgTki/
H1BAE0NvzGX0j3GyrhmvrGR1cqlpimk7NthbcFVOIbEWW5K1A5XTaARpnKdccXduW5YNcu6DEerR
+YcJGd0g6xUMBOmx7Qcp+iieunMSYqYkYioH+WK2xBPNYso10OenJZbnfDOlnCsle5qEtLgIt8KI
aoSljXM4fG/T3HooZ/NH8dnaQ8/TuOlZLbb8zzOQuOgIP2f7jJ/uq0LH+uyLehMMSMh6TWrBQJTR
JK8TJ8+PyI3oowjVT6w+blS0uWqdy9IHFPwuFXhnznRI+PW7R/34UIvo/GCOCJSOU4MJeKLKgLkB
AIwQuG3SxdHxZjdtFU+yJX7qwgE38yyubZ0KSqWIi/RejjsJvzW6Lo0N+PUKpEhOHGQ3mra1aQhJ
ehyI1WUkmKYICRmkwY7Vk6DjnHXtquuhmnAVLI5n35Fm4emJVMiF3SVrB4bgFefsOY454UkYZ8sO
AsvbfRIJjSyisE1RES9snfNANdSnYCJ/6qcFVlGb61/W7sro0bWP5PFmcABNMrZycfT9G3QGvQF3
tb29a3I+Oj0/JWnVynkk/hCJ+WYD57byvm1olfGzK2Mzp2ZeClYp6puM0wFhZpKbwLPOldmMJf4w
r91NC5/EoIEqbnLTQfb9Eu5JxF6mtYhf1rv0q5YjAo/1rD/iPN2nGFMW4/n0NClfAGuJ5F5XWW4v
U2zwhPaVUZGKA9+wfvFjshzL6lJ5Qw/+nN3ngH3iXO2LYLz640SZfXxLHFpC8PfWRd+bqZW0y4h1
z7vo2UuLHGaeDCeRLr/GBlat8M3k5Lb5Ek5JYH0K9LdBf02XFuT0ENDxu7OXDM6KS4l9IM86xXQb
CYrEeqgU34y3ffMrLyjwM79+HD89m26EVGXF95oiLlpXmZi4e11UOxpFnN/2Uh2yoiJEVVxhdi4n
qXeeFLQXFkt6lBhnmiwVn5l5FmE0r8ADHx+PkaxDRnlLr4Vu+YfkSjFibIjDFBFoHPBIdgLGqgGS
GLp5Xf9pWBmePQkcBaKR38FprP2gMqOPmXPAVO1mZETd7RbaeprUyFYM3f2VdgCnrcW/E+VdL5Tk
/gzqWYj+yY0snWw1/qO4nnwdAa1V8QfQqQThpv6pQS3BikOtkuXXb76wU2LhB52ZHUaBHa+nbHSd
i5I2boM2gqM7IE/PBmtWPpnVVyb3N4OnnNiuE1HDFwXcD0ecqppdlJVUmc1iQ2NEDeUAzKCoQmlO
s/kqVWl0brQT2Fk2KH3C2sMjIDRY6jzs8PcblxJQkpzJzLjfMHbpKQSweOgdP1SanWLkrQEN1ao9
iQQta7Pe+NwAYOU52xRhVNciNIDMQKzakizwFcI+ZBMd5TWjhs5knjSmyM11bNSqEsmjWru8LG7e
Y9ReJsrp+MNHhe9wJv7Kcq26E1caT+vDYUK0YjDZ5PHmmBgJxU1LYlK27+DsHl0dyTxpA8LxYgLf
cF/ckYnI6+ZTZFxIoJnD2HILTUfR+WVIowcO6VkAEZgYXNNvirG8DZ4xCKjvq8wo7ZO3Im0BtQvV
BycBripdC94OZDPPKZRL6gs7FJ/mZsYAOs3wh3O6ZdTuoKHfBRixz02xdKzgLtumq1I4j+SJjCB8
Hw86+0YuQWnWWkvecQ1yXKCDDKDR65tJxJxQafss2k9Ido+HApDZbpcOO86M8Ljj+cr6moyCeBcR
KVYic/Peudp++0+vnopAepj9SYsIjRKnGqzAoddHBpqPzSlxMRMpUJThUYo/348XBbuKg52IE4Qp
kllyQsbyCjR/rhQ1L8Se5xY+YKbV6CAy1s6CCKEsGN8GGDdnDF/i3/LbeVnO5lJRFdcFuQTOsmPz
fA39RGVih222+GPnfL2J715mCXxNDkWZcodymC0hIGflqOkexDU27j9G9ZpPTiJunRlVpQbLA69c
5cxfnm0Il1WHppYelTXjelaSaXlsb1SJHtLXIgX/t24SPH3DpClDZAUzO5hbgIHApicC06/N0qQV
hLrN3NA4j13HY8zLuU1cRuvBrrY3RM8dyaCfpgQ/ivmX9e++wpWgtAc9J867+v07nI8cTRGboaRW
9bQNl+UPc2MT6hFLjMtMUitUhyyZXXg0pnB98+vykUlIl888mcj8UWgdt5rT2fh6nse+qm3U0mjb
fG/0avEwL4yab9zlQuvJL0IwZyKIo8F9zcdNLrRvHdRa+va3MbHgPoT96J+DvFKF90xDCIINyjkc
9wZJYPnyRvf5ynCPL0yIj6/pZueO/h+c92hkga1JMjTMFkY4lmtBo0TCVf1he/EXKhXh6ZgvoHlL
lYyj4JNNToUz3mLD2uG9kmwzwUmo0kP0PaiKXo6wubtBpugTmFQaKQFfKROXccemzeGyQNTNkQAP
nrgteClJD5Pt53aM+jzPh4xPVvJ/zB+0h14YBh5JHm7XZa0k/ztKnQYAf2hpkRBZgOJ//BjW4/Cn
svrJ9pxhfw649vTPQ55Wa/UPv21w695yLNwAe2oPiFSikIAvbf+MbqR/MmsyAwTHVMtAeJ4OQ2gx
yD5XIIjwpqvSEU4ssCB8p3gbV9m/ekFCyBrmwswaW+YsWpry97mTxCtonvzCd5ThIiTSW8wIiyz9
icc/AtJC1rS0vaxdC9PgSJ4I4zeZvBPrzj56l6L+YTE3LicpO7A+bDU8NYiI+rchMfiNHsCDJRYv
ICbebizvloyu97OXCplW54t/Tm0v6beisNU/yM/BTVhR8Gjn8EMBlyJq+G89v24EmnWXrR6yXGeJ
/rH88AcXzZQ90YPWxWGeE/KvGKdA/rCfM4PiWtef4/vgDpit9QPlgohnkzw0zkiAzvQjyX8XXAbC
o7/aEili2httkYmymZ1yldexp4eFoIPr3cJFYrpeF2R0szXUiLUBp6HUJ72WnHWylMh7L+KzBs66
NQifB2R8e1NpL4aFH+zP5tUw/WysZwMpps55tnvRSoIxAZEAqV3wIPVcccLWKYfKtOEkdw09Knwf
wcoBHaftEiQLNrrGtK6Crv/5oAkzyD6UDwYwmryz/q5Ebhw4TEsJqJ5+tOzHNA3BUiAgfC8ilAbB
iWqhNQ3W8CNDUX5CxU56quahzC7yMxF2T0Ehhig6ClMtKQRL4RvMzoFQlgxD9yzcYmc4b3h00wCm
DdhtMAOdR8dkelkzd1k8GKk/UqCBUikz4wXKUPC2wyJaLJ6DvGMy4+IrA9jrE1eTfQ+ca/qnVM4X
QmkTTM4TblU4iMu4l7PXsQ1fxEgMs2p/pHfN4XN2m8+K6BCTp1QnfomMAVNz5FaixgRQ0z7HxrQB
3H59kPUBj0M2FIkk2RJJs1aHr9rzGzqHzv681e3ZrlkS+tJ3jb+hQq6zDL1UzCfwITBJ0tlX/5pE
ZV26H0LC4wWcWEb4k5BKL2F/UiOiKRqrF3CZH81oQvks7a7xf3QHgFc+oldZHfnwq9P2AnNFAHbd
5FSJRaO6j36IQTqcGHGO6VK1PY1lADHZKB8kcQAGCaK664Yxuaaq99htFWZVGU08TgIuWRGledGg
Va1AiwFMHrroFdAQkuc+kSAXO+lnmaeGGztEXRJtyTK8laAX+W8hE+hCljckGdA4jmj6Qn5WKafA
OV6e/aLFcywf9lbEbjy3hkiNDbY30cWvQGu/MtXzBqhS9MLjhvbqr5gP6O+oqIakChu1AxIZyzqw
3F/uShVuW0jJsTEWnLNZrKMOMJGBxaf+XOE/KYybvwkYJC+tnO90cj9LQWAI9nnOzevxyIB33F6j
MwXv2sO5v+rHydLgJU7mLvgS7IKRPXRMLg010sVNpEKsmqwLgB4RO3G6kFBqlbaxPhe/QxUiR8eX
tfkeBJQxjwW8cTYwHAEfg4I4kHu36pKJG8Ky/CZSK7HYf0a/NCbSdYsXweCMghIx68H2g+RVTqA6
JoPGhpUfDijujZgftjDxRny1ouuG0v31oVpbIFYoz/tuli2uIeNA34ZTlgSzHPXoJ4QAXa/F8NqJ
E4b6Ity3x7TyUiAWoHgjD9fWhlWT75sElebJIuD1QlaNweCryk6yakkr8M3r3Pcl83OSsptofCjv
N9sDF+iievz3/Z67szTbenh3epd9J5a/uwC18lfqYDdxTRdV0pwZJDavdElhq9uKCVmosmmH9ASv
V1jU+FDdCmzc+77HEjmk4i5BHvRLYAJXD03OLdxYtzbukUCsBAzhiNj9uDuwI11BNw/+8g8HlmTI
zL6NbInO8sZc5pjhLryQAAf/hwBkm76tFEctPSRnbaf/2oWeGNNp3xV+Zx9WbkFIkmvX1REAoRAL
vfLhc6mQoiZGFxHbOf6jP07DZugCcjWWjJaR/mr4VMnRmPYyBN7OAMhfZpHlVSOsQzzS2W5R/Awk
FXQKpGJ4vpHMkKoexcy08q2LOL3RtlD7rNc6hx4Fo5HNS/wdWfZmdzLYS7BfvwoE2J1eCIH0rrwI
yUvzP4l+hO9SLb+BdX3BMV9CKSvNzkLbD41hAG75U1nZddJInR+Kxouq/EChTpbdZGKHCjuNC6rf
BSXGzdgrb0EJLLGMJkB2NrCDgZWQTSui27P1ONTkm7mp2h6asxNwN4coiG4yfRyDIjlh0IDdkW5G
IT82dwWTjKgyyKyymX5VCg0DnMm8T4kJebFQctbLoAGHhe76bN9zYQrzXmGkpxCpCwJYOVGPuXEn
S01APlyZQ6NUcCfD7iTwPvhcLRbkxfL+D34/vsGpVKMASGe9Xyndm77Aqw7S6/OYRNMDy9VaapX2
2uhI1o1qkZB67UL4XIH7g5edt/b663TNoLwIG6KMlmNs+ks13Op3/FW/nIY5n/YGv/Xqs1S578dg
4NAW9Q38abvJ22PUjx9DKteVhZ99+84u4IxdFlju/2bFGwPvVBLpG+WhgZM1YiTKc4P+tEq+NueG
pRPwn6uwY93cuApg5OzD+Of6dBZ59SeMNxrHx5e6UajLUBe9tjbBdO2U/A5Xw2myDSmywYZox9lr
8IsrX4h5kwL0ChclzRd+tT7I1T3/MuU2x5JRNe63yOYE1kDDqoQ/GmtMyU8I1i2eWqjXt0OnIacQ
pzb3V4Zapa8DTpo0J6LrerWCQAig5MHKpWvvjg8R40O01nqrLjhGaNEAWcMuh72zVTqN5kNguiTH
gZrqw3Fe57o89sBLIGiW2T9pGlob+PjmAswMXK3THd0Dvxqna2JpWdXsjdC5krXv0CcFjqbAazI3
LLa0uRlfNeSQ2cwMXRWROGuYxOsqOiPzkQK28XqW6NA7msxDvfWEtPTxtaUlmrg90utfB3ap3Amd
+F0W79ATXu0Wtk7AiRqnWnjZXZuQJmB3rDXPU5ojqxQj7PLB0Nz0X9WExx3WibUxiBThpYLZ3uld
PRD78MNpfJv6I1jxwQiMOLzwyW5b18JI53yscZWa7nrPxOdT+4ShnSplOIKfQLnFlE/kC1e72bOD
GQ508DABCvl09jhnxwWSdRUk4uqXZr38OcWpWQzKpKoJ3PkieOB+SbmQ8QfNUsGMzNGhve27/fNn
2ea8J8Ey6abRiiTtjL+DjGw8YK/pdnRk4Jp2bG880hFApDQ+4bqS2mC97J0WQClgMDIEW8nKp0oR
ECVKvr1XSemzB4s0xtH39fz2B4t+btySguh6FJVWI653wieQisdVPi4lT57d9ThgPQdA1z9bIqa1
zZPZujcJs9MdLku63SZ3PQSSCHaVA/zeV4EAq3lxOMJ0fu6MXndvhZ1o0vwwT1eYTiJphdOOT0/q
CBDZFdzpfJa2hstTv+mufhScizD+vHb3gPw5jpbE6D/pFUDTHhGiJG2ww27FxIK9y6sNdWdBrW1H
/SEUJR31MtynWQGzr0SiTeg4qeWjVHkEX6ISghaHgvIzmXKVyGBLFPbjUddgiyno8Z27uEg5Vnus
rvIm/J8P788D4nzFrGbowAL2muyzo1zxP1nqAZjPsM/BjmENwTAtvlDMC2bD6tOapt1SB9wpqpau
cnzqdN/d2BEmFXf+f/rhiT07KtMDm9hTVTCfar1ajhpyAApg0DvQfMr9HzYzXMnBxjcEhfftweFU
0POHPYHacMQT8zn9NoEnSzcZSKlQmAitJ28Bwz3eDOgwfX8hc8HhL28x1KYHcr7ZKKBQcvXFzXJ0
aUi3XQ01efIszABbrNgNo/ae9y94GMIfbk8SpOzav+Pv7f72lHDDppZMZy8vK9RZIQi8LT1NOByB
btwYvqIhm2w75Oh/LWX7WGMN83mkuL7Euv/5d1Byj6yTds3sGS4yUGbAy7ab8fP083T5dhD7CNSv
I2IGJJoNilTB2y96N3Cw/xzvfsuwNCe8g3Nm0paEZTF5UAdkHzvxX/YtXUlXNrlENv2Z1i+PyeJ+
jZZvYrt+botbJvHweDn4YXPDS9nMCjvyuOdOtLUwGnRH9ugnAiy6ebhAL5+3UYm4LhFNVRcZlt5o
Ouy04c0q2sbExUsYwPZz8dngtPi9gb4ljnEiuvKgOSk0j0Wg0Cbvh1EH7wEQKa1snmUKYz1GNXUf
iReUK3LERtMZ85+OCmEOU0Vn57yL3WEWK9lg4ePQxiHlS+7avrysCqlSPqROXlAGrUI8Msn20AQZ
tAOVGSXVJAZH2S3KXNOHwa9Xq8LasW8xclNGpn6aLTnLvoPR0KxTci117rl5q9QbbzJaWdKE6+xi
HvUFk6qdSH4EzpUZ/MGX4x0WVE9AOEWcGwckdcrexwV7G6Z7H4f3BRNIimgbt9MPrcXnYk1Nyhxh
5OyiSSFfgBRbifd+W82nPYszCwb9Z/GIhuKywqOQSQvuEde8bfeeCCE6gavjFJsZ5u6lKSUAjQOP
WH/skDy6xF4mXH4LXhLREVNdSKccUVgJnEHQQM4xpkQhCqR8WcnLRut+EOECejubwBDz6qiiQRIT
SN0R4nQNbtW9DJmm009aWgG43WeC6CeX28h5EtIsEzH/nqxET0shKgOFZbMvJ/qyEhmv1hAArWM5
21ZjqOeWrHOtKPObvBjqml+qpTVHM6dtnFrZfhptFQqjvgcfBSp8etQKNylOYIYAQcTkQeHAyb9P
QeYOeiOYCmFNVZWIGSGqZCo/lST2O0T5nKplCy74a7wUE/RFecVikJ9U7xf9RJsaDlfA8OsWwJni
RlL5IRATR5GeBBzIHDKAG8WxuMOxNbX5EmT+lEIjZbxjkJ9hmrYjc4WXAHGTcrryyKgz8m5uc4ct
HA7E57VdevW1XdYZNHi4FuLkMhuyWwv6lKtNnohytBtm0D0T4ba9M1IRUeTehw+jpAWv7hRFI5He
oEk1/Xa1/Bso49IseDbPbXfcPvwGM75fdo2uLqVIQpMe+9YNyY7N/ghTZIe54nW/p726ybpNXmR2
k8fmmnWwFuKEupoaTJbXUWe72PQl7PyAlnrkzKTCmirfwiC+12tGVHqhA+v1eC7JpRy7MDk5WGyh
PoCZZq3yVSGNnAfz+yQycSvitasYL+JukJdk7vBvry7oJEvqJhK0sW7CR5Xjz13RaID4exDZKCBz
CAExt87wQkuF3ZWuihj/nEcYsoSpSlZ+cau1Xrfwe0kxL9N++JMzx/iqqIFD/HxqqaQCsWvHu6I4
QJim5VbNsqtkSkff4W0Ng+XnP11POm/b19e7Fu2A6RlTgsiNHdet94PJ3O1bCDtVKPDA3QGEaAE5
apDljI7Ho51ZfYy/CjCBblMZClHYuOv+vveNa3N91GSiMQAenLxgId9u9cI2vAmzPeXjksVol16i
ih7v4ThFtMPNGbm6XB75vNJ1x8NnCkUBDwiU3YIEp6DCyujz0YVsFYAZHtvlyvdxqdJLamUtvLKP
HWu1h4gu2RiFAqxPiIcxrMllhfMrEFDaNfTdkVjzBPConJZ2xvYnm4+If0R+jhaCoxR9LzCNj6bE
FcW2SzpUQCZj3YxNVH6J9xxRXUU2xSmBkCm00CsVejnQFpEeWiv8IM9f/EuV07ehIzvCR/aoh6by
fisCR7ce2pI9ugXOAiha7ANjVtxYw5WnSCoMH27aYViEpzC8QnaF18znb94FV/FI1jF1IhdBqAA5
312fRtXPYgkikZNTiWnMuNKM5tA18nzGWzgEcKTrzW3twOMRKZ2a/MNOlKnapGYjCakltVAsgHIq
V/Wzesdi+/GcnTDQpPJO9aQMiKFassGbTsv+6HTOTWdYKqCGINoFcoViOVx5ePWb4uBFWbAHNhW1
+0LzyJQgZlIuYrkgJJPizU+x0Bpiplx3dITVdyoMkQtpFSDHUAfP/r/BaOoC0qBYUbTKODA5ZoIt
Acy6HyRCslzw8yULzYy1AJdEo0RGjYGsYk7Rxh8OuW5lHzpL+OmJfDAZT83MGjq3Z3/lQkzeOTvJ
CTQbfFGRdqtE/6w/mFGX+GVibbaA0nNUOtDDrgNg/F9IFHDn1ilijo2YjHLpODwsawyvu+BN4t5U
UwcU/CI9fdA/BlkAVbVxLS42w+xvmB924MwOJDi82odemM1hAe7419KkLjIJzyt9NRYWxn/ICUUg
L+EF0V83Wv5c0/KAb1abrC2rGrMwBeM4VQvy9XZ9urw6vYN4NsE1p2r6g/wZIxRAuPRw3HHxh1NT
BVg038pxCjYPz9F3r9S7QCZpqSxhplGk7U11bWLW7sl4mTLp4Gzt0of++soMSZNTgRnKIX/JdQFx
PESMbx6Lp4OxDl4xOcNFCmt/fsuagls7YtZ+by3Z2InoGzThZhkI9C7i3ZDC8qQnSQKtq8YFlbGV
DYxHSWDa9yvSPWOuWefxSqNbmOXckgG6t7rnUlYMRz04IlDMUOg11otFwuLeJJPoDMrcuY9QgeyQ
tUc2QASfvwgbzsyQaAO7gnJNibHeE1j+MV88MfgWOGhjoIR7atOMIgaXa48W9eayJywSG4uKCLEx
vm3O9TAEOakElk3pGVZUyVIsAPxYXZdcE+mYJv1eueq7WrlRbsi3FhsIJGY8EvMRtg5+NMz8VQyw
0/DqOxOWwgMvczVdzA8JHS6Vy/4GXq+gLIj/jAXteNjTcB7CIQN2GPCYRiryWt+1TFDDpw5mLsnE
y3/JF1TWioSXrcW+yZeK1pFkZhNj4mLOCMOBhEwAklVTbrn1em3s6t509Ozd5OiExZolwdPnpbKA
XmFNtUsBMntphYF0f+HatEPqaH/kcJ6RV7ye0Qd7CaY8ppepKgX/Q5o72wKoGWLhI/jVY7Cuqstk
xalHNzIpqaKkraL3OlbFRIHOUsMqq+4oLr+hqKtSPEBYX58ryDsnIxxm4h/AkfBnAzVj9NE7/ZKT
Sbf3Su6tRA8pWu3wpIm0YlaVMMfnVIrd35Euu7t6hc1H6njXIFN4QTtlFG2BUoyk5AiKBtVFv407
44qao2IATs6GWGpEyFkRpSp0tbp3FbbMzBM9LQdqEhN4nbydI3cb5P11FfGrf7B/UswKWfOOYdsL
AL8OqeTcWu4tSvBPMHWa5NCS90MvBSyYqXpDlXsKl/mCrVeUV2NAksUsff5kuuwBJVcIwKpIlgd4
lZPQYG9/yh/fQaOo2FWbwXERt+7sAbzU1n9/PKJxaDpm9kXFE4ZJgEIn6XFnAUHvjMFlG/gH6EGe
AlsvfKyX4Sc+9oUK0Q5DWG/0E6Fiv9j3G0fAqkGwpWPDvwuywmEHkxHLG/k6SX3TqsRcs054nGyu
AfmFzrG3VX6mYjFgQ+ybcrhtJOvf9Nd7yUMdqHjWgwkyqSGEdlQO7OeBn/FtxkwLDvnLjlw5dAPV
NvHC0dcQc0Ep2V7yzvQyWAx5/BP/va9/6cUOFtvViG/r35e61adcAUPObLT3f7EFSuKld7Re4NYb
pmMQlNG7QACmrF33b/tiLXOaAMZ6AFsXJMFvxJR71SiQXOcL2dDoIKfltpxwjERm/fIEvOxOX9/4
pdNhqKoA1lMHSCgmXT3ZtpgSUvExuLf5hBhPTA8b6wM5u065aqab8dso3rqeKDTCrIIfrVxnfuq/
GRwKzAIAewQGAzr9f2f/ABkwAXXCRJIEjLBwKGsbad3HPWqxoaWl0nuYPB01lDZ0BNN2lRN8jIPF
3Ro5G8S/8yqEhStcpHhKLLP531C1ML13FT8MpeDtxntK2xdORZPPKfcpTDBow+okS+ZSvQsRmZMn
iaozsMy14Pzz3QRSa/pwKpPHZKxpXoycZFSzhPRi95+731wrikh/8KBkPr7omYCIr72PHlBJ4fku
/uP0uD4twGXz/NbtJvN1aiJhieUBGpL5pi0G8z/UIB8AcOdNWvnz1QAmG2VYoHbIXnS3yXmiLEEA
9UTeUv+J9KyoHeHHPUjNZ1IxBxzMZAhKrjNh+l46zDtJ92y0S4BY9J0tEGJVKecbrcuQkNyiViD+
ty12rEMijBocWJrWwlc2GaPJgB1QtbfnOcQeGAJqRvku+OULPfugFFxNJYJRbrjMxn3QxT97qq0V
tUBShqDQ26xuhmVqqBMHkblibaZ9t82h+IvVqZaIWM3Yy4ORDQL4SFISjJG7+WJnGrrvRDtEebb1
pI1qR6GYZpG5DxgGr2dfBaakuBphVdqN9/9sv5BC9L33J6NWGhWRWmEqaLamL95VurWx70bTM5lz
o4gHcDz8cS0/856au9Dfsxncy11fxYgUbWswTVScW6lKsR/YAavBWe3blg6LolgxAvWcCBbFyY97
ADILkWDHaMpolZvXknz2n6qnHLeR3qmEadZgV2pj7DwlCf4Bieivk3qB0fnX+LgH6N//HQlTFs+J
TuiNmTXghzqw0bfLE8OohNyUnDr4/mbkjS4i5S5qKQwgkIa8P5N5upDE+ZqOLT56S8hxp4TECyQ4
RND/F+1eBebBpDK5JX8fLDEkfeeoEGSVWA1sTXsK5E1WpkRK/XilVXRXVGR7JElfBgUiIYRxzUkP
oRZ7/wQlQmqhEcDepiXH3QyrHY8SXOdX5YWgImc+Gz2o5Psp5N0nGytnoXsTPmUvL8LcXcs/ZYcN
IjwglGp9/0CjnQFzfMXbsDIjzhuZUkZJypw1cJN/ZhjMEyo1hSb9bi142uWvxHiJ/26Mh4yKp86E
k1AQCksooOh5ytrOwyrDC9rebySu7jkMef9VyJkNBGg4MVw2rmkFeflPjJSp9SXT+/JlUXhzypsn
ub6sFJLyUFJDijcAeH7QgGxdEnLrBDxnG4vAiE0ICGFasBjxXZHQDt9wNHNhKr43wfQsI5qUHKw9
o5NOvGateMK2HAC4qM0bnY66/KwNO4dHvZNcH5PMpTTQ1b48cBVSqQPgJI+sd7ONsLUNtCpzVNuV
vbHnQL5iqkvejXHJedwn66sQw1wJNhSOqQA9UdoGNhokfkuPuBJgppICR1i6epKY3V0g78BR2/I1
y43NkJlAbwfsAU5xI+9qNYhCoS5h6wRFBINHvIi9oE7uiNj51YB7wfFTKYMgHBNriZsoI3t0e4BI
c9GYCM61CHPNvvUgIjdssG0f0aH0rulnKvsAkmxUCfPqBu1qy2aIxxopDwJ5BR/CWX/vYWW5bKId
zS8W43LrHPbe9+sFh4CB72G07IVLOnV2U1JU3EYLi6KvZdA4igVOtgUpR0jKjat1vHoQiJS0b+R2
EcNoupe22zwxJJJ2nQcej5CzMoPNntsBGanVj8My6UadBR3aOFOEkuuKlsgG4c/btUpl7i4u9lll
NI1GoHI74Jer9WN0ejyPBasL18gEE2/Aeg0wY2ASFNxSJj8bGxrOYo9cmYnkt8kr9FZ0UrhbTIsW
VyQn0MmZLZrkaGCLRQdG137V6oLltI35R2yNPH+yd7cXXNlbb8imHbV3MGg7p5OqnLnKBF/n3Qo2
FR1JnRlAmWoz7cMUJydzHCU9EPLzNtfJW34RQifg1GetFpySadvENM9rgRXBKbSWmPHI6Ra+YJxz
9dBvwWS5UAfF5IGvAJUJUKSn507wFJPunNN/0XmSh/bze1Yj0z2vkXmV+hY/eGyFg1qmC6Itv8LW
bjNJMfGTvWhwumPp7IwpRxFhIqMi9gd8JUfHaOO0R+ULNpuxScrDtzXkMVhfh69xXeV0ZfokCOI7
tMwz8oDiVgu7Gw3wBVajAs/UF+Ou2iRCavMxzDh6ChnEKmGp7wZB1hFYMoytTPaMOvqE7g6tWwrb
O/A/nKN1gsNSili0ZteWW+yRv1U7LbIRK+r01vZnc8xdWNBx9xjB8EPCAr27jK9HdEZgyAR57A7u
GePPpG2q6zf1359w4UOFQLqWa5K0T30dTYn7gl4ACcZ8a5/Yjwq9IcF4C6i4w2graZRoTCMlip+g
ytAOJPVWvIUtonKr/ybchIJp+OZBp2A2MT0CwmarOUYaEByYpfwOYvqzcENlrMgKgRJ8E04jOel+
7YUSfsP4KoCnEDhrkVq8JPnlgWBAxKDggbgn0XbsewxambgMMJKckM/Zco64y7Agiu9M5vYmQJHp
61AODLTVuVC/VdM06PnOpw0P9ZLPNHj2+OLSi48Rf1JSo4DYXmls/xpPRDMH2/3Hq7+rPZ/SICd6
L603AMJD3c1ekF7TJeygqOuV1GW3+Nnz4Xdq1q12tZmMCxvPYEGspj6S1WO3BqmZG64ZO+zb2BTv
FQYJxqEd6uZ1jU/UEgX0ERZviSNUIh+Lytn6c4pm4gBSIYP4RQ+sv4RmOv+lmrf4G4VM2LWEo811
STnzIy4o0vX+n3uH1Br0Z7BPc8woZNQatJGC4LncMEXtX7qMG4rXPSRHXX6R7CZ8cc3Y99I9uNXF
IjSxjDVJz8Qktav2qlENMkAQUW2CCs+SRFIbb+hmh/+8/m8QuO94uT2pz2tEw9k2G0HqHYZyHP32
a5d/asfS6+21peMD0JDwBtdbAKgtjF57peUTGQgIXMKrX8V1BbwDgKhfLYsJYVV7YWo2ChFOHmvM
w45/28ZFISF6kHIyW6ExajpEoNepQhYJRu53iLDrMfDu02ajSbpi/llU/v5ug9KWpRD2qTLHNt4B
1GtRoehlEKVT9qjYG4/p0Krw/ctZLC+G9f8kkzBSd3EnfRqrYeglfpSDEeMbn8oqc74IkMZA/JpN
oI1iPxqBuohS1sNbDwuQsRlQJxHYxuc41iFJCHLnJvHXNRWo55wz39q7yvCB3105+TocHpb7VztX
sRallT5EdurZ6amvSjE9TGwiepWk9SgKA4uo15u9hWjSH+HWhI3YMfzKrHItS9N9Zd4TtcWUmKYL
SC6Rltkb8aBnT+te3i7I2NR/WQgEv5SvNlpZwrMNb2MZDWTcgABmFdE0xHExtxLy+xIeOjsCVjUt
yFnMYIRpqzoF6lXd0msKAYxq+TvnVKm8Esg8rntNOx5y11HN7KQpzE0TAj0IulEKkE3z7B/MD1jC
wG3m8BZsj5acDqLq+HXDqtLwwX7/yHmKYb2txqrBxeY0V9Sk8fFpSErUXmoNRgSDelXxAWnDpCDS
7CBluB+6zYmX/Cf26wJsOUDHE1N1Rb0PQ1FX9zledfLagUjl4DDdF5G5CNklbW8o55mFUcZ5UvfB
VJXk11LAeqwHWrTknJL+kiqQ6wWmQgKv0Qj5kbHqjaSFk/Ux+QmRNgezFbVR+TYTl0+XeBInK4Sh
V0U5sqECWpVcXtBW692PWaau1ujZ0EPnCwDwZeBpTi3oUXBsR1B2LFSdlaPm49vNqu+Nh2jJ28Rb
3Cl62AT8waxsaiIOP2W6dFee+S/4OuTAQwv4JhrbB7E1nNW2B82whu0gGGNFvddOxzO4oJ5SIjmR
XEjXlD3Pw29psQklXLnU8nNue6ZK8j8I0+IaEGSAVjeubbJM9tU43xnJy9sCIU781iay5x44WtFo
LUUFCHKf42+tMCeZNv8uuBNl+LADjeGD6pYwjcs6X68qMIxdxwZFsfJKOCkf+V8zrABkV6tEBUsn
yt8NrdhdrBqK+yXkXcxocuEj5d5wcYp4yq0m4fS64K1gaUKh5sXhncbsl59WN67tpFAxQo547Vvl
ezLLYdUJDxc4q1UFcrzafffd8k3297rhp1WZEFbN+Ou8jfMRmFr18EzhQxKqoWGmNd7LJtnlZ3Cb
kF6Mfs6wC41MN8n0zlGYpoksKzntmpjluPSiMcYaYNaIz6MVHNEf6rQavvBROkgbAuHTy/9UAKoM
C3oYgmjOQKD7V2vX0lfD/e34YnH3cgu9k9NVoEqJ3mKbBQn/gyAyA634nh8QYnqW8hWGd0lAQODO
/8uCYoGRHOjpySXp7KONibs1qwYmcx4+a3hUytfzqYaSS3+G9eKF6N+pVInITjkMzG5wxMVbpKBv
5WiCAsnQBCa1l1eBErahaQLHQGk5Jd7ekTdZ+Ozxsw0rTIJTTG1uBnWwrksNkZA4fn+OFe8GdHDd
CX6IqnnuZSz56OTdj5r3OJZ94bK3yj73QBG5E4ZKbYZleVse9Kk9CyA5OCLMb9PSfvdhGI1nYSpe
wnMp+9lYvtcCEkETMJzBqzALkTEcRxxZHDNyH6jXwHnjMEmvKQbmeRzsJ8h4VkE0pvHFD379geNT
yB9rJ9GDlM3NPek7Cn8ByTZI7mC0sivczN4ISfoykuqWUNT0zX3Ket/kwH/zmVDp8z7XNwgC/uDT
712KVS2TdF76nYbEhSjne9zOKzH1uo3gywHtffXZliAmMZFbbVxVqVa6TBYM2DRa+ywGn4y9teSk
xFc8va8lAW9V4pv0lEN0X8B7H1EWNCXUiUMegcQZuBHYy+W0pTAfW6cHlFWadKMwWUdze7FAsJQB
/auwYdlHXGxhZBXmDH8UWVdfakbjd72rVavbUqCIauh1/woejHyZJ+6QdR+9b9nTXgzuCVxgqg94
SSBM/fLSb2e0k4PUZZwpNtAN4WU6vRTPPejw7c1Q3lImaK37iIxH/q02XmLYfw/qWbDMrLUJ1AnP
qv79a0u7he0iRIwKNzmiUvBmKLh7i4iJpkel0y52s5E46XqIzDpR4aIpmbjLLCf83fYj6rjUmbyL
hBtJcM2/B2CZejAuLPKMtDWnVoe7wYiwZjNhHCA2HPKZGiaaCBHqNkUs2o7y3XzaE4WQE2iOnxVf
NtL4pWLwt3IjoUxnmGiLusaZkbNC7dqBxnQNNS9hxLxk6nd1SIaq9gdP3fBS6+4qhBlBP5s1qZde
HEGsWq4Bnic6ry9/xprJoFcACU10cZtxtMgl3GZdinti8qf1VrHJ1AamgoMtI/IXFB92kxLtzKU1
GOQnYqLfFiIRU18IP8KzGrhAlrZcce8U0+zwa1l0HeH7p1/Hafuxp42qiqiex15P6/qLLfO0wNdH
tgjLU+uQa1nnrAnTUsYzmciuwCKNdqygErSl0CuWv+q44Rox8RUfv0mrPdc1bKGk7ti0/C40+Jmh
jgMSw0+t2Z1CelO29mPdoP/VHn0vNy3/tALUf3kMjQDF88bHdFO5xy7JsUQ2TCno3apNYrivHP8y
zZw4R6OjiG4+7ONQbWjH+j6uQ/ksx6w2WnGSsBXcKRoqz0JiTRAZuUPpiMopw8GgEW9vfg74gWhj
uvi7ythNuQZwGVb9WfRhdMzXgdX7Z61BQYq1+iqS0ibeC83NiFDMxlgTUZ623BuUE1aq9pcLgm0F
+4pdfUPo2nH5CjUDn191PjpCkwu3B6b2DsyUx0jsPPkAvjlYv0RQS+4UP5M3g/6/4fmLaFpeIp94
L7VHuSG0ceLxzaIEsP2K9S9zJExVGlDqEXUL2tVG1Ef135YH2HylgWRBMD/dDtjgw8Q0z51kJp3E
hACmIog/Ct2wzha7YpjQTAXcpnIBRu5L7uBQzyKi75l7/m/bcqRnEddK+NDMdBFpHKuZwTW5PesQ
MwG/O/NGYJ2EEavy12WqeOQ7Pb+XQlSN+yQck48wPHvyICUtAZ/609PtdejyUpSALVtlIm9b2Q25
MmQeEhbqfMcpoU+FAwZDuRIM9CBzlb+oZ/L+xR9Jmoly+yizLlLJ0LxJtSszwS25jwlTe2ZzTexT
DYYxBRIFv3Q1+xt4ZKPTx4SN1H3ahqZ9hjSx2aDqWKxzg5v8L19tv8eNpuwtblFFK8bQ2ZTaDhCZ
TSZNa4rFgq+sYihcmrnr5CmFFUMAol5HtQIzGKUGtcS9YmigzQ2S/9VDllGAXsBbtAvch9jobrXx
AZlQEGPI3iPfeBOLPqhhpcA5eQFL3yZYk9PsVJG2a3jDo+CNG5LLuO6WeNpavTtO0bqvzLCvOmnh
8MVdj+kVUtTRZmOngNpqvly1nJpUWZ8z2vytvEts9VemRx5wwlpGwVSJTJOdLLoo1nWMUfp678Le
FANikgvXg2V2t8JsDvjZpBCaYCDoU2LkZovDOuK1Rbg6T2uCefsktNMCFSm2vqwD3KRSH8xGK2f1
wVF5brcQe/Yjntuep7LxbAmaiafQl3DcbAcN10WlChGwUGt0dTX/N9MfHY5pqhV6cTnjf8PGp4Fw
nzB4gfy1AI6qntFLaRndPPOh8YekwM8dsLW0ehwhr37vwGg6eju0CHu593AdM/gUJ9u8TmLzzox2
27sTsn/uCBMCADhEx5oJiww/qQoelHD6f1sz/XIXDbygB4oTV/qgQgscZP7/D0+laLJcYlcr3mNY
1Hy98MZKVvB7180iAueIenHdE2KCJI9nUo8FEUZCTqtngPgBUm7pFd3gW6x8AdktPmrMgyZgoLuW
mDxyV1/70LJy7OUVap7qqHOBHhz5ShvB2XQmaPbtyKKw7yTY3aNpX9uDlFXWGcnciHh5gUhPP3cI
zMPB3ehrwK2n4/XBDi5tpQRz7h+QyPJbN8Q+hd4PKufKdimpZAfwLGcW2Xqq26Kc9ygwi0gcVytv
X6KugI0N4PBFEcIPSiy8ayd8r0xjpL3Iu9KHs4b4OwE6MkjJpagxQ3WGod3rD/Q+DYyN0xGuMecF
PRutEh+wYBqZsYO1+mgddgsSFcNhTVhDeY4vDmUXmTD+7opwoYHsddv/l4sqX4RQylWL7Wc5e+QR
jBMoprKLgdCYqOUTAZYeWTrp3fvI67Cf4JICoQcL69TYyiYP/o9VhpYpzZJLDYIi7W+zAXGBGDbO
iXSdvdgAHizKn3bjzSxiDhKmrCYyq8XXL5T70Px1fnvQGHmejFKSL2ia9xkv7AK+EGOcDQRFG0QJ
jb4tn11fk7pbTTWR/x8qg4U+bdr6CwcGnsE1YltlCQuqG1m73eD6/AcYw3sPv8qvzbRiqCpFZepu
5EZqjPxeI6yQLEEBBMSL0pzSc151iTXR0Zj1QTPFNQbJwn4dsz/hDoKqzWdswWRGJmWdQLUOa6SW
9ZQ9O1ovDcdGba3JpLtPSXS4x32RBagGP/NBtxTrLOE6jRfFnUihrcUSQ1Afrd+VqhFYJJm1wmqs
K+9lFNh1R01qbFz1+YBBhzxebMqB1XIHC6Q1oBOo8P+N0OWHwUiKbSAxoHIkxz5bCyzVXzE3c1Dj
z/ZjaDkOHWWP4vwEyeqsJv1GpTrPhTwrSWK8XyZ/zGg/dZ9SPgnSUb1DOd+uPmoH9p7a5pGRPh/z
g2kOUrWus4lHapREgTOGzpNs0Nb+B1HW7+fVQLDr5d7Vn/eON+oGg2fD+UcgpgAHFoqBBG0EtZPW
ngYVH0mlM/31AghG/ZnQMxnNXNBjF8fVOx61++ajkRLWBqDmPegU6jVjajNR/GQIfv1CKt2Q1e4G
OXB7RuIKakjlqecCzG6zq7TWgF2X+hxpE0tKc4GexeDyDx9kcUJByrqOPMYNLCKLKS/42BNMEsHz
AxmZ1FaTrzWMaQ7kXN9xRlayzWA0nNionBNiB2YJCNvY4wvYyaPFEIADMtsJV6zKZCfbR2GJrPvi
vvE32CXYC8qHE3BKEJOYPX+4O+BL+vdNv2+cpcdwpW5MxhZN0Uv8I+3UzZbMV/m4zrmJ+DDYWc4A
SAeCPDjrW9k+nvXwmHOucSW6oraSE6BDH/f2Lzr78w1LuHNIHTuAm4+X1Eep8WZ+E94uOmxdZoBu
e3z/jTWr3Hpk9S9yXBaDhnlhg/nbs6EKtjikUQZ1dRQWsJvdhI9VWfd317udU979/WdgnXJYBQxo
xwWIa7HpPKHjBpwBpSMV04aMfNOS5YELWuNli1EIwEMlz54YW9zasPLFCn5tm8PoDC5smuEFpyXy
RO8CuaUgibnCjH3v9DgfXlthL2bzUUdv1Y2OZFJWcU48LlUXfmkxDkZjuRYAVMRVAHthX1zUk3QQ
FoVJMg+y0w3B0ctLojMjIPzmHjUNWgZAqlzy0IXVL8kH1wkXdFPahjC2g8mZBGnzca7YLURiaL/s
DMT2Qx8+RzOcs3a8Z6U3z8qfXAaGLPWpWwden7hqYsqF/SdDJ+IKZF4MNMGj9/Z0dh4qiq6cb8SF
wOImQBI2ra+WFr8p9uxaORtUWpXjlEqNt8rdvFuBsH3u9VlBMn/BKe7kWt5yqbYfMBYO2ODKLMnR
/4Vzl5K8CapcK2ajgkEf9ZpsV3Thc+QomVNNu6dmm6e7jL/NybKsKr1h+USNqfbe0Du45ueyShs1
+YlpASM0BNMidqjmuJb1VvCgJz6MwD2QQJFHwEGNY9qkIL6UpmqErzHJL7ZmBaIcKIQwRFeQ1/rv
LQSon5Nl+SwOwqcbuyBc9CCkOUGkN/gmMzhU8q5DValJ2jvSG/7WflnbULFCp7yaCJjeNI9rjUb9
AUSkwuUrf00lrHXeB8hpvzHlmJ4nJQs5qnZGVVQtVXGDb5p7lTaPns+uItfCzRIHvVpy8cIFnydr
81LUok4AQDuvqgrx8QbzHQL7qZn8d1HngvulPZZMDOGDDRHmKqmnKm3YzVwuUS7PU2lJIrHVbVTz
7BI6VEyuM4zA2AZeYZIAOW1ZiW+WhnGkxCw7rK/rya28x44qI9lYRzZZjFQ1ECEZIRBDbRNltj11
8yTFMMCJU5ncWsdDlLSheCDTayw+g2KmYqiPkMsfWrq9sfq1tQTSBvK4FsvZOtLsEkshEwMxyfu2
KzwERFUzQjPgRG1OuXJ60Z6VSvcVO0uQT5kMXD6qYHcu4k0PrrLGZFYeVfqJdkNvnqsC20FtOm/t
LANa3yEIhDDyQ3cs7Z8a1BiDF0Dd5zzO7sNici1oYmBL1hu6QEYEF6Ju7phLlMYbF42d7G6JyUae
ePZZ79XEpmQXtGpHNAjBkH9mJM3R+YfQ/EfLmGAX6PItDTbaJl7riKadAgbE8XP+5E7QH0oQm6eb
GUm101fo8uDCTVUNUXWuGI3k+XH8RsFTv/8DCm2kp87enLtFLnb3uOdjCeZnuEpdHATvj7jzJRHM
KUM9jFhxd/heH9r9mUHNCuVNeW4V4Q5DNQtlKsy8U0EO2hlEe78WLclEXMaNJkPE+6ijpM812aQc
HcUklbrBI3gbUtCI/835g7GWCYI99RRrGxXkodrOWAK30/lw79KMU968yWQCSICGwMNd6sLwdGNV
EtYAhEOlQagNwicLzq5BDjZJt8UGO0s59zq0jSRUTIneO9jQHSc8oYUeAQ/6mh2q+GenC3GXyq2a
bkVi99gMHP92pg+77wSAsV/qwYKSf69TaNlwIfF2sfHIOFB7yTErHRvmXXZALFgfHjc91SODL+Ht
7Zt2jGHfEJsSYN2xO3q82QYtYJKCeYFp2qD+ZRtYCU/LyVTEWqyWqgJojs7WVXqG3ciRBzj2Mvh+
Bt09NEtSYzKH+ygm+7WnQm7Q85tFLa7hy+ZsyJ9jx8qY0CfHvCyuaH2WUbudwIq7NfHUxuReKHT6
WdO3mtCOUZjJu86PbQGqtI0jlOxPFVQ8m5SghC2qa4Yv9LmOsOktiLc+h8AtXYskF8UTPtUnDkIU
mRB6tJp7G625CpD2FX9qmbdpcLF6wOHyYLvyu57dtLpD7jnbvQfq3DrywSv3Xt1BssfaM6hGgQq6
N4j71tna9gFNjVH00BTevqdsJEEcLK9AV3Vb/5+8uipo0u/QbRVvozkZLQcsrXgIEBgPzlMA9PwZ
0s9mWbwAgOSbdcbzgG5qjRhfCLdyTcD5GL0LtwPIuNnIMKRDDchG96/Cvbp+D/c72WA8m3j12Du+
guqXSD7cAjg3gCWGqO0X39DLWWz5pYZIcJx3tvWU6bn69No2Te5kd7VssE62eFVyGuLVYShxOt8K
xFzzcTaEw399fP/d7iNHU6ZLfkEzjxoONYO/3hUeG8p2FduUug2bMA4TYVVt5II930cEVptFNf5C
RSiuSWAmIPLB4KRZeODbLyPC7OSWZ+7Phqitvz8N2xT2HsesaYyeQU+nW/q58wFxnfdAWMcXNVKT
Gj9N0elnVIDDR+fAUB2QD0KHfMWR89Rsrch+0RZXCZep4xWI9U4LvZsd+LAUcmjAwCKybMsNwdVG
OIjQ7rddlH6IoOO3BlhUd9S0BHYonckKipCLW2gGmbpt1juVB/58F3ZqrzfOsOXq4LRoN68Ggpd6
m7FXdXNLFodnP/Usv/yGceTG9suHJmpp0EwjOTlZv0Fallm1++HFe2XJ4nYtp073otsynRxsfBLA
j7wCX2QnuIiPWcexR83NkAkxxl1YPyb9N7B4Lpc9lx2VurB9tJpYppwURwxs276avuiJ7yM2KCDj
S0g5fQYSm92YlXmkWBCDQeM4Pst37gJgS7FOcDwVTVqKMSYK/0+VlOrHEecp26ucIkZWKxZdTvGM
NLsLA1n77Q9CIti+mexLHigTJvRFORz+gGbeoCRWg+pJkf0wpGgjatGYmqSHNmp586DAh+5I1ln5
JcD6f2zVJEfplEqbTuRfb6P4Epli6RcVULCFy2Ugzl2BIeBILV9uX/frlETDE41CnCtwwk5SFpav
YMCSFwOy2ATPG7DHEwn/yZ5GXmSh8t+nvFdRA9Rn12hYeeT0mTnkwcTLiTP2FgPcqYF0yuEbfOC6
yU6SLGitpuTNWr/yjjLljsfh47d7o6QcHhDu/BWGGF2oCIj25BIkpBKm296JtD+OXSyRwkGftp9g
Xo0RWaRZr400miGqCMDMh2ZNtEmsHwHMkvByXGRpM2/wF/WtoDvZYcAAhNro6wM10iWrcPGKZc+g
Co2KURQBr3qqMYfsPs+OrvLX12XiAt8I3H4K85Yghfwgi8Q0o6IYAPYpxthofKZ/Hwh6gagxRG0M
4CNumbgVLn9C6N7KzND9Ja+M/Gt/oN+E1A+jLnLS2TA3GWIjn0QRv+cOtc0q5pLIrZqivTcHqN6O
x/1vmEPYr04hfXgsZwqbnEVB8Oa6W7v3sHDfexxb60KdoNIgGaYQm8LqnX2es7EKuTa40j71KyTq
d/JQuGWgln5hXIbhQDsQEKCzgd7cPQNDQYzYF57XQC0RNJpvq8OCHG4daeTNhocaK1sxLoZm4YN1
SExvRGWSjdbmzkD+ToVxfD1x+7fZqRj5wx7xG30DpDiQ4W5niLhNy3xIVOOg1EaKhOmul3Xx2jco
uu+b24pXZxEhpLRa4qRxntgHZn9VPasF0d1rWJgq1JtcBWWkGg+P0rIERLKX4aFa1PfyaViP5Fm0
jyQlohxHW+B0r1QD2Ecyy/PLcsaxZN0b8ykl3tTranL3ngU7yGYHU7j1N4cVV4psEgply6b+5Jnj
sWEo+oY4zpeF0cpxdvIfhJ6rxn5wIS96+b58Y+BsPwNatbDwk2f2PjD/JnLChqSIr5B2HXHHah3R
aPggP2OJlOKykaJHrhtYU5HYpOVmbkTEaxd8wuI7uyAMzuilhF4qAjHoNKXk9EfLvG3ma8EsHtbN
MuY67FkuP9RoNZZPha4QtanNWpCNpdKSw2Ie48jxwh9LqADnNDRUPa1LcA+0JFdogPNV8cczb+Bu
fqe24NI/tz9GqODF2NHw1szkqtS2GBFZfhjrnLz3wyAT/ImMLym/vzIrRQ/71IsscVZseL2Su2le
dGawvX5ptD/S2qcrob+adklM12IFpX36XaRoCbhNgRKkgQpHY5IJiXE4L6kfhAz+J3hC08pmUuAz
7i+4WJ8jaAXe74wf9840Tu/BzUG6v8e8BkCAndk2YNQKu1c+9NFg4qt4oa93fnSU3WWLd5x2dz+I
nL07lOOK0IF76m34Wvzp4AU5JYvy1sndly8JGJNbhLNvRFcQRCai26MZKG8rUp7XeXFHryAhy20+
Vhjw8Vmn4JftGygUh0NiJ2n89w/6nrh66p/ch1yonf9f8LoXc4t5k/5ZZgPltKX2fRF4FgE4hKaS
3zThtXeU6bJdgddcyf7BtuwSL+Bc8jpSCpAZ2aUkriFwXCDIbka2V58C8A4X0/uPpuQgElh6Mxks
zB1iAUOv77tOr6GH9xbdlRxXkbKjy+I7H0JbuVLYj9Vyacmve7kTXpphQ9BjRCXW+PZ0oqynPAFw
T903+6jT7vCyCmY3dzZX4RYPTQrIOCG7zLQK91AGREOhJqvTh1/f2D5LCa+JVG7TiVqsdZHmcS/G
JA29V6avgNQSiuBNPnWNcq4jtFhz3KckoXJRQNsZwtGrqNw6HI8o0G0uBCgpYfmjYvitKwQuxQvq
5FIu9bOXgmQOXIuQ/mVGoc5mAySVwFei/MG+TknSE9UJZcIkhLg8dB1SZp/bfedaP3cB7td943u/
Bq3It2G92SaT4wheQP6N+CfSg+7ALKlVi9UnUhCbEctr61Ss7rtqA1hwYEW7HZ+eW5O02HDk5ydN
HoWdTfpOkuwPeivS/q/0YHPH5cBmJZEQ6rP8QsDfcWCMKf7fTI2GPjEmTFnOK0By/AEokVnVf+4W
boScTcmBsY1NfwWHm3sC0+aFoPJhZ2s7JEToUSRJYQo/JtLZz3/BGchTK4+hDWRVeDOH3AzpHrIF
XP/KmmQrlPdybL+sbHTjbFn1sddPg4CbsMyNPifsFzlbP/dQkzUo3Xw1R+WyYGFDhwmcbOUkJ/KW
9n45Z0qXd7z5FqHJEBPyNmxaHzPESBgRMf3WwlO9xHtjvEOSSToTFfWalmI3YN7mk6qRK+8C6MNw
CvSUzzmXcEhYOQGiJ8O8dI9W0EtkSDP+FjvVaw471GQreeQ7zROHh4nFV3j2InHmJ7Z1BOcFgzCm
baKlyzL1Vh3518BYwgd77Uy3RY8ByCOvl1N0mhHiJ9vkgT5ZZ0EDr5qZnYaqULI/ef8tXdqAN/NU
J2PfbUU9v6y+VPDao3UMJZxmf5hOsXSHq5S935IS63qB/uweJVfEupbPkh9fVrH0Xc9QexLJlKub
0Aw/kpsi9lwSKD5QxUND28U7dh1DosbJRZEWtwTcLZrNPiQVnSOUdTwExsg1GcFLHTNM3af8JOuf
jQiesesyK+ImixzULdUwMAYgeA2pHuRizzNj9YYQ3iMmdV0l6sgjeAMSc4N4jUDSvvWkulvhPUe7
gH4er2o+60apKfwkcMCI2x8AEp2Ybu850EjHTgr9WWCAs+m8SCl/yhio1How+lNyXkckHzOSdmqJ
mJ21WvmeyNI8T4aXjCaEcYxwJXYR/uTCZjUw37q0vvgWVSYj9lUQzMluv0F2cNZsJ7T1TEudm8FT
oxUQg0JRcNMyxE6y1unpeucZ39rM1aoF+x3tw/+QmpRKzwpDW8uxTMj4rvhEKr19XN0MkYLdd607
KeppJsaM4KEaHcJq0kQfn6nV5eFyPW5kUNS6ZbHJ6C49qTpmIVFpRjtVaB69WXosvbC2M1eocd/M
JSOD6U2L3sRRdTrkzhOuDSiUsYX5F64xGutMJ55hnuAI0zQxnrpOEgcs2n1UJ2/kz4LVSTpNKRKF
BfIOUrdj1dsBI9gLGdqY7g5diMyowv+0nSm+zDGLF4xFpxlTtPsfzv4BZKl+0VSs0bYGUL29bSCq
fkMsY+3qrhl/npQRzSYHhbdVGvbY0n5o97PDdrZJr9RL8QtvLe9aWg5e6ts0BSIG6oCedeGT7DEY
GG6H3UM4RRymQr1cUB9DHXAbHhpetJ6PzAL2/tRLYQMn8fv9xqBQXhxNRgFKjGKLoNet0hZwsAFC
ldFqQnCO9qouejvoi5lpHeNk6UtkdJF749rDC6gmwZqHLp1i28PUbjwkmFQPkYif/ahwxSD7MbEi
1NXHWw/wenerVUJW0W0iBumUUygLVLRHHt1wshQZA6TNJkVjkepUobMArMFYTSnTD2Xi9Ljz0VyS
81Lvk4wV6/myLZ8QF2ujnFmE0XAkjYaDROd+vo3SeYzVs+W1+C8hFEeVr/Us2h8EltbbThXpnaPz
YI7SK0bUR/ar50j4j/6JqpKwgG8yGyZyWTwJNejWDkf2ASQusTjuUuqXVuzQD4yrfdWbb8FW+z+M
xksNpKMFNUMPTechRqFqmT/SH6p+7xiunlbS3QJlwhI1cMFewS0XujEC8jr1j+BamIZnQkcrpY9Y
yO0h/MXu+V+5s8QvZlxLNvs+xOXHG6E4HEe0Q1wagdxNaIHPdYfd1FPat/x37PpGVSeC9nRn/GVd
/eII+C9qQGzO+INAP8DoOEndfX6i/dAO7l6K3ZCDBtOh3C1tGrrbdo215w2sOgl4pE5iYs37UHfW
KKLC/x7FuwNC9JKoSroKbozALLtEr2MC1LYH1y3Go1qGxTbaFnWhshUg77IFhryqdc2oyBe6JX0b
qf68fHIGVtXclJhIEr3bzmFgbdy1fbBw+5lGMHu54V3w38hVrFtcXpi6JybYSTN6KsA6JFgD6IVf
8vLVgWGmWzjKlZoTBDNOaMZY+6QqSQOO8eYORefXqjVxL6ZwSa3Exsu1K1dJYlPBr8Vwr0GYXSZw
iRM8KJMEz+PNWhzSraNFHdnOLoTFE/q5ftiJ3G0lOQ5DBnvtdHEKYHB9rig/L9PV+g1ZABR6oIKN
NTLvfmHmi929qkVyiSLWiz49wOwCH89gKVac0oNwGV7RjLZ7s/FhtaVTprfruYVMIrYlHpveEPQ6
xhgEJ11LLjWzt7GrpS8zF3gQX+9SSZs/ZpgGJYzpyJrjU8jp5jnsrsqy7Ft/moHCM9gaEducY1C2
QC8M/B3GHwIXghlpfNZHyWSjYvfbVEmqBOpvdvcUjvoeBdMR8U3GAkSAQk+NGEYEF4Z5aE8Y6JM3
PAKWPFz/8s+jb53AWejy40ggd6lxhcbqocpQzxkaTARSxXQgim6qkWSS5AnPvspB6FBhDOLiNwOD
l4o1XBRKMTs9Wm1HHnpAYg7a6Kaz8s5GiDkkc0NiHD7yuzMNJLUVQYhH8iWAafJdZE4TdSngUDoq
y/5z3GpkVoCQVmFqXuR17RGDtpMqJQ64hm081SMLoZhGNmCw/JY2ZfM16TjinOju433nhjQUidpO
yk7T5kfcwRp9AgZMxtJtIUeIdpoqcY5lgoMcx2jk3KOFwKcaLwBQWkHtLLRjlCdk5Pc32BTHjZgR
C/JDmud/Jq0M6ZiwgrweL+foR42lohvVGYsjovKbxPyg7IuGKZsFpsy+luTpCwdz6zHpdIQiw3AQ
UoeOESoezzXKz/qdgDRrkVOb8f+lL1q9cMD1MLBKG1BwRgzFgIHhkBuzQxKpm7Rlkrrx+OTNl2Ay
2oriGgQyxOQyrrW7lqKq9zlC+7zupZiT15VxRCgUuGI32PvaNNqwzt4a4IH+zXExkdS4x/6xv8VT
2ruSK3IZkzTry31Y+bTpdl5A8ZbxqWwvYl3pXPkLe2ooq7FEL72X66HXkTsBihJXbWfkasoy/+K6
w9enjrm6bMSUIIxiioTgdio4G30Vhj9ILMv5A3hjpv6xHcJyBnB48F5SzMYe1l9Er8EdEvtyCPoV
w+6EI61LJi6nU33p6OWUgvb6gjgjzYL4njqIgAVTlKT9iaUKM7+Wq5OViY8M3KEIILZZHTGShbzd
QecLCxNIPBd6yjWq/yCvaaoSGUCyFR0VN/f6IvI4Ua5WkLekNCKBtP3Ss8FiD7L8QjXB8OLs57un
1/rwP8Kv5v6aFyVX9pyWI4hJ6NOjo8A8jw82D6vj+gNRFyjuNuKeTgr2xjPkDnpnsvZ8WtBArsWr
aNRnxpt4CVESzkLauaLIhgBRjuWu8hKcPASu4xaJm3HiZ6EfIo2nEJtGJSM+74K5o82Y+ruKXq57
ZOr6Mti3QjMPoFSnQSo02mKC2pc7VfQFQCtWg5JW6SfjjWkQPzu13VrCe2ZEf6SeODUSyVvUU1t0
c7FC1Yp+AMNy/YCn8ARwEu3mxgMqx5yvJe7ImYMHI6BlKLRqTTr0r90cpIAfJH5EmTJ+s0tgTTfG
ZA5MNZD8ZkkSOvGivFJrW/wl/g6SJ3ErpzCtq99cZLONJhGOgRvR+EdnBL1Gph/r0v64CsqWu0FL
6CXL4sI9pZKnCaOFlixxVrVS9E+dN8Pd+D5EV1qMIlzDgBsR2OTi1NJQlO6ZIjuBosjW3dezEp3d
ZlHIQ/yNHq9m/1hrXctK/egyq71PEnrzKiSe2qqSvSVKaUHPzuyfHvWvaS+VC6bIkbWwVMnbKaZG
hNRQ7LP7f0LU7Z67twLNLE/XOu8+n1tUN+AIsovxICPA3+Rz3FEc952FXhP/ACwD1TBcDqbGXEfs
ipcC5+AAIxl5LUakwpdwweID8xtVmaw5HjFK9hnYdl4/blbqhpdE1tQxZDET7IdeXvfkVL8rlnH+
vGfxtDv18SU34HXUb7HlxJWbVkHQgllX3pjd+lhK5Btu1TTsiWg6/PJDUoxQVRxttqLdW10Gjk3G
ZbSaimLkyiNblVKCjDUI9ua+lzVaWipSU0OvhYu6hgMkv3Fnzr6KbyXLlAK/AT4+uFR5k52hCKqt
/fPOlb9fs1wdxyRcaMo2iDduJ83Fr4OOpC2PFnJc1Z+TXNEnYvSVau9uFkv0rXCsBQwebpMnIoPS
W3ZAe+7VbUoJcsiGgaKOWT+an807xgY8GY/QsK0N0tpdPiZqJII8e85izI4lId/xmfOo7Td2Xkdk
jzRCuJ0TjzvBhlukwcncbs2bEykCwUfsd5GkHlp7qLHcBWTKHaSKY2uCoK4DH3/I0rG3GcSHjNsA
1FoEI/Vt/02iLummXVcbQxFdy4fxP7Nl6BsZM/sUMh1aBh8h2RtIIuO5buEv8kLc+0s3bBLCFAw0
kN3F4e0v4InzVKMN9zhKk89QSgMqKr1TkNyaBwbVSm8+hh+aV4LSdZeEFl9DCID654TwB/ni2fU1
jfy2UxLCr7hkVvfvhS1skoX6oKanbilNWhbvQOWc80FYMz7rmXWOr9MboDcMzJ5fSEBd2AefOjZ6
vNVwa/GQDTk8uF7ffMfpBcBMR3D3K3XYquNAtyFhvUHCo9XZk9t7c4wYRG0nHO413z0s3yURIVHn
x3W2t54wOzEI6qySbOd2BzseYDYlyqN+SqxuZaCbhzxipNsfNOeZ5Go/7rhmsrvBfzcxT3SkM0eq
sIzwKzeCOo4nftuZwjihuDbexJS0c51XdWULuBo2vTLtFDmF1+vfGfdn0uq1Ro1UvMu6rGIODHuu
QdjXRey9SLvWPKLWzCPnDhgxvC+Qm7FSTf+C96Hcl1b1RxMZAmqeSpi4CFQqWMUwOpeybDJx6mkf
S6/qYHXu0F/l82ZCFZAE1Aa8OSgOoihCAcxPAR0LCbmuA+w1W6Mom90XEe1nQWeyiuBV69kdVU1T
5vGWHPh7HEGb2jfrGa86oUCi96FcbKIimgQcWEnmGECIOgqZ8v8FbvHG1EtrWK0LAZrqy3DJEDDP
lfRxrdK/Va5eLxXLCDYm2vRrBi8/ZD87Xz63u4vg3bleorhIK2KKJreUkaI3WvofWzF/BI8gECdE
2+nCULqIa7N2r+uzeorJ65Qo+THJH53zBzbViWPyYxneGJ3xyLNYt3iqjNKsx51Uh98oDtYxbDzI
HbyVdqfxA56eYS5aVZ04oxO4Ih9a5Ssd8u2ShcqOn8tQKzyarG6OIdRuXFWHkZynhZIU2CCFNVFa
4sTuxi29nTUSGKdGy3bENfYE9Ffa+3l4l3DOgbdg4KCoYAuEHsuLZw8c+Kxg+4QbnirbjO/GnWic
8zIqo1Ks745+j4bPITIDdZAKe7NucQ8+pXawjNwaXrZpd6DpVrKJym7htPZa2hxV5R9gBp7XjBFz
fWtWk09FpNnQGo2hKC9IlWraCEZvCRJMeA08Gp+3Iled3PT9oNQJTs2PrMhtBPTNKMvhcsH1mOJr
oE9u9XSD4QMBu0beiBM670sN4qOWHkrdoMkNnshuxpLl5bWh0MzLWL8fLLI6M/FSa4nnEOikCR7a
WaJCf3J3OCtQFi6CkOE+nFaPFDdpwHJXllyzoLnAkHOe/MAIqVExTVW8JEAzYZiV7KxGPZaWBrz1
0CAoLHQaxWUNwyRmTcbm/QN0ImCUIBHGu5bsVrHHEG1NvTJ6eYv1sobYTuKKsGjtHmUFnBjBKv6h
+512979R3MdWewpz1l495XDTlgzGv6BY0/bg4rB4izQzWBQwjajYNHEmoHuZRGjgm6WTeaTyLrBv
xbYb6Lr3SWWISRaNbHIbGcbieEaws2STRIYxe+c4QkGQDflz7fyOE1Aqi7lL03AYMXGT5SmRuvUz
r/Gc8sg4YSRoBJF1/qN4knRkYKQMSuBqLBf7EUcKg8nYOfpwwrrBV8jGZuMb7G38g1kAj+VQ6qvl
FW+yZ5k6uIXX68WpKJV14CmhnwaMGnkoSbr4HbKPaOTsuDCYBWjw7eqolr+T4YxihukXVFci5tTA
RejK1uJESJpnWt61AtcaLHABHpJa/6n96SaFp5x/auP1PT/f49/D0FnGfPmWHdpd902arnFcjcx+
knA9OiJsYw23oS+ExCk5EueOCS8KZYOSYvZDVVODqo6H6hZ1qEm7pWL4U5Bh0vFgrGupCSkkfCdg
iwmbXO2+xFgP/k/PFuPorYiYwl2uOrFU/KMLeKU0oJsx5J1DW8NJLrzNxIDb4DBXqWAwCOUQfyte
1lfQqKWq2xbtG0UKo8L3v+U1r210Vyxw5WY+BFBlCfYqpdqQB9tc4WcDR+qAHw0/pqzMeVlSOpj1
NC2CDd1FhItpVrzRCQy++rHz6lhNY0/jGHpYNrnbh9eqfsU36dnByXlIgqe7Wq1rR+o5ZiJQzitp
JLODsXqcRkHGNwaft+UYp7jdf90r63jXT4BfQBE1hRE4QBzrUsWMoBQgStsEUV8nFu+oufwglx5P
7VH+J1ZblmMfleKUwAlt3Yjy1g/AwjuAPzQ5q7rvzOJ3rGzqRZ2Ln1xsMobuJJ4IVXY110YdjjzE
Prsq9l8oVU/NzUbOeZ0jtqwDCqz9PYB+imlzq01OV747+ES3uP72y4ettl7LVAUF9jxwh6iPkhhH
98Eo8ExaBjpBeO5gBP/+yU2JMZnQ/BWDjfwu2PMkUN6JHpEQysHm2jziUW7Zsy8Ng+yyOYI7Teuc
xIwcGaHjbZzvy+UA2aGP2qoDoJVk40+64ub5STIMKkFBGlS7oGyDGHZ2xHDvgiz8arjFOYphdzYd
TJRIcm46c15Gz5mAhNZF2UZunsC4reGOxtNVG8NDBGApeQYP6R69sPu3B4a/7atD3n0bFi1HTlF9
ta3KXIL4Lyf8QK5VdcgcMlVgqJtyWTMoK+1v+aP5aRxmP2Zdcoq8u8qbcVtEC2gaYWq+L2LHhekb
Ttl3BrQI4sV37Ekd7LUpDOKLTH2opHnDUccd+vJtFkxE3cwpeLb0fzZntSStH51jZTtGt8hJQBO1
aBCAUPL4T6rPdJorGtXAsH+E8U5OEY1k4Cg41KD0AzIywiT5/jVV4XoNg2/JeOsG/VZZCccgbARw
VbipzNvyCfkiB5jDiV8uaAyDSgY4XRkY+IxfOAtOnH36NoBrg5iQeEhMapORmaY3PUD6rYLm+PJp
SNLXKTYA+aJnKgaiKkOJuevOPkTmKURjlZxwMv5uv4/3Hq2mO2+nCZGnN8uf30CxWxCk93j0bwlJ
7FXZMCBgSb5qEJ+dudaA1CgBzAK+TJsWP61gRtVvDLoiVQY5PwTRi8aKcTl/i6nPX9EnOF62gHqn
OdMnVJpQcicoKQmPX8GAJjkJFAq9OnKPvdwujOrl25nmeLQ+Ia3aFI/UFGotGKG3P1G4ojp3Cm9E
zMQCk0/hL+vMs/L9E3QJpkD4srQ/0d/zNK3F8raW/qj2dwss3LFlRhU9o1WUL6FQwCWFCM6DR5cP
jRVOQtEGaMtLop9JtaADdpS/T6Mwu+myjRREgO75rVKq6Ad1xlmV3Qn06vJkRYrr6KH1CMX9IWC6
rwV4ev+7+BnLdWn/waGVk2BLuTVeBtK9qF96LLupdJNIsHaqWPz0cvI4Y9ddEK3YTFHvW3ANSdZh
aM6UI5W825QVs5tn31LPc0dwegaTthEmGUhdJXi/33k0qCqbYuYNXjAYwAqPOouLlOzVHhDB22qC
7BEI+CvvTKySYvtRKS7Ln8mCnGGw8hLS4UU6Pflh/XEmQ5H1TUgxMxvclXiivKVUveyJIOaSIPG4
Ov+lqtSeO2Dr0avErhY8nT6rr8kNoSgwkTxjchIBQ2Q2ZfJ4xdUDJziy9zvLFN3um4dMMI039ToS
EHotdsqrfBu+glJvwvdmsVOsx2LvHvzkw254D0AplQyNdkvjvej+u0dHDm0cyjNOzPFGWRP5CFvf
JhrK7fof8NN/3ocrZS0+MK05NYkJuyMqFmnTM5/uGFY9F2pCqprU4v6gI63Iwt7w9zuhtJNXxIVJ
a9ctfv8EYtiD4paoh6yYXI7TzdWPw5gL4J0RNxiQcZcFgRyFqb02RXP/K1XbkrhQQHvON+k5d/bR
jEHA/oG6SnNdjScVs0Dxmcahhx/1JdymhpTIcCxH12guRzfT3LdW3AXwOqbYCRWH2k/0c+CL/T1Z
uq+cYb3/LGCm4OK6xJhASVluG3QX9wkyqk0HYDohxM9Iyaqj33AkGpfsX0VvGMqgAYHOWCpsROlW
7QXWzmeuk4QaHLvwj7A7u1JQNANdd8Cu5ovbAjWEEMZfIhYNFkjqkd6bKepQxEsYDhHtmpnmfzqf
8df5JF6jLT9Osl5NoGFut40zAnL0nfNypkYzH6v3EWoGKSWTr6Ll6KHhwK0d2fumXQ2LLPJUAg8c
redAa9Zuuilwk01OcVWv6o+TGKIRmLj6trCeVCqzF4T7YVgOor4s/dFVrOKt/KQ6O4iGZS62swEt
qJzG167S1ikbLQqpWvdJFT9RtorbHlLX429eCudw0HlgCUDuNAjGpj0z/W/FK+QOMUT6NIfkkRp8
yoVO4THkXB0Xt4grR7FyZz7uUxypm9gSQ1JgKahOrsKtiNPTN7CJ96Tglw7RBb80orng69A7tsms
MloETViv13ZLVBFcVM4WX7KNxpsjNF/cRETvVVQ2e27JrasPVV+Bu0nIDRV8L4PsS4Nixrwcn3iq
eRw/Qe/nR6kA59ys2V0G0vkJA5Xo+9pbPuCXOFTBwAmd/MhHKcZ8kmoeWLL1hXaOGVYk2hozz/7b
OlyU0R5v7N7LrqBEy6A355WZJ6Pcr192FOYJMCFcJiaV/UiOxMk5G04l3q77qANCaDvVCUzTQr70
4pAmQ7w3x/JVDH7dGRtxyHjoEauoiGhE9JV0Yy28yaAy7fddjtDUw/YO0basqStY5ONK/idP0tMK
OszlLab/YNIWF0a8al7RyiyI2wR6/4WRLZ8E693G1UpFSipGXBr6u2ZOnAklqb57QcRCoQyF6MTi
ES0St5cyxhopJyQ+BucLBXDyGzeuOy9jpEEUg/IcHVwIdmCyltPtjKtKReavF4+HyY/Cva0PNGEc
olxADg3lbWhnrLD8hyMxy1xkutsb0qeTUi+KXn6umUvLAK5SdNhd1MQ+VrVzP3uYnIIlA00hq1K8
Kk1zD67S+qtBtkAZPjfXK1eVBUlRW7lZhBQPBc0kf21Eqh5A4DYwWLP86pTPUm+5DKz1qObWBvsk
lgLo+jzSZa+Ci1PXnn/HaERVWKwzJGdyKLkmBorepgoGXOTCiaUvc5/953QqpEs8BUD3tjDV9lzr
SPJhlkhtf5nAP8oSJLregfGSy6UjsIxQH9Nu970PQ0GzYAQ5fpPgjwl55pdz9wtTgCu8wgGXCaI8
fnmXhqerYZ5OJMK6u+gjnlISLCMX1QB/jy+ZS9J9B9KD/xCdNM9LGfXwoYUHlobuZmLGDfSDijAs
+HU3Gps/xUXo+WChx9GUdr14VpaBb8Akl2lKxwB0Y4c1zoiTweu+NL26ls7r1RhheaWwLCM69V9n
y/ppmgUdoQBiTJmnObOTx80vQGij9W95AKgMOu2DhhCmLsnvFkAxsH+Pe0fLbx/fhja7ypswlVmM
MNFCKZDV9mD3f+4NyYFiLXaT+lDKDYUY+vFRBRv+jGnrn5+oEyiAjCwWpXQ8k6s4pPhPOO0IfpPN
LPU/W/k/vTTIg9TGN83/JNDKOzp7Et95kFsVY4oOXIm9qgXFEkQQhrCsscnbrG1/8jTU8QiN//un
uMRW7NasUl+RthNjHvkFM07DunQP0GLeBn+aWi8lfFd+mm9q1cVFQNIT/EauVr1z7QM3kLZWM3FO
QUZtAQGvJ81GyyppGIRu82lhEj1GexUklM462wk89IOa6c1kYIG78uw22qsh7TMlSYihvgxJhw+i
eEdzzcOM+Ugt+T7tSljArQ9qV22ocVlDxkOYmJv3L06fFjnPolaGU0o5L8p7gGSlINz+0xb4oGvD
WPyFTmyoTHjD0yMOhNKYLlqY8NBPOyfKAfm+EBClLOkqzUFcibcIUOeIb0ZVyyRv4T73Dlz+NFs6
I7hzinSJvWzLq7cOPyv0bxzTGkJoRcXm8xWKZKoEPVF6oqQ9ISGYzNcnDrzeq0192o34mAfDRbN7
ZY06mCzZguBszRrE6OVnKzEZZkRVATJ2hBH7zwOOvCq4ZbTAfQuMWjC9IEDcVeEULRt7UdLeaAjk
4wAIoTDEJKG1tC5Xzx39M4MlWEIabQ+Bzd/UWasLPQ33Xh4iM2NkpAjcdIrL60Og80KXxh4lUMjd
jxI+8b8oYik08iwdMXgewTeFjp9kIgiSoJ5U+7eQ371GJXwVwTKGME0a1mZRFSPyZhb0eQ+sAlfc
eCUfABKB1leKyRpVWSAKq4dkEJ8t9766Eyy8ov+GbCNuIJcMql459AZT3W8aYS7XJba0FO9Z5PYW
0+3DtWP6DGPb54OgOtDo2eZ+a+61wiIFBn1We2eP5zxctTQvw6kN9kI4+WDdulN+fjyUA9KBGaRT
ABT0nFTc6qZbdE2yC+Q+20IZ3XTJWt23LsKy53zdtsb6ltRpU65iGlmJEQuMfWGVbvDTj+TA/Dup
YF7q+fpD6WzUtWuVnYnbYQDB8ob/61Z7b55ZXRBgKAsDnK0wKH/CNooOlbTslZJcrhYc19y49StC
6bCuOPMYahlAxKgFZbVogrU0EGhyGGDGMIlUwRGnM1EzyQep7FjOm8OmOqXmLEDs/W5yy3S4fm1h
APdguyeFbe8gyUm8NRAxSLKK+jsVnxLDvpD0zI04NuRTnWEsTe7fQ/YT9GavMgkd1OWBJjcWp759
QHIx/CPTsVjBS+tT2shrDcc+3AGSILPiLsbCAmYzz2QK2Wl70OEN6vUW4+MHeMX+0C1gv3rHLqBQ
0dApYuNmm7hMrcPBtj6pg8/ZWXZGnBNQA3issoFkROdbjW2nqFgfiUHuMUui2KuVnYbgiL+2BasI
xTGw1+AtM2YOoXpeeC+290eoWVrRFW+CzAzLACPieGaciJ6Z1VCRDN71/HuecsKxmMjt6GkEOcZy
3L5y5HbskFBWtCDR3b/w7jL07ZKhBp1Yo3cqLifNoeNPj+Yw/Uaa9WbN3IPiVBZrfTOJTgZjhZK7
eLfwqVS0IqEIX22ISZ5y/MRg1WIc8V1eBmtPdjUxVPKrZQRNM0jt9x5elzdRkb3CCYmGmXtn9Knr
KihrPG0zoRD17wqeQL9cPRQxVxUwTEnHeeCLexUihbH69jHe/4eifgz1Rxb5dbifsJa4mLgmFJE6
K9Qzezjq1P82nzjANT6kUSpxKFP0UtvhyNgubuJ827uzIgZSpQlTpPULrl1cGH+Ipr5oigwYqjUE
7fffO1c5WL4c9tX8Guv86PdZQF1cEBE7nXJ6GevVOo/NXLRQjzNKUuBQy+SMNFJlvqiVnChGnF/Q
P2qwxJlxzMFNknOoyKYVWwyorRENy0j/tEwXLnX+JxcNhqnKYBkPOpKATenBdefJilxOan5bP8tk
cUO6l2l7TONTOuismQQ9LHnaF41kV9ic8tZhqPlJvtql5xXKLsdshN83fwFpi/7U2/wqvoZ77Isg
elIOsvhD2c/hNryjM9jPaVWrDSFs8w0wSbL7kQr4cluEbiA0tJ+7muUc5pauVeCLYUBWK4qqKB8p
c+2g8vuyGJysRQWm96EUj+dd+BAAZt6zHzK/Q9ActewKMF7+fW35ou61/mld9yEk9Rqv6Jh0KknZ
9ojIl3FyLkyz7dEXTlvN/RXWDKSnlm47ceFhMZM0gt2y1uSWzjRyTjzzmgildip/nJzImbCj3wY7
9vr/tbOy9/YLtbLdgcON4NyCJRggjbmRftinQ9S6ak/N+J/TRiTScji6IQ4ZBZt/XLizCsrK9of3
jdAjJWB3eFewkE2w2VldiNKIBykn06/DEBr8+fT95L1D7AifBwdIpyArfQs1gK7ZOG2ikVmVUgMs
lLRmhMZ0sywoBHdbIKRP54GvqgxWYJMb83S2JBbFOfsRWIxM44qvR9NO5Lxi6invHAEkIIji5oIA
aq6Uve4+nyXfoijAPZ6soSef9IzVU4Oz/duemj8MNcMizXfqJzDMzmzpWYs+xFP+HBnnkkd2sknm
xwS3VshG5z7iWF/tbL9ryCEk3R8Z4Ib2+L/yxQwHhcftFlIEjo+kOK81VYiijm6JVkfXs0EnX6IS
WX7ePsn9INlCmvru6nUpCdbB1wp2VflhsxSs/Uc9GmaK+iLXvDP4qD8yd7g/IRQMbwzQQiS1nkRF
yW3l/1s9qJQXo6x29tqDdp6c28XffQmRvgE6znfAckFCdIO9A/Mc4d7DQu+5fpp419+TBBwqhaaT
naxtawexP3nF82nrdCoS1BdYJ6xWa5zoTRIpEC2nAEERL9PwcmlVO8E88JiS0E9C1EXoPyr+hWFk
eksXoeMLHHE69su91xGttIFrYRwYbtETDWbi9q5Vewbgfr6oIGIf0UMiWAc5g9sxyPorG2SufnVH
OaZwO6aduj9hsRBRlsCD6m0AxhQ1KHAZELDtyA+3XqbleP4c827sYuCo0v987cakhB8ZWirSwVaX
tb6D9lb7bQk2f6Gs3weTCcRdDoc8l4CccuTtL0X/KvcnmiTa/L/U8lGD55BK93lTdgDgqT7cus6A
G6129mvmrBObMMi9xK/zmewoBfuZZRfPhgoUMxNa5hQwNHlCkkaohzdI4F1zLPMcET3MLyJlGZjv
DBQlJe50rqgB8CxhJJy+fP8RMsyVy2ku3h8YSSfLLGo0Xha7ubgXllK7KRTmgPx6Tl3t3TvIdxtj
CdjwfoVTBYfNptnifwDaEJ2+L1sYOtC3gOubI/TEhErSxiT7uvVFvh27BJRFtHiJTV03W8YY/Rgo
r6iitMo6yKD/UidHIFmZ2+iPce6FrRZzwGTscixZ6ZJVjFPLA2IUtwxm3wZNtv8ZoNXeIg+Bf04S
uP8yqGAHNOEDJa5azGGY+zdZBtGfTamvfMuappHHxvYoBPlt06feZXYMUj2bNkxxUWJvIGUlUINq
Y//m/o0XCT077trpaogHPu6AM6CrS0hsuAsJi3qpdOa4Nb1TLWDcgkZ87whgGdOmjroCSw6jKVx/
6bG/5jwZzp7QOC49fPpqZVkvw7TzWWtvl1LZZxfOan0QHgLnBNUSEB80i49krNuJMm0wWw2la0bn
0AbBgtZD/r7Mr4DVd94iQOvRj7k56nBUPiV5R0xIAqqucGSM2l/hMGwMdtfnb5u8T09VWi2zMkYD
VRToucfEXnhqlqbdpL/d6hNV9qx9GWZiVU6Mp4wLk7KZqlTzXZPw1p7vTI+s2D25A+jc9WBf79Tz
jM+1lmbfFYoTMuO5/EGL0WyH2jVs62fyhPKBUsR6zl/c8vKsqfqZrVnyQrMwYs6aq2eSNXmK23Fv
3XcifB2zG2sXo1xjXkStHrvkaQ1NaQ5jcA3clPBw+jbFgiy45+v1okILbBQ2OoodsQwo1HLCe5+B
yxHyjVljdkWiACcu//Po5ofFoFBHEiyUMdErYFHrIsHOonqAOiQ+QczElHT81A48kqHehGzS/xsv
w7MANoye0thFxMtj3gzptpyYINC+skgzSjpcFgsmcPwVd1Kcssug/OG99i2UuSLc5GpRmEAwfNjs
xnRQha7q6zKPSAwUY7C3zWLSIUzEPpdcuRTMoYzvVjYRo7zc0JN517u2x+Ez2vsT/h91Qu5X3HtC
Bn2icho4RMVduFbt1loy6BrtKVs5k32IoGJUOp08Vg1ZrlV8+Y69ue5mpWrTRi0s6A7CZc9zm6A7
slXO2p+diNEHofya0Q1u/J5bP9tDzSnBGEK3u85hSOYH7r1o/n5UAP98sxT5RqP0eUhsBl1Td1qn
FJeNHCKdL/6G2E03FbPL3ixwMkx2450giLVUaEFBppvoCywTCst23mu1UekPnDW6jcq3R5Cmfmd2
P6zx44HN7ZDsrPYZeBJAFEHhseIemIzBs+xo4o0WSOlYF2CZlbuUyJmEWhW5+v2yqkWPhQ5U9JMa
8pcxzBubw7cR8bBHYjglFc3T4RKxVlEVuwSCW+IP2UpjHdvY7C30PjRHXvKdA+DPAyz8SphlQb+N
MQfOryTXDuw43k+G436ZoLkg6a/DZtv8XIGnYY2JkelbTNNJJigv332YGjzhbEnP/T8P4iDPTV3h
zWLqF/Nozl+rMIwcqcG7TbRJYij5NtmYCUezkww84qYv8A5q0ySoO+NbbNGJ5+jdzGVJaXmZK/XQ
mVEzD33RljnV++KSwsC/Pdnhsing2dRO98XOVv+a/4LjNtEW6QG/Kd2jye/vjr+o+LZeB/Frc2lf
QAP83jayqnMexf8d6zxQvGRH08QU/Hy81lsYQsxwK6+iQBmByhvjnuO1Bf37k70PDlJXcsRTFroD
xeVxNxjRAKVlR838PPEdEhcq1tEsMtI69BSIzWfUvcPZQOVfQ6p1ICTiFWZ/u1XGXTAWdVL9ePVS
Spg/LRpISrl9YfN/RFvCGoeFAcsXxq0U+V4EscHNX4RYY8auhA7VYAMLb0aAh3aYuYfC+BQJzlUd
dh0eorssFvFtoXcuf/DB+IYeMQDWgzhqzPREYXZqWiyBOGDASFLLa+fSNrDUQyES5VQBA37+U/W5
aDmpbHdEx+A0vDRvrfgrev9/5Zcnuh2e5C3ozKldyVi0PJvoMNJhw34fVUEKn75o943TmHdBMHi3
zKDFIhizjAflcsrl8iVKiEieHgZaZIo/SALs+ljz3NqdnZ1IKGqqsBvm1TfD2dHLFXjuxZrkzStK
QISn2naWaY8xrDaLVOhs0ImaDCUMrcn0l5irS1H9cs1ZHircHEufO2K6eua1NZ4MwUJ5TVYle0xm
9WT6ZpXA7VudsvqCweNz7m9zcexNZh7t7HNh/WVMXgVj/nWqTqU6p7DBSsJfdVVBOmNafTTMp38e
LmcFYN61YoBqFbKD7CSVHnLxVth0LJji6OthNYmBwcrnwSr6pY5OyrJ16cvCLROtQLarKD8vxM5i
A4fLz5bPG+6121R/NPNTqqo6exddiQY+6MZzv4VkZxtoSJVKZjPKTguhOJqSPuNvfhOeYYtMV3xQ
+TOtBnPhWUYROVIiDNPjXY9zForYJU28MYC8EkQsGV4x7/ZFG3o5Ic5HmsPSBVcH1CnrFoRXZIrm
X0T9NYoESecqDv6amYOoC/z2PR0tpyYSSxvqTemNRTgSyg/Z8je1eQpMMHwCc0yqSyU+ZYbhvWAb
k4meEq5kgVM/Cwt3FhxaOpMXMe37foBu8Io1HV6NVpE25n4hPSJYbXNl7Roj5yqS0SKZNhjvNENE
t6yzJo3EyUR288/54FCd5DAKoyt7/tgeIvXwqYeX2+Fw4gnZArMJSZ3PLNVoSsAatD5BObDcm3x6
3Ph/PokuC9ZmcDhP53s47r6LHfuWSZELDNWVJ67aNzahoRgDkMCjb7AWjoDYQWjWQhtvU8g+BtIN
eTHvl+jaVzcPv6M1F88+aio1YlpQWFSthMZtQUeu4EL+WDfze+tYiLpJHE1tKBejM3LrQNf6Vuvb
d75TMS5BS1y3e+pfAf1UrUDKyFCg1gCuqBRLtN5pvDXk1PZSDmSwyDdts1P2RiLU8/ZmGvFqvk7s
HYNaFxrazMhJ1Xqo+U6P4Ku7k96f8ZntvclxhLZPQn2aoXbMFX8bfKcjflHpfBKiUCwetfs5BhQF
NzrtHjpDRglKKozPEO8UNQiMNf7RnMqmN46GzRSk6zUDSW2oD08cvOABtWx7UWRpuyFrvwV+cwvp
hknli67xpPAhg0CglNxjYBvfE9nGDtAx2qBqyJT38oCMoFx/pTpdR4n9pfTUMSBm+ub8Ux8PX1lA
SGIvPL5+6tfA6FYFlWC/qoVPrIi2krejIOW0fSEiItrNDCMGFiWRhN3B4615sFw0xYubUbaFHTk9
ElvgaAwLCIEs6HusFtn+feNu8YUcwA+s4BBAto/118P8IvWpBaUiKw6Ax++eJ7bEnV6/FcZ8XAPZ
GL0GUfHTj7vFYpCtYrAXjx4yceTpCZTS3k0NTrOWV/GyFcJ3r1CN64TPxJL8Ydk5MYPxZPwR3hGM
FLgJ+cnuL+6S8jXTzFjE9VWPq1B0EWGUehLEAvHdq+yCXktej+iKQ3Ycc015ItR8mh3U6lj/dpR5
Bo7A6bNiaFRtwVOTYprc0Kzomnu2JNPXP8O6Jt05NmOntR/bqyb3Vdlg5UVSSU8gknzQfzOaxQne
ie9RrmaWO6UsMg9C+a2V/0fPFYXA18bUCy5k2maWUnubyaxZsoe1L4KSCU1a/39gzAC+DRbDfogv
unQagAZqSTovqF3zTFq1a7wRUDrJG+KNAzIIgmlWQDSxylhMsSFpZptuxDBu4U+LTEaUO9zRez+S
aU/vB7isw7bJEoLE0KeokELh2NlSUBn6xjhaZwnDhktrPN1plA4Jl+Ssijw8HXHOzk7E9DO32K02
WOeXZhvBwkumCGeNssR3eUVVqKNao9EoA46jpnzeWzUPFUHfY+HezZga13i8BD5+zTzuh43zI+BF
vJw+xz0nHJR1Ui7gta1smPo93m7ocQr62NatHf0cSiCNQ0P3Difn822C77cAycZVlcOHzIT6h+qu
1mVjn1vIFmPYvpyg1tnAvt4cRtB9edX2guLBHp7edRBGXuoWvqphNWWlPyeLwNCL9U9+SIcA1vjJ
Oc4Z7LaUFuRdt2z7km0Dlt6DHPAIdYW5xCdVBGUb5Q53R+9uAmfa5kv7kXtl4hLYd7fOiuNhBwfl
b+4q54TU9wT33yhexxLO/PlXfCKPfFxSuW4bYTpWV35xh5xGgNp4gncLcbqo0Z78stwBilTS+RjD
IXP1T1Y8qjoRIIPvTaTLae1Jlu9vZsfEooyOcdsrYd4H45G639fLLScTMMO+R4gzDkoSpca9GjO5
S0wD7d2EIVvhX0feFcDTfWvNxVEz/cNOQfCbjydsxl3udzwaYubmouQaH1Oad+dYyKeom3Oz22uX
abt0k9Pb3qFmvpSq+biEwmUVErnK0AEMl/T4jj35hq3GxakVRbMuNU9qB067emlDmjS9YXTob3Lt
JIzjtX5HvtYA78MLrs6wEV4kaT6JOTKU5AkIqmysERK0RyLEnLPqmqRwP7dYhVlEMJar+1as+FHy
EZEyuRd3nE/OydVftXwepL4hjppixJihPTw5xrs8S2ht92NFHitvdrbgxTlJaOKS3ydVi19Vab6u
jfYsrhL/ikKkt16H6QXolb/HE6XwPYUESUdswriV9nQ258If7q9F9hy+0v1vRdyP8gkpUFjXjAxa
lhz8h56M7Xi/Ad4e1w6khQGpPO81nKSuHl80SK8X43xLWZBMbUoEQNct4/uRZRvLHh0wW9SfGO3J
EQf5Lrm18oRibwNnBEHsom37kXFImvuPzlmVU7GqzJQ9nfM8w9a3RDyY+g2pCQZ7J83DtUtc5uXX
qsEPTrNd9hJaCl17hd39CQTEJKJloqIP1CDdKokr/YMbzX/Jhc4uvJs5JVL5UB1/8LCpyUsuxPog
WwmBTMOiGgVUGhrY9+ZGbL75tgAJfNKrZ5wuFOAGaADaqLsfhsb9pcdszRfSKbswIHGGNbNZIyo6
F5kBjMD6I/4JgfpTuIXqppr2BVv+tjSv781cjuPsJnDI+UrKcongoGy9uiVlg4VmBk7QvyDb33Z8
DaeYGAL5VAAOR9+z8lxzQzz4C+G0MZZieqlZWW8LYRPOK1hxpDRqadH2uNQSGMtNAo6R2VAElTTN
7l0XZmqTzlSMF/D6dUj395b20WjFyIw90tbz+Dp8vmhjp3cYaHNzIb/P1sN2mz/nC8MYJrhsU9ja
FFHmpFRdxugDBBWB4my31NkK8+nQIsEmKXh8MSrZjCkNtD7KB/SuOzGuPo9Uf8eUMdPu3yxm9X3S
jSZWq9hoGuuuAcoRQJtc3umfg4gEpHAgWfr69rP0gvZLw1OPzI9yoP7/VZ/ze3qyjfGA3HkocfM3
WRHF1X45DtYGJDjPyY0c3B4DvZaVRlmxaXWjDDG7XNJ+MpryUVWWAueefPqoYQ8Zbe9sOge92R1B
NIvahDbtbrR86GwUeoCQ9J96kqaiUuUGX7MRDmE/9eGIpdVhrElSRSBTXWfKp56ykc4L1CjgijAc
mhKEzxAfEmmdw6wWzw49DRcpt/FaSMePHvGu3U4XQjTyhG+0Di8pJnvS8kiTR6iFUafmYxQ+cBm2
f6l+VL1vlyKgSRcG+K6ebIb92q6CFGLYrMKA+rAegqwUiRmONWfP9lv/i8aCUuFJS1/iqMiNOxhW
l/vEl1wM6ui0ihOk5+WdRC+diVthIiAcbp6rR7Tk99AhJauHLWyH72E3s0dms2v8b6Ofu44ArWun
sBuEytpbQD4K3XrML3Ky4p/0fO+zOczzyM5S7BGoxKMR+eEIO5es3OVZkQYvoa/gVdq9UfFAoSeO
uFIwjE3tFxrJlrm4yS+R32krDgk/Et9lYW6sMx/mfVdLiQKGmX5cjWvi+p9VqGz4ct9F1QRANTeE
2c21d00ZmneYyVeGN2zkFz/GHJvKOvQvb2ANT+Zr59n8FR9vP9sKy27hr3wrN/UECsktyWUuNdL0
TgUHhblWoGIjPWVa4ATUXrAREzmS9j6D49GewONnw6wpqOlPUlhTWK6nWd7HFOSBOgNojtXnM6+n
nJ+BAni8Bw42zVsUHIArobC50iWrVo+wcI6ZRsi80vd59gMfU9vL6NNYJWxbGQ+lX950cU8AVHIM
TEV+umxCGB3TKcokZM1GQtw3M2Sc0gTjATQqAIuHIJiG73CjtvGsIO6c8hNuv9w0DL7sVOwW5UJQ
4+P/PYwLqfPKD9xsFIYus1eTxo8MknGpiWhX0sj6YniGYtRYWxjw8qYhmfu3/TxjxCYXLhkOnxbG
UWq81BYgSiUTW9Nl1Lznpza5nTIf0Hvpt1TlowS0nC1T1gBwfEMBGvnHTNDN3/nBuChTaKTRajWL
bOIk4vhOiWOR/wuXdDrFcCAzwUsXafBJ30hM87/lO9VlQxlh+VV+JUd/DL6A6gE2iR2w5XMDq6DU
nDty70xIxniNYiLpgX7wyzJ/Y0X3xuh0Elc8qDGGE8+1mxa3d1/9TBbSskk1mPi5+PC/ZUB6g7RM
Iy5RzHo+lC/ZEMi/g+YaXdaU7jnM4QEe3awdRKxiDfS+m656tKavZ3DsXZGCzjayS0TAj/k9ZM/0
tekyhy47Y+z7Spa5p5cv02oxBvXSGRHVSAOdD9oZwS6eUvYnoEw/+0R8Jcab3cpuFa9yNDHHwve4
5DQcy55jR75dNS8BONNhwpj4U5xf7j8YoS3zz4kevR6zSO6F9nwzGG6NCm/8bWWztLLWUJjwVHM4
aCi7hAPe7IYdfF9JxxyxkGRd5f+BmMtlsYvW6LYJ7UB1wJjLsmMwzdam4B5vpNzS/QhA6mu29O0K
63oDuYL+/6Eq8MqcAzteVmF8wOvMq/pUVjJImqaLmXwNrR33ENbPI/XcAIrazJB0zwa8UNkSppLA
5sTOaVyzPukUDfx/z1qnjCC6aiRoafIMNe5zDN5SMGToj+Lk5Tj7m5zEYLh+Jds6twJoyGiiWHB4
sVFFOIUn/jPNc9ZA8sfXDoPHSnUvPXBsoQ4Kqdl7+GphBrm97fRC5wNruPhrxreZ+Ro4DQoQMeyN
YpKCLtQDojzMp4gHFxF6kBVI/b8yd9B5hZYT/4/ACnZZT3H2Sd+ATjrbks32LTETZRCnjyxv4Nat
ixq8991U8BllarfL4jMM0Nc+47XZtnMeu7Wf6P7mTkbayxKdAbyfaevjr3OCMrxdwzvEl20d5mRV
JYPG/pu/veyyaPYpdfXcyciYsZ+hHXEZiqhNt2DoU5P1wfHqyp6+7Seb76TnHAmPqEdSkb0J3ws5
A2TeZcBnU9zr/xO1O6WN3NjfrmiNtgphzgnRlSdd6w/JfUIYqDU9vPaFAhot8qzdl4FXc4sVsH3C
wH+7pSzX3DazEDZYCiKi0+uyoW2BtsZCwvhglc5QQ9QZkOZY/93l1uTKJOvTO9qF5tdMaD7zI7+D
Bcxlg7+YJB6fDjgETI9nXUwODF2sx8mqg2cvj/HlzKMKOwHElYS7yff+byRz9zVRuN7BMcTaDGZC
FAGt0j3RrHEpaZUdtw45rzOPG6wHN0NbE7+kbdZsy972/STsuz15w/vsBqX5CIiSFqjWqJsWlAui
REIGYDRnNfHEelC15M1Dq0hM8GNkhhy8TqHt3kruEAQydTBJ98V0rndJrB1m9od6D3ayFEdOh/Yy
iEP1DNlR+foYU74UFYAsYt+4ZNWQkLNvJfqH8HayN6T5NhH033/s8BEju2HNI4A3H1aqX/kuifjN
F7wU9Ajt457l1gN5AbtsN1xK+J7CjjsfxqBejMSHR6fFFjFSYqeQWdF9/R3kpz5Tol4rRAiIIaVK
ZWNt34IrHsrgyYD2kxSIAQ4FljrDnToUhNAIpoNAdXgXvjzrl3MZa8ii8eqzUI9fYCEiR7E5DiHK
FM01GP15bBvVnMaQhyuiSUpr7fcYcfeW6oiWv5KYecl1pYIeFbK3p9HQtwuVEVRaTtzjMR3tLfV0
ISHu8BgQ4iZSbni4eoNXHcK3kvzOgcFxRU066yd1jMirkrYbx1pwKv5WrY9qSInyf3RR6H+Bfoi3
OVpeQRnobgwvH0DHzCuByl1ywePvUx+Hlz352XYonAwZKOd8uAEYrKeMpwcld5PBpIpWKgcRxQlH
ZTLCVRvcqwlnkFUHZfP6oN5xAVtZSQ6sRwY3Mc1pKQ1ZjQDNG73fKIhstOMDcdhI/2ZObTrqpdA3
9hY/Qw5CGCziANlc82CIdA2jQd03n+6WKeqDQluzrWzAVxRrtGgZ85zicjWnqvKdbj8MrzfmRg7M
/fFiD2xvd33/XazU5Xr/UPswtzjit3/F6BF8dpF2Z2yXEuuZtOaWlaltUmFnqtqyF+qRdtY/TdN/
j47X2PjjLzLlyjTFXJMRTSvI1C+jGpDThpkYgisb7Xilkl6jAWX7Of8p7gR5BE41j+UUOQtPUl8w
yOeECk7sNq0YwmnToiFcNVwsLVn/vFr+MoPNnK5J9PMr9wV3gJXmdc+eiD4Az4r5KFS+nLpPKpNi
qEWyyLwUK8TBuLQOO44ijNJLb9sfu/miQ+VgCR71kbntWBxUH4cOP/hq7KNhIa7VGXZ3wPkTerpO
noXPVaJB3LDPvBcO6BVyp9wGd0L/N3T5WPPteuHkhc9txnNjwlFqs9HHQWQ+PJsuofxpR8Agp9bi
yx9YKWn9efxIXKSKuVQZ3OVu9K730r/6iJHlp8D+ow7yco2GZHVWMUFo6hANChbIRi1Eu5qd8dPk
PbHVoZ94tPrf+bdkee7EPUBQB221U30PARFrdhYopss3/dUaiwpZdARSc3hOHS/9FKPj01BoQBPt
02QPXKBXkN6ped51/g8FVFPrJdFx2zJbQ9xuezDxDschLH0oCrKSICA2CRNLtROJ9enQ06XB0NrX
PirHzAJgFO5Ww2y/HBEHawLQN9WsfJeMkbbfOUhCEsAswfTS5no26fo3hLpoBTeuOnF5DypXZIyc
xSC6s3Rdgg46x1sdLuMdhk1omiEqR/1P+IFk2yF+Bkg4nFyvY7U4jLdaOt7h9axooB8N2lF9GcdJ
JgTsVmQCA+cspSDedCrBE9fwBpakUhJ4sAQn0Ddf0HPgXxJIB8nij98/+L64W711ls9qEClxxjZH
mUKUbP0SlsjOJiXQCbC2QHbj6bX0bDKOgzkFSTZz9f9cusrqUmzYOPqrC/wCUTnj4+giceD6e2wt
7ANnjweruBKOgaeBA17dCYJliBgO1STuF5X4J50OPBYgrJEWs9LuDGMsxcr6Z13HBZC76JSGBQBS
vJeG/dB/6CkYzXbp6ym6WAy9aaQ4wfBQeHV15ex5Uj7CGMdlN70rxYcEQGgqeqTdxFT9jHVwDoYh
XPprD8BCbBtd8S88xtWOru0Snob/Hmufty5y+gLzgzILdktvEX3OD93TNZ23Y5QRM/EjcvwLPcwv
ws6F6a3oNTlkIbdoiR4lJzNRSEqhibr8Ms9Mu8JqkiY/YcAPC/+M+aP+FAHu0x5GUIRxBpKC9V5H
sYxXi6HcBbgF6crePOL4IF0llGPNCy39U9RjJ1WgNBmBgWCYyYL7xQ/Fc8Qp5LQsIg/ZsAtKp9fi
+2PSx9UPTn24GNZn7EoyVMOOBTyhxCZL+HGfktD02FxlNuSOnUX2ICOsNNCZIVITSu03xsPUfA61
2PhOOeB8i/v8SFxMvPA5un9Pyh7F/CQaH5kFXtbBGy27mgOx0eyVbfETGPBmXE5pQ9EFD3RCVpR2
KaJN28i9rPjyIBd9itx8UmT09cV0YGtHTNVL28d6FG0rnvcUFnai0bpNhz8U9YiZR72ipAK/c//C
KnVMLg4Fw2tBw5WOh1STMS2uHDxkfh9w9EmMWBXwRtLBf0JRwWoU0c7jDJ+4/+/wze0GEQckSp6k
GNSidohJGxk0NApKQpJXWJa3B3V1rkRMc1xuXANpQXamjri56WeNgoYIg/IjAeCfw+pD7fIjvN5e
3I1b3tH5gyiLHUm0yt4Pxpt66BlWkSM3euUp3azdzcQoW2QYNg9lLJatyxTkcQiKVYJAa0OKdbhg
n5cjAajfb6HUiorOyrkxttNauXjDX0L0K3DmeBU9YTVvF9hW5GaWp7OjE66dnpvorDr80Q9dNowp
YF2HHDjKUQYgBKiozUrqPO+FsNAw/T/cUng+LIlvvvBox+1pv+JyvootrIwsn3QxfOfenO00No4a
8GN0x9OlH0e+GjpWyCWEQCWNcu6VaSUaCn7802IBXtNyTc8f6fC+jhXBDPTZqvChU/7hDl8kv3n1
rp/XmC5UinCYVg3Gi+uQ1DYbldKeJhN2gjgdf7AMwW5MfPNXqJu2/amaC84p2QuqhSrOm7uVTbFb
+Ts/T9GcO9P49PFCBzL1EurYbfGCLmompyfh/FL0rOWLxWrZQOGkbdsmegaUaCHQyFhHqEuTOFhK
Cc6LRPJjcD6Uv2C85XtrEUTA5+qgy6bZ3FDEo4YdkQiZk2UmHuatPr1HpzL9VbUBTyTcb9IDaxPn
/kpeYzRpd9G2CI3qWgD+UDZG75YZE6iizeTacx1LUpqMk3CqN/d9rwM5hsMkGyQc/rbhRk3ze5yH
LLYtYPq3qHrTXKZonJEi3tlPWTFtUK2chBenoHYXEFveM42AfpA0URXuBn6gP0Yt/TB482m19+/t
vldipCZ0cIRfZhhEW1l7i4kICKV5kYjy1qiQ/r+OVPBwRr+TJ7gq8DKWPbgxaTm8jlaXsh+DhnU/
caEBSa85gvGtNKIhMUqcDPAXZ6J6Izhgw5KhOz8jpWkKbW66cJZ+GVuzGX6klODgs6kzqgD3zAVd
tAa18uzLtiOtxomZg2C/ILxft4+2pOQMR0hzuHt6vGXOIY/lbb32GcQxUOoj10Drw7LGuuJGO+UX
XOyUera4LQ2lyDAAPDf6Ivs3jcSxHK4ftzaTCbfywLYTD5H4TVANO+DQIv2WPdnqi/j6A7UobleY
fkLklrUo1g8YrENaTe+/JcsMo3LtXPiB57COIRc0tGE6Fd2dnAWYGQ3W6QWfb7Tn39S/hVmjmY3a
fuq4vnZJJpF8K1hniMqMZfYi6sclGvx+gVMLdhuAugIs2M3KHaxY2uFze9bHeYMUVR/+LnbNAiD8
fHxosvzlV5WyHk51RX5ER3WIg1t7Hc1Ekk0Db0qKs3D69t21or7XcRHWXHpiH6P3UQ5OL59f+s21
nY+TRMVxXI2Fr0NcKAMtzoO5+rtntaLeKnW81cY9brclLcgMRwkkAYxXiUuSoGPHZvHEOypzFEXO
4zTYta45uyMoqVcp0m/ZH6Jawhj592AJ/ohO1w4brhX4E3xpMcflQYIXgxzjU6ROnTLnMr0vottW
253WLZISSukbOLcQ7NxZgcOFEzqRx72Y7zzaAM3WgPuxI94N2yPAo77n3G4St9lNdhUvxm2waTrw
wCxa056kifbpddS851/YHcug9J7/6s+bmin4sl1+/unbo1ZCgkYn3+1tRt8401PRvk7jj0k54agZ
cI01YLfACQK/PKbPZF9ArrYyAebGl8XKaJycCWYYh02NRFbjGVTZ0D3PGQikQrRLzxjYM6TJ0MW+
RnX7xY/OXNK4VYHemaHSkDTS7dBJ+D2idjUO44P/nkFIsgp1nvdJLL+MdXqjK2O0nsAlb9Sqn5Vf
+7cR3YDNi+Q0iAYVQs6dbVI+RpP0TEKD2zhl80TBJZWjhjv8b601n9sR9E8pZ+1mL3LYiYp2+sVx
kk106eZziUF6R9YQ3FiC+C9RDH1rT6VWqmvd3Fan668KOEKsybmLU0hf+VmpAsWODyrE/+vO9abd
lfJAFZZURzqifCS1hJXYdKWDegHE/tezMSMyzj4E9t6fo4Vn6EzIv2rUpE8grnT/jb1u0Fr4gdd5
zOwAiBkXBP+BlztFwSGg05p0zEmwhERSUAOlJPUf44QvhWmqBTmblg8t/VFS/XRmRycqXuzGNCQl
fkZE2KSXBK3wMpCBBia/g9y0PJGrAdli9bhRKdd6pX9kWv6948gS8E+WLa5iGHf/NwbwmlMOOJee
KnVpCS/DwGX4AMB0Idl/he7qH57ix2DWiiBnb27XWhfu/yrmacXf40ICFG3ixp3IjUsGOYYCv8EI
+yHM0tEzrLK/W6wqjeeV/qfs97b1TsqPMHmR2Fef5Xt2hpe3LzeX37rj6MuIAk9E/eMnl3YSdCtu
QQZZLbsO1QzmHRi+cfqUsn7oEA6PylyIec7DKH4acQNHHqbE2GGioKN3+q80l48LlrCs3VMnE/bM
BmX5WRs/o1HHQdwU48V5rAgQDNGTlmb1obql5uEHd4NMZ4LX52I8KrMLtSpjFcAffFCAxYA85TGx
nLtwh159eTFaZ1j9sVd+J89SE+0VkaJ1AtaIGAs5f+SgDQljbu+LiiCT2mCKzLVww6KWZib/Y5VV
RWMHEXcItgFYukl0Yf/fzPIlI4kKWau10CwT+awM2ySnrYvG/1V/2B1aQ4kESvK1WogzPgglhTzD
ET2FIa8YmFJ3R8Lt4umt7W0gomVVfVLf1gUmsRI4TS85jVVY1smEpWEC8N+SwTP4lSAZaNZGDHs3
SgyJTCVe+Qp9/FKzwS5477oaaPZ7IHAJrQyaB0MVxd2xXoHqBrgFBHfm5/FVjq9mkpN9VPo/VSbw
2hUkimbejoljbYvzAmrmaXwJ4mVrSjtpY391Mx+24iTWrGsPJ7xipttEWBfrt6YXxEDIvX13U/EW
JQDE7BrTDGgAAG3RDgb/dtSiL26XaYJWf1crcxfab51MlUTvZksecorVjq5nGJeUVUWNka01Bciq
yatcol0eN83f0PbwEr0GNx6aybBcSrLTbX4NaYVr5qTcjGR7npPiA9w2Q0wwbF7/yZiVipk2cIoN
ppWhm8tdy2GuxxNnmnLANEESvgKqlHH+fzDT/LYqupY0LpRTNdu7ukRhF04KbzPKE6c9pq5gLTor
H4Pt6HLSJcp8Ciy2Pnn5VFAsBe0G9kpumQYGWLiBS/WWwTMHZDxXS0SnbFvA/L9ch7VO1tbE90hn
CY7VHW0dqDtCHbKdOTmmWW00pWGG6eX9Ja9EO5wG0pCpfut0ZpPsUrgGpD+D9ebQctJKdDTzQbRZ
3IVR/pe1TPLSH19kf/F4l4hwLdM9Z4klAdGeBjNFZMgulnc7wxg0Pf4oUQzJbqnqcF0CDQCzuM0I
3Kvs+WKLQf2efWvAtd62o94qoz+rkRKZjH8ARgDGGEJ2cYN1BmJYRZhsUi+HTyAcmpUCjv2b8FKn
I0zcCI+J0zPhblUrSeI1QU8tn1olzc69hqnHo77ZFo7eBGmrJQ3f9qwPEXSoXwfFPLMKZ3AKdnMv
6M5jVKb9hqT7U+KBHhf2VQ2o4uBVECiJ4YNwfWCQUPh/harnq7ezINJZXUdVIhNFvRV/RX7VbttL
vg3XDbNoL3WeWUL1Ep/2VUcM6XPQ0/n8JQaNFvusDh44PB6VH60UeL+k4FW7dMk+5Y0WP8zt5WBs
oOOw0ThAepe47A6blLhzNKXi4zSHpLEuw4Z98lZni7MyHiWjesR9d/LMC/yExOX8CQiTauNLwwD4
dWsRPZt9F5opzOOP60xsexQb7dtp9Mr3R2ZEKRusyb+Y9Wy/XUMQPPdSKSyQjeNv9VsFnt9PdmFK
twR3IaK0AVgEwh2lZhW30axmuq/AWdU/n1L/Xxo2sSglvQRETuKabe6aX5JkOnPTdXAbi/3O8cNt
sSvkoRi0FqWmXmxOGoxxoY78kY6SiHBDe7EVEjlQliSpICct24JHJX2fT9QCzHT3EnBURgmFHEAZ
5Q5rMjBnq0G/SIm6eB5cZYYrLupH9vlVFJ0pJ5Pi7W25gfAkyHRJ0vQElVRicaswPjSUSkOimJaY
4gJYxCI9Hk4PiKRMtvS3sLFoAwEdaP26bmOH6LYfqU3YaQUqoIf3VjMOeMgVR9vvcQnWaxyZ6rzk
58rf1IdZteBAF5riyHqiLnnjhlqyAMDs+Gb2UfCNd3lexlLXSyKj/UA74NJphYyJ4vDM0zXnWDUm
2EqLdmMQisMBo8jw1DIQsLLaWX5BO91gZonU9Qggupzse3pDYZuAPbgjt9gOZsvH0AU4Eq+gIN7h
q1/rNc2lPmLagZE4j95AUSuQHETmruXsULavzF10jojMeStkKWu6cQ688pisuXNNAUI/77jJV6Sy
UQRa9zUCVWiEBLNXGRh9rAmMY2l4lCaPpGGtCcazJB61I90dFc6lBHbP4kPlszO5YAjhpKdowiNZ
jaeHEsr/BMArw/qEnh3DZTCsxiJ8G9cunbcl9/5KzfqPNr3fob7NWM2BNcILhaQafWgbcwCgXJos
emrZIgE0NizkLKQKBfTJAtRJR8oBQex91/PxnuTx4kWIThqV2lhUrnuP7ZB11jHQDi9Jhk6aH7kE
W899rBrJI9Bwe0+FhRAeAyRpiuVBUfyZkwH9rSgKxEzraktMAwM3cZkWH+7D7SAJ4D8xF4smuAXV
/lWt1RKduD2rui2Q4wanPOBl07WBngElAeEJVBK8YecOaxbqXLy17DPSfeIGdtsPai3qqhj+J84R
E9DhjYJZjXGnHdnkK3/eJNgdBindA20IELREv0fJ7RdII9WueYr3jgmJFUQj4maSJBwiLx2VFvE7
0wqFCwVCigFaO1om2cwDqsIvMosi3TcjsRf7SWCLYVUwkX5rD8BDfr0Bc+o73V1JD3CAX3EdJFhp
QSNetYaD5kUQ6PxZSY2oo5ze6T/A5Ds6LTeLdAQWaKRV+mgKShEz3b8eYcoPSyHodff8wHmQqTp+
+LVYhQp2MW/+O9KCv2JtAcsjR4nXaUosWkGVPlUat5jQtuBOVZ0ve+vs6tzbnGLm34pZ4YoOWxDA
3EPJZCHhr879KRFbAHVeDwRKwnjxr/dUqHGu7fY9WDYEvTRTU9Pep4XX7tBFJRqUbvBUa52kls4L
h/8iDvJXE9kD7jnRNBZrnz/t6tCLNuZZvg+uzybdt2XnOw/LjYzmPTaahjJrVOZW25TsYsDENZBh
nT6+Sl2vcDmJneD0ktIteEzw9wFasBTjP+pp7Wokpnd98BREhhvfnUIGcERZNRmpW+CNBXW8K9bc
j7HfWhaD2C80B5Y6mfTStas+Vzoz9KV78KCuIDHucgZQOQMoarz3Or1JYImMJ0y6eCFrWajIXKOl
82WJmDlswfzYC/IXwjmEdxPo6Vbmp06l0bOzijKsYIClOXyrzp15mes2qbOMF1FXckV48PxJg6hy
3okj7ZtQRLFAJYmuA7XqaPb0UPx297rmMds+WChV8O1Ta4LjDYRgi1clJi6gnNSzW+B78SfGzc2s
4vZNW9665U4z7A7gCgCuEqvGPZWOB0hWK4Q3/rnUh5xWq/stdTNu25Z0RUB6pWETCKlYqyR+VVOe
ou+Jmr5daCGD7y09xqzmGJvw19uO7p+envDDUjsvZ5BZdvYEcFA11PKE233QEIWoJx8jvuKmuHRe
SfbPLAdNbAzs4Xp0KKdTO7j/WCLrDFmn++TZPFJw5osh2KvPlaFHDuCq0z13qJIPjqSU02sQzTuU
9sIw9V+8mt4kW9AekdDNs6NSLLZ7luri8Asmgrna+Hun5+td0kj6cS8wVnEKmGBeBiVydxBDP0p3
DmCIQGSZjNBEbUiODsa2mOw9h7G+6jJmo9tSmZuq8g4l2RJH3e9lfB58N5Sxu3M27WZoyIZjFWM2
g7EiSaWHSl5G+V3E2n5iUG7g5ovaEcEiX/SggNbDRwioJLXiaz5G9BAdtMvRFP04TqK6aD/238+1
QWscqLxgBqBi3L3j59L6r46pOnDAgbxhd2JLVdImBxXOUYvX9CjkgLfq9tPPEswugSHm7JVlqdj3
BZr+0ChV8qFhOuQKEmUrKAC5Uz617SO/NyL93Y12zkcBVm1avfGpVE1XAdBL75yCupGGVnNsfH0A
ANFd+TZs0paLZF1Bc0+E1a3ljtd9evpZ08IeVlzTqOWhQoADSheV8OlaKfwdiwfv9c7k9EtS+hNQ
AmqRz/UAOyq3oJDYFYgsmQnQ7nl2KQNOl+dEsd5/FCpyAg5ix2q99dMeIQ+hrlvZ+4L1lZHBUdwc
WOhR/j4NpnDcWRuvwYFUgsJB0GdHsW3vn1PZBrOJ0+Whz32BbM8X054LcwbScqVkMQTwHvCX2LWF
KLlAOXFUFISUwX7E1ziz92n/XXeDZLk5mpqOVlGFqCP7K1B8CT+HwXMFFMlT+f8buAREDjZIP/5R
yycoi89Lc6QAulV24gDTmK9ldM/KUzVqNZQXSArkNGqBDMBsSerWWcFVHsAmCKUIuVeTohmrjv5V
UkB8JdzKop4h4slajDIGBhcaMBM8S1/7gUYetW2N94o5HdX+s05XnmuqahU5F1uaAXaAeHtboB2V
5ju0ecNW7tW3L6dFGTXacPrz7LcWxyXo8V/5uLNYUD4bliJP8P+01m8B/yCflHRVr0d5XtcgWDOj
H1XXUtyjNEYpZIrn75Ovo/a9C8AD6CYBykxwPtiEIuec1BKhOdN41OtSyEIMXFpBQDJeCJnfX5Xm
MbCyuk/UPvSzogIWE/prkUQpzEuCcxCt1gdbjF07Rx5KEOoNgqntFZQGj8w2gpK4SmWg9CdbV7RZ
bZ8BFC+X69t0TrakxwTeZbkKcNRCU3S+20clBGibPB/fB6r240zaPFNP8XBEVBoyrUyAD9SPq3JB
8tY8SFp8nH2MI/VrV/wTmGsjMmDTn7QwRn4EjlbQ+i1W+J0TG5ulrN7TzBq1w03gc2BfSC0D+tz5
ltT1Jv+qUlMtCThzd7pGNOjcfo54yrX/1TkwcqNg4LtbFD05m31RlpLI5iPapLwXvPD/byPKxrdZ
UlPS3jcmGhhO0Tv6Qw9EXbGTVyxXK+vqG5jimFr/a6KCJqqR5SblqxSEFZW75rqga+SA9mXJ+e6O
I4hg+rR7kAkNPLpc2edtsz+cCWUVzqh4zE8B7FiSMLAmvRrSXX74cj3y1PcnKzMqJohnPnGRuABI
VChGh5YBU1hUNsQFdERaPjtXhoa0vFu8CR/92zMoHv4a+XSHiIUj6MzL/HecbEZl+0MJra3hrJ5F
XnqluOdIKILNN5xX4lKjZCkxnsC0+wbM3Me/xd1Fwd9+gqnNcmFgVESKyNh3gW4yAe72IpIveCxg
8zO2c1Fgbx1pcZiEPAM+GH6F9TNqR0r7ozWqmtiuf7/2dSY+aHdXHTnNdkptJUIRViW+NwXex6OL
LHlImPBqpgPESIGyWHmw3WsBJeBgwL+zSUIjs6hYULdgTNHQT10AVE2S2ErGcTqS+NlZ8ZHYyNT6
v8N5JlOkZQPlXVQpFOu5xdCD6hqW0/66RNEMeoxIY4z3fNTOM0nwsw6i82miFjvbzrmPXW/QlF/0
5eXDHCbGkmAq8jL+UdYunXaSt1SMp6IMP7lDj62uqUAPPC7zJAuaMiZXbRO4fNPBtfGTBHZ08OLY
KKfRXmMkEEAcAMepdDsiRhWM/RX6wOyf13riuJKYW2yANc3um+fAzZtoZXM3makqBgVI9E1XSctn
p+t85S0Eg+xZ5tnowdyCeznSH7qj/s6m6t6tQkLmxnOp1BYfbp4C4c+SNEZ6IlzJnWZHwh5mY6sE
wat7WP24qYdxJFUz3aqTxrH+UVffcWxLdlafxpfZJH1awZDkNeJarXN0nCocisLuXQoX+M8P3Wyc
RMg5wOPU/VssB8+Ffd57NKsjzxH65uBLiRQlGDrTUwioukj3nWd1PoOF+ECvVKmBf972b9YO8sD/
qoJN16JXmedGMyxqSoXOIj3P/Lkr3XdsvmgCZHzdmRg5LXJ4bIAcxf8V2NrPHqyFdsXLkdHNhmdj
iFzuDSSw5Gg2Vkk08Bw9+QwG4E+AiCaQe5V2Y6lMZIsJGtrXMGvl0W9kDMz26prOYe0onPbY6VVd
Syo8+2aHJHslAaGCDdW+hcXaQHm+aTbjRWDqlPiwxzl1ldIGo/PnqrnpT99fTND63gNlb+1q0sxr
FLY+xrT8CE3FuKsPWpjHpIWo07yPMKZXWtOSgvNWdtEmpomXcGRcwQw0c2U8Qf8DGmNya0Z995Kx
IA6nmvKykIbYwrnKxcKUWByUUYqLUS0/cfLPUYKmWkNun9AuSThEG28/IdMDo18iiX7cmLypRPxi
5VeKHAgQqBYd1TyIBjQUstV1ZfJZdyTLy6lCnEYGj8D0WhmtU+c/ZvmEUFEmPS/b9cNBHFG6bDDa
xgRu28DBVlXJboh9DsvSZbmawJ1jYKM9T7i8jpi2Grjh8saNWajrvybgV+HrOzuXADfvtwN7NDp0
gUi2nANO9Z9WvDvKHG9teSQrPdJ9uYd8YOwIeC3NOnrv9WENHtxf+5fGbC3Ox4dV6XEbUodg6nlu
4sTMZ1Md28oCOIOMUs6zXO8LHyQ4/i/jKA/9IK/uHz2otbd8jp9eprr7HNrBWdSW0vM3nCm36tjQ
AgiSdNjF63RD9Z/a4uVdH83FDAF1zZZWqemVL/ydxDMKHh2K5F6Vn5HPYxQJtPaTrGIEGfaAhV2v
rrLTwo2HchCkE/ls3IB7XlFTcCJ925bRfZxnaqTCbHP4OK7r6Bajh2CYfn/CwPOIQsJTqGZ/gMnG
oik6wsqbuVomVyGfPR7Qq9iumS4DfrgBC0+OxEF87gVkHrj2pya4x10t3g/Kl0dltKjZYw8fV0kc
bMNODIVmwRPKrfG5jbIRWhB7XBi/nGk8m0MRFT8EEz0o+mwJFD4PuZba0qycGBI4XlRtyqbrV1E0
6MKv3Ky2kQ0JkGV91S0sc1X9eUAOaqifn9sPQyGmmrhK7RVx91yP2QObcKhQs8hqfb5k2PqZoSIr
+KjLUYtSKBJvKDDmD+fxiAtzKezS0+pQoIXdqPh+Q8jCKgjiFovMOY+Z0HAB97pCdIPjH49Xp0Sh
h4qo6YncLNUKt70f9+p+zktmzBXEwqIULuQJE0yrdWH0mAxZlYTEjXOrOl3K64m2rC3SQUs0AM+N
iP7P630jwqzKrf+8QCzehpIum3mL5fagONIvaHTWlfw3NXLkbIu+EKbxoay1dwnOXwmffsVeUohn
ceq1ipxbSK9ayzo9EjfiegyQb0Y7B+OVn42kylBLW1K4iseKAdmp8juxl5qMXeZ2/qhgBt0mZIUX
4xxahk4xlEKr9cwrNkEMRDFHl2DmXsX6QW2qGJWhtK4dXTIvc5w8dKB9WO1BRSDnaZV41UzJjSsM
kfeMHV5T83WsZrRIt4u1A3Nj+z0f4wRkUAX6+T85RQqNV1u1kxprKy4ory3OFkvrs/4ePyNKTZcW
45wKPssjXWo6A5U8+dIbgaGRT+oZ4GDu3Gsfx+ESCTa0OB5S5de8eYKzohmi6MTEIXvQQRNP2eOi
zh43YTWxqpr4l7vRFOhRuvwVSPLSIQ/GRc49jV002RddrzUYyai2pC1xFf5ljxmuwXL3nQfLNsyG
Rgl3Shge7GJpnzsh9kQFIhnoBWgww3lC4eZL890L+nOeDQ5GpBio23Yzr9PZD09bsy51xO29P3jx
fZ7bSqvT83ngze+NkowYwHv1lukRMYKSJsglow6F3ZIpDk288tH9pwdsukLAgAjiGHBg9pbZxCnU
f+UUFtENiDyL/UKorH+zGotA7+BbxLJwWDIRJZ/6UMRcRPXfVBBruf2Ig/kJ9SgAvF4UEFe6GHhc
kmEKbYFdLAmX+N722K/Vbzd0Fxnt6dHVHLCbdrdNdFAJ7aEjo2WKh3LeYI1/IGLuSCzOW5TktikK
0g21nO0s5w03czkAwHEMlRLjWHrYL7gdyNm+LIIvfDf0r5ASZtimdsUftGwaZ8a17XIZen//yyiU
1FgBCxG7uEOHP7tXqFcvr32PmzU8CksEX3hqJLmq/lE/r0LN53BLgKiK+nS2NRohBxN4tXS1pstO
LED2E+NZHaWdK2R6+iReqXP+e0e+zHVHWanxl7LrDUado/pOmddU+p8K7oPxJCuVZlz4f042LUvC
ASRABmPJwemnzSMizyP5iFStYfaw1YAVmMS2yTfjifu724Ir1y+dvoqOWl0r9C0K8Xp4PpuQs64Q
GAnLFAzKAUnGvbB1RbaLea7CWGXNMN+EjlyQ66Uaby2eeFAs1ayOBBPO3kTsyiVLJ2n9ze/+YiFh
UiLq/SH19ECRfQAjsiZ5KFlDHQAgiwm++2k1W2MB0cmxGqSOnmbx4o9r+Yr5zUccBJnxTJDB4VAD
uzz80Xnane9fzB4geOjl5xb0j9flZx+bSx0MyM7/IULs9WTMO5gRfvr1fnqGi8hzX1vbFr/SOrzO
1wyJZrJQEF1M0R4WmS6bAmbOUR+uviVz1Q3wnxfvMsHXQl4k2Ro+xFaBoJklmlI+WNVHq5hIOmGx
AY69Ft2M5sWp1JOHNBMvefKu5LXxd+fPqedU9QdF3kUdxtEIVq3W27/fhO5a1JkD4CVw29on8uHJ
q0HMyWNfkd2ko08rwklbMvJiIZJEEY6zpc/91ot3VxZDOGqAdq60n7cDl0EtK97btX2kXwKbnudO
aW8uKlTyhxKnMTaU++TDPVx0l67tm0xPFe0Ol1cY0L0swxKV5H15w/Wj3Y5KviDLuoftfhThC3OP
k6ivRPTWKkJfu3u8xOujUHEEgkPmRjutAvz9o2TX9BU9sGBfY25vo4aoOXJ+NmQzGjy/GTA9B1mr
MU4byFkSAG3V/Z4N22owV0M40TtfwDfCc03RX1vWqE4BorpEzqOpFDXE6Y5kWQUyx1FuU3O5dNCL
eqL5RfFPRlK9ofGXo3zkVKGzpViOJNpNE8RACbxuPhJzdSOBbReZRzz7eTecYe2FlHXE8DuYyncQ
QFFFTTyVIqz8TYitBNwFXR9xFfMtjg7rjGNYtAm1X1x5yvfg/32Saz83nyWptK51I7N4enu52BlU
rz1f0tH8n52tnX4QQs5PwXENlJiCU++F1DDodsuLml8puCBe2OsR9DZro2NDGYhk9bv2ydh+rCeG
kpFZa4Gh4xHI03m0UPoKMZmKvIKtwCP125Dn2rCIuoh1ySdo6HpYmyMSI9+X38TyHce2Qp2iDohu
9pLr4a3CbEbcjDWctvmANYnAqZQ6R2Z5dCs8iZrv9C8E/KLTk3HxsJU8qGmkpZKqOvpbBgF60nj8
aJmCemR5BTMKcGnUz7V5folVceaEm5BBCjkholUoowkfgq1oSBusVWRLded9Bm2Ciy/wfjYxXGHt
+yRYukp0YdW1Wg6dL+03kl37tl0HR/lnmyHVb4divyHny7qIo6LUlVE4WyUMouNasytgToTjFAad
wk7gGQBAGJK2H4V3pYaiQAyTOfY2cEn2BMwlAbp50b3bHFfaZILe3kfgyczKM8yrt50iVMjqsRSY
y7Pa4kbfduO/8exgSCso8a7+X/puTHc7pUD0jFyvcU44C5hEPYuo5wilJwqp0oOA79ZYtX6sa05E
yAeSaT2DUEt35ybuEOv9FBnJlzu6SO0LIlNxaU5f9X+cMgXW8G+KMqTULLbs5tPO8EWtarJiDScZ
4i8Rx+xQKbhYhDJJ8dIG8OZIKK5q0e6tIDNkH0YsGTLI2RSuMrjHlVjmplS3CYkXFx9SgrVlEJ+j
u+w+3so/51WB+17su1vFtxXYnUhq9kAFPEl+qkW0VSPq16nasYttKsyAyYg7hZPTaB3o4ADAi5/S
DJIJX1wUHY4pShsl26s1h+pB5WP5JhrnyZY6Y2F/2124GE+/F1RJPgdncfO4xyrH3pejOkRpm5WP
1D4pdMfJ4QYmTfQdfpJkz7TCN19H2RSzNZgIwNtRRhMrej/UnzvYUnoiNObP8ELPlqPjw0ioETGV
4ZaZCQYF6Sdaup1dddspbpcfdoOaCRa6f3EFkUbxxCj6Ipx1bgSTvVKIO0phahB6/ROaCSbCf1Je
iCBMD8qqgqthrBg6god+JGbiBwJMgNLfr1hvvUHNqtC/fiJA133fB5G9xKd9gDRlOFf4OFmDs91E
kFTNTBY6sTQRxkp2dm63CU5QQh2jnAxBMhZosHz8lD6GIw9q3KAjakYjDhB5Bt10f79iQWHC/L6V
wEdRedSYcmQZQGRWc/c0HWp0LBzbpGDb4okO4HK4lSHvDzAh5dJqMYkS7igaOcW2qJt37R142esC
IXJW2VLBlQda91KQ+utUm38rP5LnWNMJ1xUppBwMsZPd277dA5qt/Uq05+HGjppHE84NHXczLUv4
1RfOsBFmv726ZbjcKtIgghrH9VDeq75/DtzwEohz7DiX66lXhrC02KTiAyLu4w0QZIVnWhuRReuV
+jVMhtJGZYr5AnpCwPz1zVgLxsJOy44FwYQLR5nT3eId+rgMj4Io6lAfLung/uyHbTjLSenyts+N
AF30GWIacEEqqk9bXfA/fV5AYkAe3bWMdZ3QLPFfbu7FkWFoIvUA32GVVfoe5rdOUf9juD3ceS7g
5OMUWT2DhMGRLSeKJbFm45OjLd+cz7Ci/JuHpFpXbB08uwtgutovw9jUtg/oyRh4GKVv/SY2CiGc
MhIQplm+2NuoIPBS12xOy7CJZPk/BIN2jYcTM6Xou82jfeQvbbSS8bTKliC582R11LXb/Wq8FfMA
H+INY4qjDuaJhBG+EPU1Gmsf8yb//CIKA+Hou1FwkSW772Y7rrOsvWIaw6/n4cASsz2/hDOu0QVt
/SNX6lEKVu2kXOiFw0eRl7pmHlroI4j/XcC1u0oFfqGGW+sdfNbXX1QtV16H/jxE8Tla1Nb4nNR0
uGkPE2vPq1NAeD4E9CNNjWK0M54pAtTvEisrr1Zh/ljLR2bjagseCuUbvRULe6Jtx9QcMHcN6mVl
21yS2SMet3xbS+30diZZ6UKdtFwPa/JCk+Ds1cmsY5T0YMoHp6sEh14HqcpHMFRvDNXPiSN+cKuA
gBXIQVjuQ1h3vZe+hb9VKbYmwX/TNzeYldprQOfCDcf7gbvFCA3ZlkW1WD/mO+5IlGMMZUNOyfOD
xnL3yncYyGPL77jKRqMOwWgoWriE57c4rwxaYrJipQF2tbDwk+IPnn+Fmmk9lYmamJXDp+iJ5FTO
nzf++6wpNSy5j95eyLykQLogAuBHp4auOxBpDJkLQX5h9yiOtXIN7v2+oFQ4AitH4Tljdf2npJoN
mDb1Zv7Hts6xUQEI0oUjAHpsLxEiOAb76o14DjTfkFdCKNqp//vIrTXq7aPyODe7tLNNjgHYa9Z8
eo6Ss1brF1TEhx8O7WMF1YTJXxsOkTrsmV5WkA24vOwibKycv4MkEjiZTsF8zLG0C5khG0Yp4cBH
YyO474JV3nGnggZ2dSRhZLZInNySJflgJW1GAJv9CTSRccHSrTose11i2cfDkCZFVnKPX2M1bLz6
LSa6VtiSU6+lWptjA4HhAGs1VPexK9CGi1saFLgRCFnEmSXLhpkdnxyckez86hXxjYiIN7vB9xNJ
BAaFKGTOybkMl5I13LAgnM7+AAM/MEmlYEVre3Ra5rTJYSPHKenUicgLFGl1DdHuLq6qqSI3OXCf
OrtIdUoobZyUaos5nQJ5k/HnbVC+PNW/LLUU3WSKdBrh4DZeQ+ungtnRIyLRwUb4HvHkZbGaINmt
COJ4Dh2rxSnBgyXFN8NUiiFfzdH2fr1X0c0eBXCDRYCarNanXs0A4Yk8Zj3S3PFzo7ohJnj0CfxI
idbKic9OAbtVyP/bMPGBmcO0wLo6/GkJPKYQ2Khe/zmqTw9CLCYu9AWW+drg9/wZfuyeg1fRekGK
0OkPPPHuMqyTJIkg9UFa/TI8FYaMtc106gkyS6Z0pPsBKdJgpGNNxOL4G5USE5GxSi5IyLS0FzCc
1RMz8M1xu1ygPJZ/Gysn5brOKDt7MBNyZ4ATdBnPdH6arQqp/2cGEZbSEcwvKgCSV0yvuFPfi+gl
I7wuSh6STBWKnuDkIjqI/f1VcMjX8RP+qgz/mR+FDKhXcWxqs8/1GJK21FpWJgMpDb6uiXMOmyo5
ZqMqmFOeYxTkpaqno1M0yDr79pjqyOSaqIFT8TtjmZ8qc30wTYWN6GI58coooXBqY8RNRaIGlQ5d
4ULkW2nHLX9v1Dt4jv9P2KgAzFx4y4CIFAWgxTKt2/A8JAn9G6nO0cKsfLE+wG4XPWBRlbaCKjXt
xZ4HPoEECOa1NTIQwtVICvok609z1sCPGX6/1b/nNFWyQeCEkAEDO2M7kcrtGgU4JF834l0bYDK1
UJPju5LGxY7TJ756ezhlHzgIZSEuAiPcKF53bKRvPdqzoAyKzOVPemE7dGHZ+eS6hbjDTkILnpYG
l7lH4NFdnvkZTQD58Ag+fHdxgITlX03nuC3xpeUBkL4PE4+AHfFS2r2Wraaq/tdmCuVIJPno7t8T
tjhB0WL4D3bCLnotJsWR/rVELn1oU+8O+a9Jl6BUFr9SkchBKTUMVy3OVp1vGrDUgzeBnNt1r/Vw
tUOGYp/tJ/sFWI0OjEmGD7sKh2V/e4tTHTpTT9duisu1YpwyOMFINeQByjPp9XATG7RsFqfWADtc
pRtPs/jNW6aJKzmfCuuKVdBzzaM+OSZ1hZ+X6rUFttQBMpAO4Z6reaMhDoRxXe9zz+eWYHufHf3c
eGqNFLvFdrodx9zXfswTXYXa8SwkFl2xZlOXnjJKSS78p7PCO95a5vhrKlFs5Mse5c6hQUu9BG3K
EQKbAFyTtJKbfJ8g5d4Aryg+mGQbV1a4IjP66FSY4wr9QUAXJzuluEDUX6YE+91xqFeSuyx9WkNY
vErBJT+KA5tVQN649OMfqGKxR/aZXajm+wV5RRQHCAqJJhlk0XkN2h6VOeyWJCUppcsZvKEHEwbN
l0zzQQ+ZIqGYsBrMx3RC5x4JUeUCBMTYWx7gV4z+9Hvovpp1Yyi6PW8QQE4n84XwgHcwNbYAnmN7
j8IFZKuVyGUmyIYWzLuLzHmbBYWSUHGM/3qJiEOHy4yaG+0//1XM+KIr4GqSDElltS39bSVlDwjS
ujgoq+GQsPk247U9h4ZJZRJv2a66Vf8ZCUwiHJcbCeBefZUw4uUWI/3rZnJNomTbLXiJazcr194I
A7deNmPknow3WrrPc7AD9/AZfbwrNiLKleCA2mRvWDI4dMVEXgrWxEsMq8nl6Vbm6MDA/wyhStof
iFR+Viid0RjWWd128YX/TqQyJaT29M7KW8OE5Os8S77EpBDFOPJt1g1rAiP3EOg1oVhXrszeS+JE
JYIIIrOUZK28cW5wCz5CqAshChhShDHesXMkpP5uyGqlcA/HhQ6bJpNRCdYlF/WyEzRVwxBStvQ4
HPW14ODPeEe51Cjoz1/Q5F4o+62k2ChuP5t8RUDJFo1dutHnG6VgrVCSbi4VyeY4KHVCxsgbhdQ7
0YCphsQoxJ39dEirgWjfcUJRDwOLBvdyCQJuDKL0IbqeOtmTEy77wRcrEhnaLv309gzoa69CwGPt
iqO1jQcH7mWtn1v744BWrfVm0hPiXAKcbWnQXRpnn7Pi1XaLEKuzhmkB+6bZ8dOmNcNLCZ/qxgAN
R5GiXOuNu+r/kEkvpHeZJAQoJBVA7VVRBlSik4T+xKyo2ZEariP1hvEvaqa7uw0mYhNf9V3J61oX
HuOLoI/VtBr2D3yZsWvoDsEVxxolOFAc+vDzFdqwnIfTfLgDEHhMJRHhOvLQ0KqVpqzbctCp7pZ1
bVqJamnXOeV6ZZ9e2AO0vL2iMK6dmrxA33CZtke3ifUSIq6PqKeuXwIx2yk8BvZjzIGwtimGlvej
wu+keayy4Wa6opfyzoGAb7/TTy8GHGZFOY3lgsgpttscoL95rAYJnii9IVp3Lo35zkQ3edG4YnoE
HP00DTL0SvY3wvmSdAzJk/ZcLRDBHUph/8f6va1DDJc/Ax61hT2cZ2fYhNpfOkda28pv9aGtEl9x
ifxAAuHai5QPJXflD5vwbMXPCaIWGs29YUn7jLa8LnEvtxjxL6MSPjQPU7YPqXpR33Bf4jpJfBGv
KYPzCAc1mUjVI55KGfo9w9j9M7eqEEN89RFaSQdv3omGQT3KugVlsSNIKmThJ8PDB+T7GghWRh//
yv0AU50c4uP/aEb5i9EWwhfId8TC5IDyQ9wXYZTahxPJvwzUrTOa6wcKlGEsFtFuC13/F9Iwp2AO
6iKgyqOpw0yZbQeMGVcTnVtRXWInu7ZipC4fYhIpfA8IDwoqYKV5rkrqt6wYd7PpswJG1v/G7uQm
Ql9gDWoyMkeQkU13IgwMkL2sCrYavEvesqohiDE5ylsosXsl+GuAzOZp/6ZTLrFIug2r1Lfu8khQ
sqcj8K9NKLkUpWlySBX6PFpwwDr9wBVWM1OJxE6U1nnWM07AAcJkIOCoNyI4VA/tuogiYVfd219V
vh4tm386mPG+/oiaYkMVMcTPDKl6QzvjpGtscrR9so05TXHLPWv89qDMBNhfObKFb9ij9aFqO/T0
Ude2oOQnpPtRdmRsnSKX07g+/jqcvy3ySzVodJw6kO4Lhw+y7ixWephaTxhOeKMIPJCieaXQzIws
19It7dVuDXTwiCaqHt4oMAkBrqGQE2slsfYJjPSYltJrUq1Sk2pmCnUt3RvLuMgZ4KgqevaAKHvv
S6zwdgZplVVzMS2n2fTUC7aCnnmalEDKas1kmOSjCXbSZVOHn8XsDkO5SxvaC+2eXIuqIu+QxVT7
Yiz4IKCl4bq4f74x4Qg3rC+elUQ5Qg7ipSR7lw1OFHkb4LPWr8GDkMCLon8myY+gqSv530ce0Vwa
xP1Fx3NBI0kYXzRv17mwjmrs1M42AqOvbs3BfNImLZMuRSPuvVQvDJnr2CIZDPkll6eSlRoFM4Tj
+84CqLNBrjIuPMV21ApM9NHBS/F7tRccgycw6uD5tY9MqKAOKB6dhwXKgSwnk+vzyYDTPhUU4sI8
ECvxRtjv5+Qvevp+RVuBNvhhHG+bUDaVc44XtxVcO7Z21xDRwvL9lXT8CtADRMBjHnhr27DYJas+
hi7vtP2Dc4pvZ2Qpr65bKpBYLdPK8Qta1iQZvdOmF7GNKgHCMFYnZET2jc/jITVyijQa143+wDes
VZr8P4KVRM5/yZLhtj1Zb9PVtKNnWDkiDGg8XO/YU4W03bneghos/mUnoqUNS6CfCfmj+4LtwSTm
8GU7LIdB1hOk1gJJEb7PX0hLXGZPQaWdZo8kFStG7vM2bdZAyJvYpS9rtzUIn7m0+21tCT+U1Hzp
wIct5NREHBac7bCPZuwY3MDX/vCb6olCjv0Y6eOCoc2Aji9rn1UkuUtjZEz/ZCxWnBZFCSZl53jv
16epXb+CbnN3KMoL3VJK3Yy7U8+GO4TsxP2rrQemDB2oXZZmOv2l9JqyKP76x2yL5nVWRnXXcP/y
ztuMjtTkRY/UX62bVElbrgSf+vNMi+kHxbxK2lU8fuV2iBTXmLl1gR838pSCYYwHZwgmTnd3WIFK
tsQKOd62Bv4+kAKySaQ5xmYIeSNljrW9Nsi6gPzVbC2m/IESor64SsUbLRS6WScuqTV/ek5Yrg5d
sd2Am4gj9WTHP0mzfzi5Wo46lGsLg8AOkga2NvYLVyyB/Mu1QyH48Ecvz0RZmgUbw3AZA31Vqw3i
GorOU9uZygVXnHp27QA+ii+uq+urFMe9hxbXEHUyXc2qor0PwbDy1dYCXVnrOb4UuHoo6ZkRmQIR
g0yQEumTe7FVkqE3zZlr0tk7iHYDS3SDvX7TPgh0iNRbWtoTaNwpTTrq3E5kWyddba8Z5uIEcF6E
n3QrubHSbsTBgUstZREQW9nxeNf/LqmDQ3VSOc9gjum3N/rnm4/iWLowROc32vWgNZK/M/Xu8xrv
6C5Y070w0c/WV79Jbn1yUc6BUyG4GGvgKqgpl0c5dJSKbKNjQ+EzCXU7dzN2l/6/W+obZGupIQOU
AbgraDWYIKcs3If+L7PhIH3Pzzzsuyj1Tam5XJgkrGBHsFsGBswTSK4cr3mv0zXw+EBXSsZR8og6
O469Rfsfqp2JqHVGBYi87/1/G4hsXFjzmx7SGIjd6nquRVuAg36Iih/4nnIDPbbP09ByuQh16uO5
z7AtYNGWT81gkVsNQ3CFNEQsAaVqUCF8oUOaovCRzTX12KZ5WxxycTbRypyza38seBBWWF6nnQow
oRZmWacr5uatgdjO6ZzogLWgBxCJ0/5ZkLTqgkJMD5DkHL6oPZ33eGXacgVPYnXeTqOcGaen77UF
tgdCVZqFq0fAmSv5RS8Ld1/jPQ0JQgDVSApVU8kMuMwmueQKfMnTyxRTYg3EXhOMGkxQmKihhWgr
Jf/w+WgpnbD+Ml+UKo/4gBzAea0IE+d66uAulomvfXZfEWiOSGdnmyflmUtm5SgK8AUCB94FjSmw
dUwEcrGsBAqM7Bkv3ZWAlpXRHYC1jAlkolfbRO/sVZLGaFS8698m4ZkWPoINmMb47Dy+vii/oUp4
ncKBUVa+imL4FHEcwlmy4rECf09kP0M3ECtyptNGz+4Jj0ZVWjG/DoGKIDZIuHAJ0CWpMO9+E3C9
aQeFPLrdH00Nu9WTA8DnqVI7mx+VVbmjzrieQL5i1tjVVCki8o/KySVBIhGVZB4FXx+IBwKCAs9r
MfUjhUuDIylwkJzjLzLql/5oEGQ2yTMY1/chFi8asV+GQKkGCZVg57V3JRoR6jbxEsMTRGjvvSmb
hYZN/T3CMG+fPQqFwc/rPobRO4YHJdyQTlkOkrtNMTIBH0LCBkxO7yjp4xsy8yd0vS4b06xnU082
dt3+azng6YocmjUJcxvBRVlEXS/3H7DJQ1L+Qoz3nCjfp0f2KKJ2D8qBp+77k3uVMjmB/TdAHoY9
4v3ECuFGnrfSWmeC25/h9dsmzswazC2ce6QoCXz9FLq2byd2sHBiqhWZNLMhvDGjtu5Ro3+eEjHe
TPkaaQLnxLKuycrdOZvPynZ2TtFp8chgnYPFCP/mrbpz6VaoUfZ7ng5zTBK3Ca8m0IcsEX0xCYhj
0/zgNsHzBtS1oeRL9qaKmFlEtauiPyN3oYDVW7O3Ug3lOadsxbMPmvLi6ub+C2E4J3x0Wzzi0N02
/xtzqgofSyDAALZQkT9vCNS9Y942Sdu/NWjtgB220TjNK/zh7EBdYVcUFy7twDRlvkKt8YW415/v
29KkNpOFOPisxct9T0IWHe5KD66nvztZbEa/+8RvUlZqgSQQsaMsF2MRMFXV4immB+o0y++UE2yf
oL0D2CLXSydFdlkbm43bPJUi34mjS1PH7Z+bYqJSI4wmDMIIfDJ7HFEzlthQswZnKHZULVyg/jon
Nku/exJuwp3HN4cFMFYh1+1KDVbHTSxq0iDLWSXvS9XXh96Qy8O++Pvnkkf+WBM1dULtbaVjDCCa
Ak6LCdkIa8+BX9ZtJDOaypbx4P+EVrH7+Pa7U12PtL7D8siSydiUA2+gvw/Z53AgsfZhK6I8VZ+K
ssMs6T7N0mwchiq8rXCaFS6B8UhHBu8yjCzGfyV4r+yDwq7uWHQ6urDORJKMcK4h0oNZtv5Z+rxc
UhEC218TSAAxvUWSdmByrFx4lRxL2ilhj31kxKRYb0O0iiQQdulrWacsXEp8FNJZt1JlxReWwkPz
cB5m+SB/hitdDSYenDbz4PG8M8UH3AutzQJI+zwhiYhbVkeIiuxAvN3NJXcPXJG1VLKrr5dyslt/
j7m0RKZ5KktNXCKu7+OjbyYjVzKndNjtPf+oYw4qaTbcq6eIiyGEQVd9Hao02q8tcPiKw6DQBXKN
KABQWfxFljzXJo+qJr1Pn9mcFN0NkfRme5BBGNGb+p91a21N64Uo77EMCsHuD7xGWg7dCzyR27qY
UdvaYF7OAD7G3q0ZvOAUEi08PmR/O8m7pnH2OsdR82UxlXiwuXNA3oL6UjDvRbmWXGemxfOMbNyU
jJK8lD+lDLbp72Rg0dsjRytk2iau9v02heP8yqxEg/FPimJZLs8Yu7/uIDbu9Zs2yA2A+16l1wRd
3yJndwo2x6lKYyGc5B3eoYbBOwip+JaID4uJTGBzJy5Bb1+Jcu85V4PEHfhJw0VKcnjEvu41q4PK
qU3egSKBUzzea+r/Ajt7TzF27HXdYnKh3PNs1GdM0IT2yflhlQx3rbdbSUFOx/3mhuP290dKnyUy
i7sJE10sde6TYyuI8exKnxpd3uZtBynygnX52FuVjgUbRJ+jSqKUMGkQmvX69W7NlS9HNqPvrUl8
DCXX04yqV41/ffCnnoEBNWj201iSR49XgCXld5Oj0kFLmgX9X27THH8cA0utym1jBo/sbt9clqxq
c1sB7E1QfqJI1MYIRanhdsa50+DWhR6Asej5EDnKXdLNzqt7cO9Kso/0cnKQ+mvWeTjDR+3gTmZl
/5XTyRoRmCfK2HqRM6M8YBNUdIW7ZimQGWzLKqx4uAA5tu3oWWle4/2H7B2CjBE8ih6fPZjN0NBY
EJxcSzAU3joKeuFsYFEvM/Tbw6BUzVQ/oLe8/9Ijm8HKY4trdY/IwMTjHpzeDuJCistMnMCxWbEp
jIa/1X3mrZ8in9YsuqQ5E7NEq7cWE9rCbHZELEI3gLT8KN8cfjqaD5G4wpZ2cUxBDRpD5oruntTG
u9jkrCjFs7ol/q7ecNqaivAIEC/TR+wucmIivflpCbRTM6FQIeboW/HQ+rW2PogIyuNN9pO/LlKL
fNc+/72B5PPerrLNqmSkw7oI4Ag1im8O7lvBHGryKmJ+5fc2KsznrT3pJr+k3M+6JzvTlcHyzxxB
bqlynLP+7uu1W8gXPlqhKtj5MuPdt2bTQed5ROxHKpzO5Hk5af6O11OD2Nqroizy9wyRBJpDqWbF
VQ0yEfQIVA+Leo9k6Vmo/J2Ndk5Bb61c1XUVK8boRvY/6Vj2WzzDkdyCRlaOR/Vuo0y7uYTXr8y5
gZkIlu5WZOA9JMMbXtXMwwaT4edKzosWg3+qrlJsCCezrAKblF8+x281Nstuu0yBJF3ZeKWX5yaP
PlUQ3TkJta068q28eAE+nAYkUTpADfFdemEuXvtUvRL68JMjWlvsX1x8a1jO8qj5+kqmBr8MEh4M
ZI8NogouZ5OF+RTQeHq2q4xpEsHpEukgd0XxoEU4mURoO4LjhXc3N9mheUmjFp++0j7qLEU3qlCt
gbj9nr4281/sZlLNHX18l8OSX/3TAOpCx7xRr+45l3z/u8Z4hAdqpUwrMgwmv8r/VhgR2+Dj0lBR
YX61gwsKPs9GuRf0M4ijRxR/ACPZAnHx3f4IIW1TMiRLi06RCqD9pHCRSlaIEB6eizarNes92lPT
kNdRhLf6f4MCfo5RXOniBdxNjeeNgYxDbc20/nlCuC+3jv/YGbbCksrWAdhAhHbAkFm4956BA796
phXjh6cehZb4TvAX69lzeaU4Qy7uPUmPxLVq+WfDeaNuB3FL+tSX9IpY6DOmH5GXeELEzpOkZ1jW
aZbstxE/n6yvLup4CwjihKDvQi4ppR/28U+ID6HjcXxGp3PX4O867iKh0VqFqj/A+q8g7qvwy8B3
FnQPMb3PbM3zGwXPL6Jdm4nbEw63QmD/7hNvsvKBbFoUF6pYSPG8OAeoyFEVzmrTOhgueT434lhk
moVYc/3iakV0RFdxZt62VEky7FO+hJtwaj0AluaIStQxSN7Vgl1apvnDcd8geDiKQ3XRSHpyPDS2
viOir1wp/2tEzNMcLTsKHNv+bEUU+Ur4ZwD7Vx2LQ8Oc8fHn/leYn3VM8cKxcNmxMt4ZumdrlpGN
QLkSQUne7QSG89J1XLmpln+bWvm908HCvlUZxwjLRw+P5nByTp9wl/xGUXju07O8ARtJrFv4iPZo
02+eU59/urtSDL0gAmgEAWssHLixvh336SWi3g+RGaz7dlxjBB0iORPVuZtJixUMZqzghIBYCkmK
oXBfvOHNdNUKRXm1Ff97bzokpEWqIK68ep51jVsaIO348OrgsHA71XV8TvHg/eBTCpd56K3giWuI
uIxo2dSdGI6ybtyq9G01QGPYlqE7/kMQKg/ic3/EtQ3Ttd6ItdLi/hOhNwYGHPQcvRtz+AKNtzcU
tEFqlduUhPvv/EFIs4mccSgfnc1gJ41DnrLBi5zLDZIr38RawP7NU1feeNw9WegaFT7MZcXDMjQm
lTBgBhAxTCFPRJiPcTt3R7xmHWN3f0RK1SoP1Q5gxNGqwSnqcfjIfOYoYJTX1z3QOs4mrwTajk8x
nsNDTFcPPhYwIC82VXfZeNCfo9q6TymtcbeCMxT0FcEDZkBhESSAK6YyXdF/Fkv6ag7QQ9x2+aab
qEMHUMdh+V9OHPz77mhoEMNdvHsGJuaZKotM7e+GKPviuJuyIKahTrh4CprKlSV9af2X8fYPNPqe
ZRZJvvFH5DiHtYmMN5w4eCp7smbiRGH2wU+0C2sTopMQc7/RAJUb8+HhfMFIkKWGoiu9LA6tfbGw
e4BCh6qy0hqCWbT0A3idr3ah+SaNabyJ71BpsrsryLeO1aTyS8v6WSP1Hzd267RvV9tfm92RLT9J
utVYFjf+nDM/FZoGq6iqrQOuV14lvUhPfcM+vFACmr3JVzgDZ4t+5/BJZ+iuxtnUrQxxS/IaaNPB
U92Z0Vug6dJYVGN2YVq1xGzObSvbNd12k1NnIz0HKxGGZi4NkPnNJqa7TQ2+yJh87K0gNlHfa8Zw
kCMLnqOUUyTosJDh12ApSmAxFzxjhe8VpeVtF9k7vXfXWuKVLE7lM6rqG515Z4qnpyBvFmOF7GXm
pv70ikWKH21IUpW1GP5HADzdJqFRqzpVD2Nn/FEi0tLTo1JGx9tHPHeYpx2izLL5CW9cDSpebSrZ
EnBi1GXsQioSTm4TPvLBg8XLOS2kq8eQapQodjOFccw6Bn0dgL19KE9LbNFK9dZo85LAxK7+ZnIK
A/fkTlUACo7DyAFqTgrYL8B0s69kSYp6cIqo4ZoB+JTvVmPpPyEi55MWOAIr2sY1IkjpmeT85C/M
dN/5eRHdXGRFur9pVBdF54FaWN2CKrID2BS+40aKaJgZdh3I3Yy+ycNzEwukYX83FZZdE5trr70v
+OhxOyV+5leIeNn4DdO1v7erWwzAYYgibNIxuLtu5u/pyx8dWQfY6/GtERzX7XJl7fKI/iO1dkUY
hr4/HkEpKfaOQBhq3vLGDB08CFRMnuZPWk8FTik0jMGjwv2+3gjsQAQGv0l1XpFL59HqY1j7pWze
dajEfUfQEe1nPpCCkXShIKinVEGR+PNEhGIyBL6oMeQDOHwHaA4uFULA65FbS+sShUFQknalrrq2
oG3HWeK+GTIbIJw+kJaTxoQMhTTR/ZupGdcsf6zJjHKIkRmOGC+6R2KCrzpt2zlAge7/H8fIF6RD
dknL0azWNGg37pf0kiJmVO1mV2tGSbWQc2D+4jfyyGQ58gkfEAnz9r1xMHrxM25wA8X1hb22SMMl
R1WrVnNWydQqEr6H0T/EnyVptLxtHt8dVWJPpgTq5zk5mmSoTuGdGLnFTqLyY3vE5dcQRRuKMe5a
+vYwmE4SHAM66qc8ZnROwdmze2MVEChpp0aI99tmAeP9SAu0/mk5pJtgCvf1ZddxluKWacO+WKQX
1pN0kqPcQL42wPrb+Tw25J/qK4H6ofSq/Ev8Xvh9xogRoqR82fsCqqE1lcUKBxkicmoomMycs/1Y
CopqcdIRaOomL6hRcOXyYKM/0qouETDjMsp7+5Nj0i76aEcgmMotDd8nUxrJRC3lNIA9F9TOZCQ2
kYP2a5hgJ3M5pCvfFaEuYV8gyZwj3nhM1VAzZDUfRwYQT7fFzBOXZxuEPWC4kE0/xvwd48IyrzmV
p5CauYCWBmgTHSRifIsg0WJqRMabitEudavCaSqGdwNCM5iAR+Y5zmSgdxvEhrDrC+zLqpRtI57+
wv84f5qxoELPdSHRaAAAc8y9uwwdMjtgc94mMMEhkFYtjjmWVGIQ9lcduxNsZnBt3/E6AQ5BBPgl
v2VUQ6I5SfFFAXcK6mG7xqE9XXiLwPWBZdYp/mAxPt4cs91lqQEvI7L1FQgOzpPiquLF7zvbdw5M
NMbRtLJME/PKdPFLsrtY/abIwivmKD+9bquB/HRTFcUUqReoqDeP+htYTNuDrkpwWZOwR5uAT52u
HZnnUIql3RD2Mbd/Yqe76TFBxbTJ5DuqIfca/XMKuLPEO84rJGshvGFvfeymtXZbK5E8aPJVR3BB
rXqCndG3YmnnkRCOttBNuZPID9fEj26FRN7daSPoCKzQKDixvrWEowvVZGFhmocsWQT8fECxBDvn
SzCXFZNFzrx6tpoI9Yd7gkEho24t7rrx1ZgFb6qryxFA0IT7VY5ci3lb2k+Cg6VXiwDYgcRCBH6+
YQ3kfZcELKqmgIgvEGwtj/hEBb2dMujevnPM2pfE42dPRmiUJaybj/SMiKq7Osg24IILw6a6xrwB
IrBqmlQrs5rit8N2OlpHiRgGOQLSwOvNo+bF3M5m+d2+fZxONlJHJZyyeStUMKc7pXcZCqyIdAUA
inFI95ozQNyROepdLSfUsrBvVmUiKgnlKBtBUQmET9LBVY/M9F9gV5/bthdUKno13f47w5wPy0Jq
Epy/5QJcEKcZsRZZ+bEnJwBKXz8hwqx8er3JICqTf5yFS7SMivu6pQXS+cd97E8Hv4jQwo4Vpts4
b4j/WFg2eJ1szNbwJR4Km5CBN0Rk+1ryYjqxAe4SsRPFj4z0NQsjYZrGNP2rvsY+/nB72miH+oQZ
Q3xceLpCUu2P3Oui4SDCu9OYWiWFlgV2wrQcJ8sf23gGEDIDq/vsUd/3m5qKTWGG5YmhUVxHSm5Q
3/kc2GlBCRCyyYs4P62KDK9Gj0l1tuJJqW/MXEDEq9mEmJ2JQPxuW8YVdZzBqBYKIZcQkjksMyYy
UUjKO5NNnkPD+f2jC25fW5TaYe4SG2guC8nR7iiEo6LcKGHJCjEMfDI5sDRuPP+j/fCSyz76F78f
cPP8/5/L+OsDNsjPcokBwyyXAax9Fe3qUtouUcFVCq5p/sOllPZySCC+d1KmSTEXKd9pdDK/jIAd
zIQXe0odowm4p7aUlDtVUx2VAWEQPaJzIjbeFwazKQjZ6ri+ihdusgjoWh8V4cqSwPd5+G87aYJU
JChcZUDlVpUU/t3lbiUg4sq7US0EFx9FfvMSsnANBzHDDx9c56O2GPYMDwzBCvwyrVkAFB4MshWi
xFT6zBaYIBDeIwGj/nJuQWzrepCAKJ8rvI7J/ELLVDB0wrXY6ri2Wdeg4zrKm0tZH8vc/bOduGLI
DGlewa+cMXQ9LDdKfSzxFrIR28VmkyFom1v6ZY233NTap3CtKU7Z+YMnv8rmQbUBWuaQNUBPODmY
+RX2b9EIeVSrzA0dfK0+47Npt+kkab7aVra+W/Qw5Xsxv8noD+mYT13YUlg+HCb/OYgl68t4Qapa
R9+ZNivdYyQgun3daYtB08D/E3jcm3JZsT33uCRRdYJb9a0NdY0HexrgU31XINKnVKO3eTlNwV54
cpIdmtiUZvYMRMEj8yqjo+0He4Be0/bLAE1oTNMRsZn73bYINnUdDwFlr19BcqwHKV+VKk8SBnCM
PbBB3vwEumslQjmMll8oFhc1jaOlXS2MeBgpuHiNLaAHQ7hsGxacqFRzADlt4YTqNLFaaeJn3gRl
tP18qES3OjHM0NaIwX9tVxxW2rAlcmzOn/ZgJR+7iuejG8nW2YgYzbR6F7+1WmwV+vwJemDsPU39
0xYdL1Pp5JKr7WwdTj3obgy6X2g3edobKziKL5mxXp0wsRYczEDD1wqSkpzy9z/ERwPnBfDjE9ES
/Z2sY5mdn0Tbj9BGzjujpn/NNNqfrc6wIDmDcAUWGbXdR1Z6WQ910v91Tid8dwrRlulKqqIGFx8M
Cx5R42i4PvwmrrcRaRLbEmntwMwhZ12nLV+DIyXezwPrcQQ+2ePGSpGiwvW8vVUGK46Jv9ox7ieQ
kDBeRbOy3GqIyvk2cnppXd5D5wiRFrWR7lcfWsmCMmxY8PHKDSMYslkYzo2MJ/XuV+MZSovm09Yf
DsIWPT+0/Pa/Rx6pJFLUbbswJJTI7L+LHeTyXRf/5SI243jT7nYptLHwaQNIQjDBalc4FG/uoNZN
byatDxmK0yVNRWAIAxdrCRUtJeVsTOA00zISlVRmI4M2XLckyFGWd6Ggsk6jvIyMNfNdTUzFeCNS
/GSmLsCEel+7RvzyijNfk1gBOM4/b5BF/qgmc7CUQbkgNwFpKm2T2uOa3yzaqQyLvQwRerJSBhcQ
AWoDuZqoe0dnIUfxZGXQNzpohwfFfU+zGECIA5AZAAKGbQpkRBBwjt6oVspX8F2jZ2cmW+SZXIGr
TCCKTBkp5hn+xpljnDTuWTT2dPcae71vH+QHPBhjR56IDqsAA5oVtIH0Dgp2eYGzaMQzxmi24+VF
n3R/2eTfsZ4lWSSIKGNMJhbuufA31zhw5gOnyNLLTIyd7dBej0RiNd0wx/GgBLqJIbQkb9NM0H7V
XDo9OQwbbznhGf5wPRtBllHgrNhY2cgtVYeSkGJ+ttyNVgAtf+6uSL5LoLS+R/+l83nzhII0qRFk
F4YFZ+bj82nziCCVBPsM3EY5B2/ch5Fkqni+8OVeG10+Iq6Nh1WTZoqasXHVVTgTvgNQnAyYHESs
Niub3u/HQienNL7t0V6hgwBy98M3nZkXGn+7qbEGXZVz9vfYI6qNUz2HOaR/kJujTKdcgG4MtccI
VtahIUm5OG70/Rb4cgvyiInktc1CbqVAEKN9M1kX26ntzxkAoO0gOfQ9wZ5z+XaU/jjKv0cflZat
QdpZNe4JH2qLdrH8/cxyVowCnSgpKnpgBDZEXYUy/wJz49dSJlzmrdICRxC6Yd44qM1zmPRRZcv2
bFaIvOzTLi2AVrOYlyKngwPoF6qTYIPUMEN+iXtJgOIXUJbh2Q8IRvUBE6x2pWkgKR0aiAVhN7We
zCRD7SE1hz9hcJQJP9M98xMO9H+lNeonSd5clyWvdzO+vk6vnkAdhAL+ghei/3w5sCZLDTwDkmkO
6/5VDyn0qZq91y8XmVW3NvKniO6OyOSlixHHIfBWwcplMMhdY6P7VIU548M607enQI7o1wxfVnwa
G8SwnEWFgcRFjdLP7NJ/i4X0p5MB6WYHJIJEndHkgG7kP9eoiKlnFYjGS1iCX7301giLFKAuMTBv
rkuf0fvJekiZOKgf2AyBGwWHfKcgRkMPklbp8lxcYpoa9wcyA65nPiBnpv+KvruqiR5StyplmPCP
Fo6Y4G7n6Vmfq9BwRCv89nANcpLnOtU86y0CymyN7r7lPh0IVB8uRWRmIuMTqSDxBmn1GSyQdgRv
HuD+PbVmJ0uOc37ZqWLmyByNiJAr+HjbNsDQouOr/czjYp7IWe/Z8KAXKWo0CmfwGIQrkZ61vgAR
3/+Pud1kGTbDZnRTGnbHO1bkn94ZztvEJ9BA/s6t29Fi9iFUQIIWztiMLm3g/pXAcUd/1myioqkx
m3FeGkxeXDKB/Twm3c9JIVIMCnmeyIAPzStKqPCCLDyaMYNN1lL3Up/xvtdLRJahCF0kOsa49jUN
KTQ1+kLQ5oqngP4zNl5kAD4+6eJu0PXkJBfv86TEqKJkEzrq+YjAbNcOgPulCSZJvVp35dDhsSot
/XnvDQpOVW8IoRXyto9iNoZDLTkCoXqyNi1qwbzZ+OiS7uHfGl58uF0eAPxpZnKK8hC9A4yL9kPS
g1LMmdQTRLL7+e2OeeIHJBAr7+A5o/DbYj0bujSQggO3IhS5edm9CfbKe58s4iSL9Gdb1NlQCyi+
SX10ZAm0BgcSgmAO6kLxIRke1zaBMwbkdNFJa1JL7sNAR9t5Rb+LdMjMI0A1Sm06e7ILiWkh2Eas
JI6/4Su0cg3Ng8fDO6AOpoUB45bpHnserenEmkQmD082SqGBDLL4YU4tgFPj2Buwy4Jh19H2GaIN
cIRwZxWj2Zzcb9WqTAszNN3LFLND5jrrzQuN1d9htvP18JnCp5EtKC7Yyc9myOVwo3DMXjYlL/RR
6mPYHaXccauf2ztKBH6gz9/8rDMkNywnH7Cr4A506efHVeaSduF6gDbGujx8jxCj1kzLnijcyoFW
qvkDDi0LQjNJVeBZ2RUJOC8vAD+6tihX0lNNj45d8eGs1XjSxaCDavsEfhoOGgdL93CmnyU+wXUI
R5D/JDNzTZyIsF3ekCiYPhMeFp/D1ZyRYFuVYP7PUV7W5IcLFo+J0lNOCZtyT7+YZGEzrb0kjETR
/qtc+pk3yLAKJRnFc1CvgfH9xTp3n+z1DlWw9t1ZZXEj/CMIDEqC8CVpABC6N+15WDuTninL+FGs
VKlg8I8fhXwOZB8oaH1h6mv4dElW2YdBagmK0D7NIyBU0PWwkET483OmHC6+rLu6DcWMeiZxOeXt
SAscWTyc6+OoLhWI8sJrLhHMkBC9dGekGWcUJFX7WNWvGr4EQwXRPOtZkOxAZ4ffjPfARMAs+Ajh
0My9mub0kyTr1hTkKA6mHpuYki3/RD+sz3ZJE9Apmolp3d8ywlR+aGLtBYB104oTYoVmayGyPYE7
FDgKBpHnpsrKLpG64QZ2/9gPdSsPxL440/q8DdgCLooTq9cXTnjcMRkmsI9DWXZZ4TdDvzXJ7yV9
SAFMJUNAVDC5iklk4seovoXlLWfBuZ/8BhjFvUZAeDdlV5w5NNGcGVwWzAfapsUzwlKHV/oxuESJ
dNSB1r11uTTZNeCpXxlt7S8NX4gycg5Q4H9fIUIPVO7Oex1W3L+jn3wkGc7Nm+VorjKSNNDVHeoV
Q0fnOyXRPQwhbOakrCAO61HTClY5lCNRwMDBEt4ioveh7wo4bQfNlO/k1uj012GWFIcLoZTAzwyK
Dj2Pt+gfPLcefpMJa9+Ja4yCHJhwNR1f+dC9fkeCzZzPwibMDAeyKOSda2osdYglfZKRweBRUVGE
rZ14tOfsR6Iaci8ztfBdtuEDUBsFQbWpWu4N6SgahM57fkFVIoYOgEtJXqEKWFkblfjKZpt9tfNi
60VEsSQTXHnRjgdSuIk8Dy36g8pBTBPxEWlgcK8WvpyU9GIiQBUqPtjX8UHuvjHPiRgrYvzWnzbu
lUooQVfWNmS552MEoC9m44OER+LjRxMqK4+6z64BLE4sureYajYja52GvtEGbdxRtTYsUn+GpK98
s20vthhtHMK/f7P2BqcKemKjeVSrZXW4BXF5xPfv/jWhqZZHpq2ZSc+vq/38XLlPjv8rbEebQhvh
v2AqREExpGQ2vSZcPYZ5vRqf83WMJlMGHei37BbNXsIBAL5md21WCwGEfVnlb0X0dqaxqjr/dqTK
qnKLaAff4km4rUP4ULd2D9P8ZyNf7XWcM1ATy7LDdlMsfAFCJl9pw1/J20Sy/6Wel50sXbGZHj1+
fw5rF2J68cv6MhxXy7d+Wph3OdHUo/l2j3T5VwNMdyNalfNhPXqUljumVvM4HZRkBqnL5KqjlJXK
ASztBuwL1WRPfzbVQIdvhaN577gIkstrPOpR/XmWT0gjdPb35HDmFFzeb75/nsSLgxjpD1/QYazy
w0nkt1ITxnhDJ+IPkNo9wMgkpkDamj+uSLtTCc1b6ooBR19+HHTwDFeP2KbFHZmvMonnnYIpf1Ij
vuqiCGk6TlKMKnXmnCTBuR0hnN1D8PWi0L66zpTNTGX+YNgvZ/36hBly1CsUFiq1aD8HM3ULhqQ8
mp6nEEqzUlUbb0XhawI56XK85mofopZPrXtRLkuk9HTuJgox0gcOiFMFwFXhKuE369RMSoGoUMY2
gC1wFFNtkXcFMaStwTUTzeFb1Lc6AYYt/hQJs84UPgz+Wdz9qcpPwNvjIX/OI0/tY22dpBtalk/h
VJ5M6l4T2SBzwnt64Uj8C8mnodPqCXI26B+rLPS+MCAl7tANRU7EwgCBZCuErQsgMmUjJLFL0FBU
jMTDxfW3UuXZaJGVYrVVrNljVXpbVb+zaj0zD05a/Iz50KdeZ7hJLu/tQmI+ykHmAqGscbRnfZNX
kQiBUBKtV9LJXIfqlrfj0s7KHw80Jht3NCdmQUjpyEoUsdx5HXmn7PW+fnPgY16Z3wKkSpvyPxDV
gpFN5V0w7hy44qojwcPMHbIehz8nkp+8joO9zKwwecEQcqxcltQtFZ82kEpHn1B1I2Cd5+ihr56X
rZme/tNqWiw3JhGs8g3poIb/aCZ5HEBainxlfq7XQloBU4snEIqcJ2yC/wxL69WIQRFyx99EWnEW
Rn6eiBC3ZBQUYPo0aTU/0PraBklfoJgn6peX0r4lISFiaLIHcVVd7psvHGq//DmZdw6bN7OCK4wy
CNF1b+OWPKwT32ExK/SRCWqrZ2zulDfDj6uJzcP/usTBWLks+vKH+U4r15UzicxmO7bQIrBSfr/D
BIUZ2IE6wg5D7rtONAviXGCRI50fsOEcEeWXmPdJdU2JQ2qPAJzdGxjs9r9Ng+IViltfKMWV29op
PxwTvf/M1GNtwgB5WZKvTK52CAhojyj9sjWAmpP1WkJgI0NCal3h+AXzjEKN/VL1YwJ3ZUOSndmy
QEgilo6qTtJCPDkXge7yrQ6We3JvuXlbVi518uAWpQTm8OK6SvhotRJKjR0vuXR3aBuLXm5xObgQ
EqbA6IQYiBaF6NQBfnlhz9VZEDzFCOCTsbnpswFTf4InhWKAOMLAPXLDyywIX09aMQhUQbyga+bN
JYZgwzoVjZYFisoy9yHY3UKCtkq+A3nHqJRWbw3wNqEsGUCZH/fJPWw878rB+7JRV8hHbsU5yoZX
zMoSmGsIr+8GZddYGlNYVlBIBuGoEZIZ5sdBSem17p/WZOJbHGtW+ZA6L1CjS64louv2AtvkX4kc
4eF/EsOudjaVm2e0qtFanfaGQiAL8LgH12jBtlAzZJhitdWbjOe6vSrl90IjvkRDpX+9g8a772ox
Jf0fOo1vdHdjOD71iRQhKAYPuEZwf2/Fvuw6RXwl2gQ20UeaGQfIg2c/IuCUlQQHyklfaNv8G7DD
iSweUSXkRrlA+r6pXfAC4c2zStNttJaKXTTzBusOS/HtXVCa5ON26ZF/6PMqyt2dV7KHp+aPNlSO
P5zMY6we1LD5N/KN4zlHkoILOllOYSrXRZPdBAkqs7Fkhm3jEqkMfMMMt0fLY4gGNLVkzZFVBeEB
R1KjyBpymmPZ2Zccumnvd44vafLU9LoebIGQR0zQsDGNDHrx6B1XpDGSWn+NGpZclJlML7q0D647
kolRSRxBo49vGW7sc4T5GZWLSmly19G3WaPZfOToEQFzyN5jhRwiKuHwlOSHpW6CyGyf4hlMFD7h
XHPEH1m+8HiRpdL9VEQy7NF6ZqSmdISg66KquaQkg6842fDqDUGI0AN36ia4AIraxVITRLHTIzUb
9D4UVBImbew1TmZ3RD2uFeAbTcSVUgxHOLMAnxcuVOkwxtRrCt6wvzFi31fWJVK6cuny3QIjTmdd
gfCgu0NE6vo3IJQVGGdJiCwm7Qvv0nketPWuXZ4gkk6oCAaH4Lh4dDHkT++mTV31CtdkDQzEml2J
rfl3hLD/gHajXnOBpNu8eJlo4qQLL1g7sCoWJXe9y+YeABWyrQrxQ5s37B/eXz4fx8hfBy9FgqLN
AwjKc5IaG80I4j/IGwMk2nFmKMeUKKjQmpOFVHqcpueHOil/JdCHBV87Kk1cSGVV1/eAUDFiUxYc
icX4OQo4Kc7NPzF7cSA6Id/QjJLQaa2QrtdbSupWpabR9SZw0uVMDDSJAqVeopYrU8XktPq60Fp2
jiaByyseTcugSus7vihmTL2rNvfEvmtlTRKEHzsS30DMjZNzPtue6IgdEC6tV2SQRHABTHbLaPpb
B/j3AZq5hrLtpMnAi/UsOb5S20LUhVmKbrGz+7JxJibkSDp2g4wg+J6jOge444W5xk4oKtA6EFSU
4p+v8eAr9hJRyuM4KS/YCq9FLOQWZTQqaolwUIHh5d+tvr8eF9vInC/s45r8X41v7uoHEqH5kcPo
OOvhw5VyfvUjJ4yR2QLIUcoaN9r+X2BBpqzdfPasXfMwh3el4EjKqBYda42DSSekfq334RCcdCzS
nHqRZwvmTPItBMMIMSUGDSx+JgcOrYmnHeoiWZN05bzy+USHLoNfg2XyNnhSk0I2Cs1l4cV/RJtc
YhOL1x/DpQGhZNK8v09WuA3Bj519rTZRv/cszHAaGF/DDmuSRai4CGm/MOOULo/8yp6g4fC5fYDW
mLmD+35K4bGYTWrntQrXA5MqzbzyxUsjWNkXr8D9zoOoqU6E8vh/G0Jbf6Wd+qFh3J4Ns42INy8n
7idA+r8ESwZR5rpKYonOgPM3BffO2WsRKggObV2KrVa7zA2c2jt4FOjlQMZDLTX/1wW6uMxD02Mt
kyIULiVlaonloOKosfLCATr+2Qcz6tW0SosFe2Ak/gHs5CZssqtRwKOEngxCWs3Hs5CZ7ObyC8b5
qXV4F2QhNrmk8NHaEG7nYUhNR4IqSbE4Kq25tyo81ZCJMFLH6HeQ6EK+w+4GINRsu+U250pd1mtX
kXU1LQUCPkNtfsfL1fDlVWVmvjOFHL30u/vqdC5yluSe6M2qff9iFrcgvozguMEuBhQ9URSOfBEq
jYT7H5VK5id1yoDwk8V20PjGxtaPq2UJzesPzuTQVheesE43W67EVqQhr5YPCnO9VE6NzMF6y5sQ
zPGHki8pDU4va95AB7mOiHBAX12GV0f3eMAXVTpGa9VHcUpaG/TKu+5PeNR+4jyWz0ZMNicilHPp
6AIj/y8Evz3XSDDJRT3oyf8vKIyJ9hwtP4QxKXmdl5p1fSjf1YDDk6G9N5OpGrck/59h8GbpHGxs
VS3FbkbPPk9saIywJtbvc1jZVAaqkzUzjFfmJLWNj1gImwNPt4r81e0+LtBhS0OjSlvmu5Oy7jcJ
yiuhAgb6WeJVNVa+d+AYrfDO+yxZCXNUBUZlcXMj6jaml8RpnZtkr7OHJwp5ZGeNqxfh1MyMPRjY
Wid+M9UeNxReuEKH+xhWnmgpkHPsWSkYvwVhisziuUQJ2wcY1bSJ4GwTi5m/jI/iTldar5w4Xpbf
6yUbjLCfp92hPkOmc8M7TDDzXsPLMJHC4PnSU/ByjEsyL0KUWTQqCtAvKODfFIFGLqo3BBaGmfgH
hafYV0m+1Gx4Cn7bP6Hpgu1wLA1kubYb71prCVQvlQGSIdlTEnsP8DJTwiGAi2M1NQdrGxIxilBQ
nhP4uXo3l1TRftc+ITE1G8D92Lw0jfn7VW6I2/xdn/m/pQ6jEaXtIufwaOOpXfmhY51P9kQvkCzs
mev+1T7poq0RbkGbmeHpItsNUTUOKtvSvBvRL6ruieJ1Vh85/cZR8R+S06RpBiI/KF9AvhocA2my
/FtdR5+lZa3Z/KefJqbaLunuO/0l8IJCygENOkWy4CNMElyD0mq7QPk5bjcqIot9oJa0EnucI+gg
6miO20IIQwAaP9brCjZinOCGH+iVfHQV0jjeQqqlZj/yjq3m43h3v4agOMzsgOoO4VwFdvZg1CxH
lXwaBFv+DMLLsAeR5NTUqhD3OnM8RTzpZ7OD+aFTITJnHTrx0auMYpugi/HpbP5aGBbXJshwEEiD
xzUuxWf5bpCiNo8TqIHSqcZUCn5ZczSOXh9AcU3EYA+gZEZ+LljDX0dLx4Dnop7/kvyVVmt3ZiaV
cag59Ty+JnjPDkbs0ImPOESjBv+GWXOs0JoqUgPQmYOkThQG4Ed2umjGY0v3mDbvJPqU1BNDSO4j
ihZD4AEQghMOyP+IF5rwuh2ycC52v6Vxqzg6Mvvsyax/RFi7xTIlQcam0g7Ux4Dd0a8sHSm1zoib
PDtoVr1+Nx3o7W0++uHbmmmPP207fZWLM+ju5yaDVVwYL1zStudXWDBQWuQNGp/Vju1HfoIv6BYm
kLY7iNzqUut0JeZ0OGf5bZJZ7Yf8ZKOphl4S0n7VuBoceyjuyKg6UKwZJdce59qDiq/wGizHNMCN
YPHRNTiu1fpRsfIWgYyZidHhWk3XaK1Z+tb/0udxxkflIxIRnDyWsU/0qQh950DbtevgPbnKQE+I
hhl7bnNrIf5jyf7WAAdy2XaeQYcKbe2ZK+3FpIGP1EpOnX49655aMsikl1ox9gZFeStWgron4Vu3
BURsWSGQMWuJPw7ZJGwhFYMnMdiiIlBqVAnro+uEgboQx1IEd/FmfsV9lr+J+WoYnRuaU/60lVOj
e0T++RuA4WT35kYG2RkRsljNGPltWhag55XZd2a0YtAboCL+TBsWr0uvU/hqsbpbF6RlThMYfJ0s
X5go293OY1R1c7fMOsWbaTot4hJ48LSGdFbffodUaygyEtHuj7J+Od2nSdW4qnyVVPu31EKr++qb
i1rRKbb4OOUtPO5XXS6gR+bAXKutZk7NqcEYOx9JKF6v4aFf3SpXbnr+tCF58x4i/lc/WfxeWUFo
L3E1hGRKX52FDUtuyWhBuNwOq1WbCvDGsWzmewfknJqbXMVSK2JGX0UK9pri77whDeLBDlVybPOh
RMJHEg4UeSUxL4jr0CyHHe5ULxb8hDpa9/AN4WW8zqxQ0sP2D5BywrRsT890psWJPiPgtYwoWc5s
HafZfJvAU/gXXVer94uaGpALkhrmPMb/TvrLhx+ggrIjCo3CicNcgeFY0+tbs7eHSHb9LSmUAbIu
8ls1/jSoF3n7VoBnNfwEWRWohS6XlPyOwsXhvGuqxCoWk6nq5b0XacKjUxOIpU0sprAnt3ePljC1
bcOTFcrlRI7o9dZtNczrLLmrBO0/713YJYJqwOD4x/UnmDGWVDE2inZ5+CwUoOUZJ4gmDm6JFj4j
u0kMFhVW84wfV3k+jAybYSB1xVF8oH9km1TN29QS9xhR0Ea14akJ6CZNZYwtjqDHuvIcc2OSHFmD
v3JYAJIDFQzQMr03yLqVZzwT2MZmEUGywecDGqYVsBN2rj4Uu2yb9ho8n1jjaqDaZe+H9hqncrhU
TEEf/+wzqD0WR+ehfQn6mjs1IeUVDyOGr5dFL8HuNP3h/UIxw+oOihLtGb1OKiPDlOH+GNttolSu
3zHFLwPCUjkLOPArief5E+lrcR8I/uF0VzGcmnkQsvL186JIMuM9R5hCjRYN0aRQbfpljgfN1EMh
5rR7wfDIDZPTVOel1tRYU1ahgt8SBfJVVHux2issWLTYM+cHzDQDOj4wq6FLjFHDuC07GKCtlIX1
stg2E3uCiv3+o/90uaFHUQtC99Cku65lvFHzzGMGHNnnbPe8VbgCBUWZYNxNWvfWcVrtdnGiPpv1
K8vCuw/0U+3MhTCZIH4hWlgkOw/IxKVhpT8ql8XjOzMMoRm/dSO02nK7SaKBxnYnymJr8sniRu6j
0/bKKr+y/OrWHOIYmgTFq5gNXqwjLPy5u5omCsikDtVKALnBCKxMusZqxAQ2fc3PzEeuDmckI0ND
QxVRrTAWB2q8dVXliCH+F7SXRgIdB4lq0b+AoYOPA+/hOKIKRaOyxLWUthqug5733R9xXy+8Cvux
jibbo5oZLD6w9EVpjmGkLwm/Lp2V+5kZenivBZeBzAGWqSVZoIRGky3euEpA/f62yuv1rYRAN+OY
SXNh1I9+tdAsZw5ZcOSzoiuSC81L/yNjn0zFzLabOF6nNP1UBEXZQRgmgIYgV5H3qyDp48pmhr8i
+GTC3TAyVZw6L0aJq6OeK7gWWn69NkoojBnkR0SPXUTHLdUxl0uD7kcwee+TJzdc0In/rwKb73mI
4Xsd/lK5iWemqx2NrH0VMYMq2fVerPfzGhcdvlCHidT/RV0lnjbAgm8NGmZBBW5V587qERq51pf/
FOkJfYmfI3tDGdBY/efzEPXB0YIpDmP0nLVyzLSgE1q8aU5R5NJR4lmH5tyaiEUKErfcOffandkt
K0BeIXBWodZlVlm+nlWMrYzXoFxxKQR/FqKzxxnNUpz+yKltbQQLy2SNldLcvBwRfG0/9rvqa7C8
xoESto3CgJb3LRCBy7nyv77GD4FI31g0IxWtB8m3D0ujyJWcVQ4dkRXM0g0ZtG8LLJzbYCvC3bpN
aKRv05WSBG1wcUMLUm8HymAP0N9xdzQ/XLLE+LReA37Ov3s9fUGSxDcsdoMxLG3qC3ggXfr8KvGT
KDsBIkJlU0ASSysPeL4kDdr22DDWUmGOuHI//Br0FySzhmLz0yOEtLVk/sfrLBOla6d7RZAaXjJ0
J/r2Mt5d7NbStAPCbxL9ZMbQMot21wWgvlbuL0G8VFpggAGZJWrpP/sXH1rBR45jiIntNZ8tbNYl
XjZeLfLxws2RcrKzf5H5tAikjAkWpmngqHe/M3n9KTnaL+pwjKJ8VaLLYYcG+HzaihlK77GIhRz/
gvpYgxXEPvjAO3WkRqD2SjKee1R9SFubhJvFH7LVABcq9RUf+TVFIfMkZ3cKCrpbyifNmNRJtI4N
e/boj+T1z7KO7YB+MpQbSBbu8FSkaJgLsaX3IOyAPn7WGG45KkSYNfGgosqIZTmC9NG0GKKEodKI
J3wMTzlgIhJHQ5J6powJDbIHBiBhL2XNJMnfF6OOoAOGeUgWkCe3uniKk9X/RvVgCY9Pqz8TXcFq
CfBtXmyqW4esjsQvkR5fWxuzoiAPCzjVgxcCvaebOThnzNaomhqej+6r4hWCnmXJEsaP+sntg36G
dy8ghDp7MwdEQCvk9wWlcVl/te+SmviTBHec9NlQJbXXk1+sUEc8K+wvDI656Do0T57o6/JUqDaO
dcEKlf7PJVYRZ23T5R7l4RKwUO3oSElLi8m+Dnfv0dzA9qaoZHQUnL74D165Gj67beNwm7ph5ngY
g23zgzXK3KlELFhEpZfNq4zzX8WYK/Fj4Y3yCoMWTtrCnS6XxJr8KVNud5Nj1CX5wY1aJrEIwYIM
Kwu5hD2FDiKdkglPsOqJq7dnVYiOU4CUmGzFImVui4T+OuuFIeOnm9Go1xoQ0slFVYa95uPxz/YN
XMhm0heQXckWBkTK7hccMJD/WNeZmIXdVovSe54toFuyNTe8mSAP2C1R3ojUy4lzC0BI0zyOCrK0
73AoCFXYIc1mhZe3Wk5nii4lQFT91Rp0X9LWA3z6S90OJ7o+KdFMbHWIXzUXNRO5KUhaT4V43f9g
tt975uo3P95ZZ5JjUOtWmuin98AaRYzd4iccXc6wuuPmeJekVz1Ol1NBn2LuGaueMGJFXPVxE9Yn
lUMz+uP3mKPgrxFus1SMlcxvPii2txF/RM2GKT1U8vY4b+mXrzmLFu7NfrSsqSZXF4has6j652r+
fKYPVJvU/UWjDdto2cwcSZ92Q5S2WmZm5kjMmXqpbAiV1vU3i6ZKWSCA/gQ0koN0JT8VjN0uV6Q6
c39bl0LmCs+/SmJ1LPF0uGRzN3yZrrs9QI4PHZ3YMfuszmCfts5Rovfjan6mf/01s2D61FqDKISD
2ORrelWo/m2Yi0UsAM2ituPcfHpvh7nxlxsSqJRa4j9oelyZnsGqqd8T6Vvei5hlMNRym5DMx+Jb
n0w+Kfg/hzh+CoH9wh0Mj+/JSvYugftnhPR9blUzkvZXf//yFQA6svdvB9ayV5wx7vOkvRo07glf
/espbVOLdfrjKJXAFYmO0lUr8VoNFM6d6pzzVKBLwDYAqZoVqQIE/XEuqqO98RNpthGAyHc065q4
JqS9wYdmEhCWgpx640mbIO0tPDItjFEnDXrMIaVD/bx6D2LyZLuDlB5f0q/e5J3VEUAN7dWS2kac
WDkExpa7kxyDYGex9YWe2fEl674GdXQU9hFTwkxyvgF2EabC+6RlSEZrSRjDMeqYQspqeRwP+OLL
ekEbbco/4X1/ob7Ma+S2STxC8MHsuiPVJNLdmkKEjfOVyXhf+6H0kSQZscp9YGPUYoZSX9F42xyr
GnOH9m5YyQknoYC1bqJNNOcz0Lh+H8QoClfVwQypWA595FJhEoAydwEsIiu6Wy7acfFlaFaezDTk
wlSqTZvCm11xrW3tbb3ZFFIir8NEuOAKI1wOeFaaj4/Zm7BG3z1oLICS/Ul25IXl3laY5lET7isp
m/oLrLSsqQl3LZCcoKgZno2rMVFHEkUNywvFHXSYCRcOOx3tRnH98EEBUeRaWya2mGsDxsaJLjnZ
tcYSNqqlDPvkVFh7Fq0n/oCAJygGIvbzHoAErfH1KsqvmeG+ud10uGpRDvUgV9s9x5/Y+nMhJzAo
PErE+7WpEaaTUfv1Rt655naPZZncciTEKjUTy7G7Um1XT0vE25Un3YnqkF6zyQYcQHpM6FZkIVEp
EcouMAMt4h3ZQYJopYmhzA03RbWPeLYB8MxnQUemmlfMhdyBkz9NqpXBfyH9srwbs3wPvvaPUrWe
670sMcbHuf4bR4IBcQdidbm7BnSp8Tiof2r7ZZdv4BKY5uR2r7z8028jOJ9ZI9yTToeEw7418P5X
6bM2NpbXuhxSDopExEH3bBjWOnWXOVTCcqxp8w6wWH+oe1OnslPxrU+3dGg1fsNuaYBRMMxwAKRL
dRwg5zUAD5s0VuyspDM5l1qtd0YrEsFos4TR8GFeJxfEKHHpNPsB6KB4I89vlayz7ieA6LZ0Imlv
LkBOk0AvYc+FlP/Mim1sfexG4Li3yl9/ZZMbnl/WcVmaOklCkEJa5qCjjPkrZ7dNevRsx9/74gd1
QHRGfecT0w7nneRgXPxRsC8zJnh0qvz9a63+ommokb2JmRH2iIi1bQy37xd7yGrzl1EvsiQ5RVfu
4VOyXzgkMCmQl7HYA36+SRxZyi9uAM8563I84/9oCGb8alrVAEmeVoucMzmVNC5xsy7JpFJ0L77R
qeqjmMoZopRJJQr7xE+az8m6yOOAoJ4RGCzRzgKgeEL+scLQv5LuqYVms2B2dR8X/KDjFaqsYXRt
2n9U2U8WdnsTgr8MPHHpxD9e7QwqY5plcWPPcIaN6Ixv2sgcrpWaxQAAdFb/GYTdY/IKdWNOMae1
6fCZHugSi5uNQgqFnSL7bdMUTWUzrNhTjYiznXwpzWG8EaNyEVXVeaIHQJyOJSETYXmg4S4IIaen
PIBoFJJeoOHGO7PFaAHtXkt2hcJlRlkTSy/gyWl4918y/Xy/utmwDE1og3wnpL37hXtfZHsZ17/P
31H76hsBoxUpxi3RFlAXEoch/bo6o1hBIx6BgdfwVF0txCqDeWvcS8VrEqqi6zySQyNWsWKtB8Oq
jhSv+s32JCrW6oLiqMeaNyg+jAC1YWxskcc/AXYTVNW3nRUjvDPofJB8xlJ9paAVcOBCxZPjdLpd
Hw8VWDbn/CiDmltCR9mlQ4xPKyI9paAsy2molKD3UAXE06l6JKkUU+9qytfOsk4i02lEs0L5vqBr
AyHlGEd7Lnfdwp16sTyYVJh/BunToDsYpcVLufvOsS1GI2zh2QZFWIdzHzVPBYpTXG5kX+76hJub
2SzHP/xOhYZ4K1zItZjVSx/X6JMwdowR6gpDZG2fpUcHDZsbNZVtVvoU2VIiOyC1LK6TgESL4RP5
LsITi8E3ZEHvsSlUhZlTXD/krztEr47TAE/zxLz/VFxc+YdklFenKCf2NbZ2TFMgJj/+eAR2AkMd
GJwLwIn+LuTsQFwNjFTeS1UAjDPiQlg1BnO8zxwvGwv0ckddkr/vB0kaBGGLVxl2wsKEUAWkyqFi
Ba5I/uNKHL4uWySqKcFzF8P/YoZbHFiZTefBhktAjZIN93V+u3eMR3I5T9C3mwY/vV+4zN+Ys+mv
/yTESEi5d9/rDDHAr9/Dijgkj/Pq4te+NSjP8CqBxfMdr0EAiw5mW9SXYIwDiufdf88gCWj4Hnqa
G1zY+uUvlzCqNSdcr/PUmy1CHmyrg77eboXEJzJkMLcMBKXvgWtXbUSqQZ77+vjK6cl5dv5mflkC
Ltp+wI7harCWN/6uCRH2X5LfaFGgtGSmZFnhEIvJkNjr0MVkn9+scuRvlK8wnzwqOZcwFpuxPPwt
Obq9VLEWVYgVC7UbBm3S4ZZmbIFKJQIknUI57yPLA7RdTX9SBKD985sgWsYSVPuR5OifYgqoUdiG
Zc1MvzxT3kYWWPIZKNjHAyWXVlVDVAqgJ7qGavcB6pMgTwTn8GUaUWm/+q1r0YzMrd841ERrj/82
49j3FSHUiDWYaneZhLKcTMdQRRyiQ/tqjyQ8QKxC+WE4xf68pXWcb/S5wgFPC4ToGw1waoNhgr4f
BZGOKO2jZC+PLqHwIijpj9/bTlHa9JJYHYar7Fr+fvSBq80Eg6WcDCwsxv7JStXo80Jn7GRs9INe
l4+hW/1xnbXMRYmOWRFrsf0r0Id6UUO+inpo9NvkNXMO42jvmo+YVqcTzpHfnQkSb1EE843hAryz
7S6gNP/P8rmSAPkoyZoeZ+1YQhAjH6qysT6jpYIztI7yRy3sfJUT2215yCdN2S/WI6/eQv5JnEXH
x8UWa5qWvz0RNTVwYEelOcIkl1xe8fqfbiubcS775B7Wqt9gxntWwx2gtc0Vv3ZEhCQHVQpkBBkc
Lyv1ylw4EIawg3hS9Sqj5S/ixMwa617fO730PyGF3NKFzXkpqG+ZVnuFUXDsO8ndPWaRx2N523i+
kqm7rBAhp+dg//E9Wha9vFdzQyP6ikBt+xNHdoJ7jm/0OZnQJPsQET228/vUSQYKt7RwfzskBegD
RTsuNVZkNMZ1mCwQd1B66rEStBUR7XF+0ITnWTk3Y4e56MKS/oAzSd88C0EKStuI3JwgfkFGq3UO
wgxbg+oFMIYyX+7uo/rwhzB6rkFgWuqcDkg+R/w2dedsFwifqZdJnxU5w+aY4feflV9iKZ+r7HVB
2yoEBJ3Bpa82n/b+ir+2sryY/nVRKnczM9GxxtH8QvMnJM29vxrJy4zaTCv71KRSb40VEAAL1rEt
0gjhwDQFeQpdN4EFRW6/EQcE3auKsbjUVkCn+LBZ6ffv5yolAwYQadj2Gd5u+18Pkhyzc2jetk+F
bDcoLNU8o+N/hnbwhPVYFnCYG66GKbSxRX/FF2AHxlVr5NysKUh99BS/5xdEcXKgqjj4ri/ycFyr
qnPdXFsEg0wHLVRH9z5StjCHb9Of0TLFoa/3G0LxrpM/8uAETAbie6obIIvQ0Zxo7NJIRb5TkeX+
sv7sNkVd23+Yztjox2IrlFjNNq6Ii3mhPNvQRltK3DU9rtfxvHCCFaynnb5g7M1M811OGXtFsUjL
ic8vuUhwuVLx8fIV46ru0c2XPWZHYyc0eaDHJtIrlg4hfcWYCL13ymp6U00BWMODrwjAhxHf2LGa
4kZrlxe5t2ufUDIOrUzRMgK9zNGcpzCq0NGrYT7wF/scGdOMmTWmRqwShs9lOzYFjnqaSv4yj9Cy
5nXignOJod/0ZumOM4wUjKjLE8uWqO1WJtWBRhHL1G3hBKuCyoxz5OrDQ4HjZuu1ZRYz+5S3WP6u
oBpmqpJN/mUGbhTeR3PDgp7aSbmZ/NpORg7kh78ydxTqV5zNKMquqeeQkZzTcXgzM0GUiixUV19L
n3bcfwrVy7vMcFMEntp8fpqNGTZFYuwhObHcJUxWePeatjCWJOtwaGDplnvf7UV08+DERmGBarc2
gVMah78rQNjg90PZ3kzTqm28MxAZRYSog758ELGn/1XcVcrEkMCJs1tTxa+hrhV0A0OX4R8FQ0hd
5UHLZ4pwffdtaYhEPJHy4V5K8SwHxHydc6SK7tWFlRke5BRuU2xSr2nD6NR1b1JtScH5JXMNXMJ3
N1ppo/5TKBWC4Zz8MDAzM53rrGoPO/VdahIZlBIBIcIWKXCXvUy3jOv5yMuaWupZsQik3g4B683O
eC4ZRU7CBdz0xje337gYiz9lpwoRC8El/qukh43mk1m83jzZQLRqqeGzsmXcXaPxvjcHZ/mfJ3F9
VTUSHmkkSZfGBQsHI70IHSv6TV22/ASW4E3Za7NnIIj4aY5u3NOBfug1vgMZ7vusBjEq0GTRtBrA
ej+ogPOepBCDsbBmwrznTcf2oGci1vVEKqJsFbsvN2rxel1hPoJNuuttVyNOKAhiTwma4m/amU9k
g/EIqq/c8nNLjEshCwt1n8AUcFI+PgVrOf0MBY/veRhbb3McW4pKY62hC1ZWrVPQ0xhuvjkgNypW
En/2RB+hBuNxKqiZ2LU0NvzGmweEYGmf7sf85suTD2QWZFeQWRorICNa3+J4qEzZKjv7NvWqDtIE
cLQI3nHaZJFJikiZA6HfSbLG5Wiqi6j6EHjrmhflt86q4dwDotvnDSAS+Ba/4VHMOnTQ8TZnuh6G
4ZPipp5DKNAOlmnEa9qUoDZRUyrNoEEfpFEKLhY+xfRZ2P65fddNYiCey5PdTnuEzHoUylb/KU8R
lJJITeK7aK5sMYmBuJtJTWDShJ5fx4Z/myEuqLVhI/Jcp/vhsW79yorOksf8Uq/dPpQX0telPGNS
iGY+3n2Fw/SE5Z9C0mcMYjHeDySy/XEJemfZC10n9u5pBdgTTYIOKwSVQotEBrawPz6bphNQR9Ky
nMmBbmOif+0kr8ADB3LQZxNbQKVtPGFAA+XVz4WHW7G2rZidokDRD2VKDhlKhQGe+I/U0RXBs+KL
5xqB48n1xP7OcD/9t9Fa030KuLMIpFggkmfPiiwaDo4EV3pNQlL03UjCItKPqpJ2Ip/dRg5mdohP
QZO3fjMKniaKSRRzrhYA+rn/RxoFQ0+jUrhM2BjbazQuAaIpX9MNJTM+FgzAc/1wuJDSYbHGWIzF
fpSWxapk9aLb5aNFCXn2nPlF/53bs41WbM1GIDMi7mvdMr0VOJgw0MK4pkbIENGwhnfvujD41nBH
8cC2NNp7k/O/fdRpxNSbwHccy8/2ZkixcbAB1lrVfEd+MhWEX9gkkohOyx8GohOxRuqvxVORcpvk
F+B71Otks1w4koDoFDcDpDrbSCkO3cMQRC6OyUplGNuUAQoQ8GN0ZLO/g/i9Nnj3AJYXZVF1eAkG
fTMEtX1ousrBuYktmgyWO0KYfTdAS3ODKG6zngy7/kuxUkn3TfEKywWOsPwTDjNByrdG/nQx+Tzu
RRVymk/LcmUv7HaT7uEddgGnVRdoPPgLzsrQ4RHpjTTpbJz+5xvCYHaX8CYT79JNSUAEI06ElV5B
p/gZ5Ks25Jg4OwfmJtbae1WQLgLRYctQ0+l+w+7nrtIFr0VPSQ18U4HYR1nQlzQRqERg7YXcCHub
V/pDukKCylO/4hcC8hRCOqSgfjxBWNU+L83mdddK6V1qBafW9LyyRGQcf+n0vWet1qQ32BNr+9yu
a6TvouUf8B5Arm2xkwpu6v9X81gkns9ydjI04+UML5m0Yy6z8GpTkZ6UuyxoR1zHIHxeGJIyiAAf
rn+/HaQ4oTsuEqd1pmTzuXhzT9LMd4sybMtGIlIZK8dkH9ULv3Fygt+KME16hLnQSs5P2Di34ivW
RY7BWDg7Zv3gKnYpYR5PfdBOFIL35J8TC9ba/GjNvVWbvMiXYvqHIqye2RPANsKLC3YWhSGMFdkQ
Udh/53b6Pb0vtEvOAqMB/mV9qi9Pf8f05ltuesky4GVMGaZjW8Cerl0qprnHCtqU4MmE1/CQe3a0
n++XCfPeyh34D0J7fXonH9PHaLatVqDFdPYVO/haaiZb5ma8WznKvP/l5QC2WFYUNmvORTZZ3m8/
zZch2ouuskQHXuqATyO0hacZgjgqpvqr1V+uAEZtUKFqmDT+HY4wXFGR/gzVXN1JzNqzaGDCqSpS
qxwmjRM3jfHFVklLjYk1WGqw2CAcelvCwTQojpR2aPnNYYXtw1OHmJ13ng7OmpfjeiB7vb073Dzt
poGsYZmiZPj4BgXp6+dCBDkPaSNANqslghRsAXqsX6CQ9nzsHJSV+bUrXCQ5ujSPYHbRHUVsx9us
re3ZJOib8ZbYu7RPBARqR0rQxg4V9cvJlylbRNbNjZzYgYVDoW87Zx3Z9ItlbguaynFOBl6YkWUx
GBCu2hxr04uJc/XyEyMc+G8g48oOmhdFy7gpVZBWwlNMwlUXhjrEBrdCRAVkRS1PYghahsjzrTqN
p2U8DmNWdfJPdTHbvx4CYE4X7h3m75D4qbavuwNzkqzAXE/4RVDzRfAmrJPZi5rrZ4oXifln2sQx
RC+CKS63vzKcX8x/ToMCCl+xySxKCQtvBxwoEmLEtcKx50+VT0FnB+K+PG5V3uOMld+G0xRpxFYd
qM/nMjo7KPrFRlq+nF8Va6d7LUfh2ERTftn6zbVepW9l/XZe5Llg6rbZOyO/duFlYDE/2jgC1OA0
B9d5DKFw96dloM0F93+wArmQ07mnuH1j7QU+naDRXoLaD+Dd0O99oPqQCluyLzwnVF2YHIeww78d
GTmHCx02i7NAuApek3WL9HShvNzMcdR7e1obH3yNk9aGtih+Y5P7PXnT1h9/X96HByHcyKgKLwVQ
FdDodYOsIEfoWo2dOzq61ezIgWgG+AaiTNbiC2VrUVN0N0E8Ic+4i6Vl/WSgyulP2QER8hYs3Fi7
QylMXxZacwE0bWhx+NW6KsD1f3YwZ3dQjCFmFwBLd1IF0/0atMJy8qPzd8Q1peXBcfB7PvruQJlD
jPGKq+wrK+g6Ie3EYYWyTbI1uCBYUGiGx4SLqXISbaezDD4szP4c580TBfDr2vw3ZUgvjZALLymS
CC5j5Jjn/55KKTdT+tib/b/dtbEMBnJYDIquOzZOSSyxj7IWc11SNTcXz54boCe0UXr2dH3NqoyV
PB6MFuA89WzhRY5dYgBfjpeClnNuioLQIiNGpeIs1r21v20kOQ4Uy8Z7dPn36+VdKlEM5KcZXnDP
ciQeulsUC0Og6JJLTf71HvUwpU0a2PO/3c8NYmg2aCVsdyI0KcGGZdghsiCcQL9a7VsqF+gD0Nqa
WsOKQRe69nszr+qQ72ahueR5vBecB9T7XrDalN4MCox/4SlYw8V6V4MjZXRUmMnVsEHhsnH810i8
k/ncIpcsYi2a1sbQLNmYM+scADJQm5QxyHUsp4bxvkAseusxLdVDrVieAbD5nIOa2knMfRX7RpdZ
4FMrxcfhr+r8HukLCGHV81OnxqPnTPkFqzl9wnMIEx1DJN0VvkWffkKObUi3GUzM+2TMvRi+Eu8b
Y8VltxDPCivu7eb1kziK0+ENR03hazxsXlcfn3KtLDSoz/n/y0UrPTDMRaZkx81rQAlUV4IQyFf1
dY11tUbsOGVMxNVZs4P+4aqv2SBmpVnDjU6KJLxbk1In/nOh0CO4+qfyEEEHeNcHZYvdM8+/kWII
rp6oZITweFztwa1jb3Q1L58csZ3uA1V/cDrM+GYN2j8PUh7oSkIoAZFXt12GYLzSK2Sgo029dc2t
ZuDOCYPnKg1f91e39jYChk0HE+5tq9pEkZPOthL2NdyZ+ruS0Jeo0YN03m7ZfUxVXrLTY+M76Att
EfPyqYS2sk6l4NdIc5XLRMREHihKmsDiz4OT1SGs1uvUBZaQBfN33xDY86a4tAgERQGyvNyNdBnW
erU3RWEecsOOPcFvKa6wd5rMi8qVH7+fturcSvkh282+7z2xSiYG+yBcoL3S4cmaZbYGeNUgCutu
GPX8ZlNzDPphM4BYNhdS3ZPWcD4eqTEngPGA3RQx4lxuXCrxCQ+ILCkvAN5a7ChydhZ4MOyAKWQA
HiyZSRnquftBRxz4FFucRU0DHmeSpb/6thHPeW13vZKnHJ+t4J9BvFXqDhgV8krhTLylg6wCMKKI
lFYiDNHrz74x9BUtc3sm3aPy7ALwZcVHqYm8slde0lz5ezv7T607KBx1Yso+pD1yD60F9mghGEjw
KqstzLwiJejZ5UHJb1qmnluHBDZbPVqCpoLbLx+afc7KtwpOwDRi+qtmXiOiFYo3E33X0sYlgXel
U4y5wkddol7NtwwVIoUG6tVb6/8bm1zARfnHSTixhrLL7QHUFe6FAjHGpoMetBBZhqgDd3nNcUsS
K8cOl+nlPLncPqlvyjuESAzlW7M+yK8PnkkvBRSTT2yQccicDztO9RQFy/MfVoy1xxelsM0huiXx
j2xrOzmqMoLg7cEUkAyiQmhe3XhkMKuUnb4HjUK9X6dQnMh9ZRuey1Nxhi8yPdVGnQhMNET/gIe7
8ABeOcJcDvqWvbwT59s6yzWblzfUYpa3wLrHw8bvvbcrKsHOl3SbNmzmvWUU3uXPxb0M2+TgBs22
2/ZLYlzo8BmR54esA34ObAAWgtqZLQG53QTbOkGOBVQquAxnwl6CFH5WAFAUYrlpPcKlqlOWnvPw
L2ZzPzUW60SXp6THMYHB79zl4exyilCnkhX42NH3XsrqGEm8CoWGILkSx7BSUayKxfab4sb1Lvc5
b8dRp51sj7dQAgKqtfDQ4I0QRiQq3lD7qUDntIP9kI76a89RrQ3KENfODNp0GEbAWoWt+4mGIMLW
62IsvUCZ+Z9vfqC3435N2jt8P5/QXXqhQOr+jC2f/gFw04V2ThkCGUmrLPQxBs8cBr7JAUHfPfDb
iztaOk6VtdbxAOfEmr7BKmU2LuhxQCpipvNCMjc9GMvh+JwmAHU1nnvHqkmCH20qagwBCfc1w1yg
KZ5C3cm/13NzLx4qDhk6jyucwtgBzg5EMsMT3BI8z1Eh6odIn6E78o+CCr/fNMEcNJdoL9ET+THy
07eEmy68DUR7nLQTImJiLFmwDpnlU7rPZeCSWj8SRrx47q/P8HtEDO3mdDO7vBT2M2PCPPnRTJOT
kL4xMUw+1PY0DSHNyrVebIBCf1yBP274Dux5hmaVoLHM9BZPnMt5ffv3mP25Zmr725dBviuubbDP
7q1xYjTqyAcOGa7HbUqmqq9sSr28Zkc+SFhpf0JpapmiCFST5qnG+au7mWwwPyccqMzM5Yz+g6/o
Hpdm7+VhcWWVde6U0sAjAKR2aWCapr8GFHQkgsJlzj5ENgnmvr6DyOkaQdZxaJRoV5Ux2vbHECSE
UkCoOvn1JMkGOG8Mji64ASg0QNVIGyGBbpCjatE8WxhVD/5liMC6Hh+mL0y6aU76sv20OfafdQx1
3KKssBL7plFp2oeQYuAp93/7aJ8VmCdfx0MRRs3oGTp5reng8noD6fnVF4Dt7OGBtomty6f/6CK+
dPl4n4X85npWD8RpJbruNsJcrvC7s3ZRdvwKeBW1kG80kohMYwcQ3EDtWpQfdABCNLCmARf+DLaP
cHZin8M6HgOIMWCJKZ0Z2VKQrlWcN7kjKhSNL/kXVrzer4467nwOHMEaUm8L1EkOuTi2TczpWPOK
M3YIv6S7EDeQCZ8u9OKqMmHuMNFo9OpeZFw4Ueg9ZA8QkNJyCiaPZDl5Z+IAunKE0c1iis3WNxW+
7FsjFG2ZMyfSppPOvwSQu51nRgr76GNy5OR8MKm4RHScVctMdO8ejGfJIubmXMJAMTc+eSVWPrAp
UDxQN+2BBqZo7gxp+K6Bx4cetYDrcSv7Qk6BQpQUjakaxwAL0E/xWpKKaZZtY0Wfpk1wBC4PZNzT
OMGrZEctMgVrWb1qsaMyYUzbhN1vWgZCCq0AjP/Y7ZW+9WWpVql45pZ65f7x/+omAzW5cJjhY88S
q6g0prsjXE5AeO8Xy8uA346m+Etm2Zo1Lcdvl6+IeZW6S6wARzcbCMQUYqFhYy5u/7a70zfveIzv
04kV4fK9zeaeAdgHCdRVHNJZpot1D+6N9FEQOhAoJktazar2xvbPndm7cNsDcyRbAXIenrLcUpHy
iJZGwXANZY7fpzoA133ktQa3o12fgwaTzJz3MusAtM1ZtJbQQ7sxF9XpEbndsmChOhdlsT8hHoKP
Yp6qkGIW/PQ7uMb38mifrIu2yUj9kQHtrFkCFVgUAmfTBkqlo4twABLhlv6d+W1E4wEwHSt2jaUw
PI3Vvjewla0kFQL/ArgQWByx/SlYxyidlQ58EaGMVt6Vc1dhlZYIv93A+fhPiUBHUGSuGBCOPq3Y
fET1f97unngGAo4m+OOr4dC1lJYVpO2szp+Nbj/3PH160vmRvcnsy/LHsVxBoXNpi0wCkNgk6zF3
Jlac33ZdOq+BJ1QgZamQxNkNbJ2/Muq3CooUn6LSIa34tHSMNwaLp9mwwHq6hWD8V1gh8mLXMWKC
43e6Lz+thasJzQI72Ydv8UJQbovVuwmgQ2Dbcc8A0jqtVmP1MBm4hF1mMVtvfom7zYREevAjD/IU
Q/rEBaLF9KlZlzsqlRbXeK+cshuse7nC4oRrEIsSDpk5pYpnPZCkTI56QBgSgRGe1ua1YvI579EU
2tpAdXFhTi3AFM4Jj2zviQLn5Y0xnh/a7G3zy77DknWtg2gHMuwpCeskZEHMr4ITxCFz8EjLYTjS
K2CsPe51ARfHS8xLKhyKIk5bSW/rinuoV6zWBnv68WutixMjbRx1zIhnpEkrbvFQc/uTtoYdwks4
/BKX3+YKtj5/DiBw1NasfWUYMHbAxZd6lCf4za9QPvL0jkoiGKVQ4QeiGwNzoZctCcEr92FCWEcV
9NrKFqdWhkTLDUqoyJIqrVd7BwhMiOD8dAaAX4gaxfcuduZKkDpTIbZWujVyjjo+A5X5sCE16kjn
DbX3NJFsKGUN4uhDIqvA6whLU+wThpoHIzijBntbzADgys2EjpHhdN2HvFIOrMdbk4YLJ9MTN13I
lvQxXEj5UdbBGkdrvAv9C+dy47BqyZ3+6qQtLGpycIzW1BFfT8A9M9KY0Oaj/jciiBN0W4bdsVOa
3nPc5qmBvpLBMLHCIDswMwWDo2JtYDfIR8TvHAdvq8OejECbtdQ26haOX+DWvDq5PXTAPGQK4KaK
LhVxNmFMtLCNXR19FnF7kyHQPEKks5+1bZo1PiFuk33CToJL3XfnJrOKvN0W4ni70hY3GmcV5o0Y
D14XZf/l7xNT5sHMhZN4vZxOd9YJi0IRN9oFRc63sLFg43+zD1PbOjh/t4WokvHwmmK+ZiVVXNDK
wiFh0xS+j9A+gmwEMIIAAY7YDpsfP4sv0SsepS5F7bf1Q32HBwplrmhfJgmtB8QR/5UZnMEQOtMp
3dHh7ey8jN5Sw0oeWaOId2RD60dKEP5YGABrRTovLNG5LGBvHmzr5n9akywpEoJyOTapxfvV7cP2
l5QAh8C/JyhW8adZJJGtx4Z++ffQcOFHtQcaphMfPaVnG7bCTY/0pmxayaxrQTU9bQLRLXzmPboE
xM9xbIDuWmNfzm7ho9VjeYWpXcfwKwV0ABQ+TDpRIvX84+KyPCUWwHux4nZqMTSeL1evyqm9ebRN
gnGcJ0A4RN2XsaU0T5TtEZ4e/bBDllszTTK5gCaztx8oO18gPpSRp+0VzgpiOVc4StHH/lV4ZwyC
Ri4DqEDmt9YG6wDb17tUkpn3w2X7TIeeTF+Ln6UjBeEherWmV/iXBidghWj6J37skZpc8i270vsF
kh6zLttriXApo6uVqJZkyVx2T8qPW4NjoFfG767NXQuvKtBpeG4pXoGnSyxPTWbU77hhDqKi/VZG
YgdXXQNJBb32jyKguRSsk+GFaE9EfPr0zUJuV5TJUF1oxy+f/cipTX7qv+kOUvKde0Eod11884Rd
d2Px6PvLZGhwhC7kYnZ5I/MIICO079lVJfej7IARoOFBvW7UmqH2vBAzkHRQUg5J0mqH7SzcgJh1
pJnnhoq4PO9wJiKu/GTbGn05i5rpUiPE2dHo8GY5Bxjm2nfBrqp0gO1+onIz6GDug/HzoKvjCb5n
dE/ska7sWGOME5zBjphKqlCzXhNT6002nZJKVJjz/fSNH0uXuisBE9EUqBJMWQF6h5OO0a9V6SNx
mAcgPWVCEc+dbXZ2hk51ZjcgAU+a2UcXvW34Htt1ul+/45qjbDcEUVb7EqlSUDPz1QGNgGUiyd9Q
yjFbXCK8R2XhKo4sTBuJfEjSiQLvtB9s/EGHX/NBpRs22WKeGrPrzycospS0bWlE8LI+XKeCwkNl
5+FyK0VaEnYfA4/xbbPtLUi138RglzblWGbhm0sNpGHwpbG8+4/P5q3svHfk17EhtWuMmJwihpSA
USR0ahat6yzvN1gR1BCXD967s3Hr0KizYMTwaoUdi2omltovnunwP52iBKA/S58DE8VV1vJoXMyQ
UlHoK7Gn8yMRtdtF5Pw/yprAe78JSkXJ8anptedMGVdQJ1My3oejTJCNBlgb954l42JncIkMXv/C
9Tu8d0VRHMM69jkX9DqtmuR1DiFWewsj+efjffyIS9PB1EYwJLyAMWhLlpRw6g7k2EfXBWZscw4c
2Qjc87DzyXvh8bf5Bto3TFxW5MLGLQHZ3VWOSHRKQm8FE4biUSH1oQddzhA+rHLj1IZXnHl9yEF3
GoIRJ/DXJvEvc4YG7l+iEfh/ddefuxcMZ4fiebFS+cFPq3ZPEA24G4ized2yX3t1ZoAuIrQzOtpG
Bp+/KxIUIJO21/lAnlFa85Cgrs65zEtw4yw771Hx3BPtAk3h/HMmvqbaPRBueHVBRoibbTW3rnTe
Sy4O2xEjG+atRIuaKkdu0Wp9fx/MCjRYTQKsV5vc5l0JSk6Q7LLLiFtLfQlFZXb5uHJQ3IxhBCIt
mNa3mReNYyaSTs2IvMBI7wpZIbZ7xN06AX2kNQ9daS3eCryq+JtmxkPkGGf1FqQn+2LQHrlPfnnP
XEV2bzH7AlGZRDjDeXSPeuiTv93ynyvcIan6Gsv1qqWPmExeqbEuO0srOiwQSxxtJzoruKgHncrQ
P9RrRQ6oDd1OcMTH50yONPTfjgkcyLLmIU9nWy9V7Tk9tRyJVcfPo6LAl6sX39SqeK1O6/w3B8IL
KrIOclDLz9VMINCuKl8O72+CviuBFNhTKNR4bO78wmhEnqdoxo6MhmQXbgsOlT5oF665zC6dFg28
IAXL9D7fJ0JF2v0zZ/4fiefhYO04yIvR3wxXMipzdjnbGTzUnAWhXLqv6/UvPnnJJUPbMnpQICi0
+BDRKVeyBdhsWwXa2M0b/BZv78u8vnoheakluL5R8ttc0U4Nvb5Ste8iziDIeW3OG9CTOL6GjzX8
i+0PtV5Q7pyyjGI9l+Hy6uh/elES2YfCyYSFLgj9XNjWT6Is/ANkaiZxu/Tq/J+a5imoJfEVycoy
qv6gZZ12138Ea5spnDMPiniPBKyjToGeWlEAq7OPMjSq8QDhdsPHxVWqGzWtCIXUzEkNnom/r5nF
4De9PiJi+/S8JswSgnHKWYHmX3aU1OoFRBJVlM1L6GxCdIbcf+uOgyM6vc0TqqrvBsLwpxX71ori
a02AjHQx6c6WOwce63Yp+99RXZeru9+KwgdTZOibRzrZaGr7r/SZ/azmj+O2X9Hic1TgqILrW6cQ
mmozqoqpX2gOaTo2Ga1T1rF3g6TUKyuPP2+iZm2J+n4wJocJJN0JkEzuHHxp+xlZOKZkqSUM9+YR
poFrYYCnGvOdkLFSr79CFbm6OeqkEUR11NIfikjfSii4EVPQk1y4RixE8gVEF4p4mP2zLfVf6Clv
BIteov4evbzeod6HlVhpAyxKO26lxNleaJy16+4nAqsl7dfhvNVgFTem4DOUrlNmQ/IjC5/2or/x
U5hw6dAW5n/nGBpOkg9Om1wnRawNdSygB0nxLALFZY9IhoP/oVpFd4t0vtlAawTBrVsnHTaQvNNk
x3Sc7jrEpeifFVKAruPXf8DKXUM0dtQaw4whoY3QyePdqGJkUWrwEiKalAoVzw3WjvEG8Tb47fgV
oLSQOy5HmKlIFu6/3qZixc3Vs/eOK0s5kPbeFF5+b8N9XDyNuZAeIOYFruh+hbs+EyP10fv0EefG
FuhQgO9VNm/iCCthyYzNltzqtFFB6mnFQ96HNv1P7KnuMQ0AkGTUx1692pEC3ICHjFja+6HwGPUf
PnqnEpvMyjHO9DpYIWz7JMiFAxbUD2G074/LW748B5cxCz6YSFxyvKsRqP/aiXZAVdIbA9c7HGKG
Xo+jd/wPCJAnYbIfo96j33TFZQQqILLXszPb2CqV1d3NKuL9aL6622v9spwM2UKrqhd09hbQvn1F
LHprtTRvh6MVUeyZ2zL3NbQL4bWPDPD7GXWOdwpkaaBdYha1Fzs3vKY5kuMPX7qK1kVvNVORD7ZL
V8Py5yiXp2JE5ouo7dY57TOloV7pQQNoeaAsET01tTeWCDg3sSgOY81ovpbZyk07IFYSvi48kwOS
0Pe2DxCCBkOVV2QwaX16MU9O7V2VEdZvjmqbV2EVmAitBSm0nbSXKE6DXu1vxYRN2Og/m1a4YaYl
7magjS+znrFlamyLDdOgMzYKryvvGfx/0/oguQSxIODtwBA4mVBF9fu9/TLqpsG2KgYggDO6a0ku
a92tsJaN+NGHKDDZLJmyvfYq0nfnvhRLn1qX3b2Ixgo1SMLVSPE4tFF8y7eYYD4xW1LxGhSc/2TU
9ZZdDX5dJzBX6dzVULnUj0nrpqiGJpjdL604e5Gy5WbGUYK+KnhpWS9Y3E+LbHmMi6au2KFWBXOI
Ii2+KewNTHDWtLXLdzmZeWMLtu6jAgJszh/nY3/D9UY8EqIFtUcFkT2ZxDfSCTIKJjnFEMjNyN0l
C/4iZhg/o0XATIeHZMx77n4G0lRVgLG3Iqrz6qSeRm8v5KUGNAOTfCklL82RJFb51+V/02ybEBaV
dvPKRVArM9h0st9SYpvot3+5uQNJZ3nhSt8hvwjYISHNEhO760UvUz4KVRVnhmKyxYJe+eaiTNFV
Uk/zaCpfElHo9nFDWB2j39Uk9XzXXjOuJmel3/zZtjatwzK4yYyzhm7oygIecL5tk5eGliBESJcJ
HxFb129MGsTBZZqdukyvKaJbvqI5VZSNMqwqhul7tcv06QRw/ZMirX/hgi2Tz+HKg722ygvt7kqd
i8m/wHrmfTMZGkg/fMYvvJUSw5wP8FUn0faNuaxdGSXyiJxxvTNqLXaEc1bNDY7s29r+Jjt3CiMS
HKy/WJCaUed85H1klsvNzev2VYxJFa7JUcEGLVzOxZHitjygbISOJ2DAN2SBSN/ZCUaJHhZsVW32
RC467Di8yyg9+BXG6ACKs1HWbHL+bbBMDR868SE8AAYdsbU55wuJQ+Zdc9i/qvAf5lO/VkbQBRTc
Y7ZLXLlpwB/EXOU2CtMzFueJWSG9xOZE1/2rwywwR2DnoBUuOSLgTHZk7YgZhc3uoJTm04HsUkar
Xz3yFaPxR3c0CeFy5+jbliRXuwnM5KOBBgsDbbSpJ5n46jtKGabXkleg4Hf7HKyK+JTy7lVxo2ZX
MuzSnJVDrFwkcNdylC+fctnnNB79njgtj+42SbPOmOtM3TE8h9T0hW7pR4RD7gluaQLHpbxOgyey
jNb9/8f7uHbk0Uf8yyt1asn2XAPVFfKQA9Te1ayUATizUHUnIWR7RTD4yIOdCjtelGzXL5dObXr1
bXKfnbNkuYGW/ggrkXSnfJ8M9xM1pp2TzCwg8/Ht4w3Q6OUij544Tj2AL6TeEr4LLIMQfJgN+pwp
NUEQajCOrdL3njubPjtjMq4AW1+4DfA79AHoG9u55dUy8M3QxBiUkHVq6slq9IgWXm4wwJhSK9t/
0v+qkizF7jgDTHfOcqKf6VLFJzD24lXRyY48Rttid0abZC7WAKwkjC4HJh6OoY3larnCQwdP9ik3
81OqeuruHz9mkxGlvKATWVZb6Ven6sZCutRQ4ubCe6wc2i1qdpmlWGsGOiCuRdHhRwCY4OS7tV/h
i1Oml11kUqb27GHXpA2FUGZ6g2KRK4lY0N4BLyh7lo4RA34wj4FJM7MvnMO0IGfHWrEA0/Zt7lpR
XmtAefDNFND9rAy6RXQ44Jxani6BpXetrecWROanzoWSvcfMrhsBeunP7L6UixbSFFmp6/iOm2W1
80o2yqqz60AauA4Ezdlo6Dmy2fnp0Sj8LM3WRhISdoKoqJt/DEdG5TCa9CUbjPVoH5axY6bDeqpG
MFtRy8ki9Igjd67t6tGcjfZR4ftwVCi39tO8pH04zEYX+mR9XaLdFDd3mxTh8LjvpI2XBa4dw8RC
AVxg7RVJhJdvhbpYMFIZmtQsxyFzYPD2PAt6IOjIi6aUHV7Rk2WK93FUBWDmBRI61yHMLJugOj/4
rNsCS3gCatntz4NixsKMl0kQWV8HtnLsLWpgQyqi8i9PDoTFiq3Lpz+3oxLfTNuwf8b6uABTvHnS
V406o2OPHIV7C/4OSv8t/wDre2f2NappFK8MVzUJ2Ck15D9uTIQ+vDo+KURLkv1tY2diuF4OHYfh
ZjXolez9JjzzkX4kk6kYJn+yrfOVDtNP+ODn9Q4F2CUcwoWktHJPZLGL+ZWE1RZSQFAxnSXY3QhF
HOj8n6cc/pNh28xVpl98Riw4gcpt3UkIX7pN0aB5fT2JpS238gTNLD5cwrWtkFbfMP8R3OU4MaYa
6Vq06hKjQDM7mlpvRP0nPuILjIPKVXbL5qepcnNfmFAjhJuGUpMVWnSjaJRPuytJeGiZQnVXhz5G
VI95r07sTV0KW8X3r8/Ep0We7XAuagHVZU5KX8Ncyd9XBGKu1OL0WnDGwKXkFaAsrTyoy0iXqYdg
zXnkJ2/3k34jPQiERi6twR6ISLJTnJWJq1FziFKhhPM1DzHGPLWzzagsXw75ucgVS8C2t+pGLNWx
0+4pJJbnjeuJrp7WWvjl06cxmAQR+36DSG71I/UiVZnfwzdtv58w1ziYRnOnKs6gxqY3Dd2pdL55
dtugp5AEIAzGX4OOH3/1eZwByRwqpoGTe0yEyoZgwuPHXbZDeG3AzKfidI7GqFILAwVTu6e/0DBp
IBebdYKOc8i4QsamKd9rp+zwtrBvhJ3IqyrCSGYCIyeIwBH/WUxZ+cs3UcxDeI+NSViWtrLKMpHj
s52RKah0lFQ97/psCKCr1Ns4xWOs4EDMsgQgy4QSKppZADOVQgDfPX6g1vJzPkK61k9nQDbNyTW4
EvujFpVPUYvney7UZNdRyC98HusIgMfF1WupdgzSwRDkxEQ6w2KHHD7gvLbvXiQLPHBXyvyfFgS1
QZ+T0te1pS8N3qvqBrjX+f5u1s05Y70qIFzwl98VOP60cdDd/ZKNxQDnxWr6GDMFWShnHOiBUX50
RYHHFbELmmk4HkbGlFZXsxTXce7ZtRiiN+NQkrQnFBZfGSsumDrgci/WS7lMWyFGYCxzECGmyPpY
IngfkvUeoOqzah7V+RPJFys4LhokIi3c5pXKQVkK2n+7hiVydJfmY2xBmvFqpDmvZewKGXr8Gx/U
PyAFi/lf1ClAwCmr3DLrTV1V0ejZ7s36uNSoCPX0rTe20DINhz3eCG+uDbYPFZFYkFga8dWG/cdv
fwgWToJ4D04T0Or3+SGis7nyU27Yfi6I3Rwx9wgqkWGury4dtVGdHYDTl2tBDcvxSXZN8mm095hM
LlIrYutXJfInaOGBD1QWhAylzVaJkKCZNs7l9AHvU89um5rnKOSgGfybuy6SLcYtrfP7qIZ0R0W+
Q+k8XdaVTH2v3+5in53sYjbwhHJrRREypKKd0auqfCa5EaJea42Up2Ks2PqbgKy1VnttrjNDSSWQ
RDVOPfZzr93ythKilshhhXipARmNzwIw/y9m91VdF5v9JXSq0MzA55fQJkXy2X3kyAXd0YKewjrQ
eiFJvKeZ0hH5irOQXj187scz3Ctq1n4IxJW/SHlH1yL3lOp73DFy3vf69yXd/oVHksCuTVVBw5/s
krse1l+QM4ePcKO+QoY3YLpDOo3wsenm5Utp/eZgoWxswRWsa6KR3XTTEe1jAnX5laDkbkU2BiGy
/ww++GszJnyKBxuLIPeL+LfEB7LvMm41zudJO5oj6EvchhOHcxmXmfjY9Iih37wpe/MUwg6E4AAQ
cvlGRynHxmWN4JgsDajrxNJvjVspp6qkE6SlZuh/D14HD/bdGzdt5fev7vMbMj4xAVNifkbk3mgD
IvyadcLyDTasqLY97XBy+GIB5St66a94vWn83Sk3x4G9Vt7pPIoV5AetqMiu9hD+69iyrdnwI64F
T8OxLxXzEdXQi8kndASs6zG4lsNWOKy7E7ldqlNRK8cUmb8uv12BIIa3g2FZRhs4CBS0IWR0tnv8
Y3lqNOj1IdhHnYPr5xlqOhHAHUBBHXQLmeV8cag+itynKBGN1tLYGd3iiM2caGLlpVq/nPOI1jme
z8Ny7zP0aMPQsNir3uw0hbI2xcrJAxc9VU7iivSb9nAfDeoRNm2VdgdErCVa/Cv3yMrCzgZ5xsra
I2DvOnFCz3KXzrc8Plg0PUC9r/7Jj6/rtTRB5GEBNegkjc4b0RQMBB+n50f87y48mkWRt93BC2+Z
1aZNQBlQ5m2CtKlX5gTFQ0ED6h6qWY0xUOIKh96z/+3FD8XihcvDb337nzG4kVzuP0pCfmwkDuSp
CkbMwoUMKFrW43iWMj+GwO/mq5qRYk5w32JeKoWnkCc2yZ7NpR4gd6Mrj/9fW2jULv2DKicAEuuu
2MEx8Hby2/Is2ZtnvhwaGn4R49uir9AnMDPCJAyQMHC2lMIz0F9z/H1RiDZEJyoGOzjSwhHAd8ty
qPVZmKXJtmb/I3xYxkrE/f4a98QIKkhPLeWXw1ksWYeoHj5Ke/I/Ki1FM8LWc/Wyn7V2VGH6crdu
PIWbye0p9aVDRwfT0JbZgQarfJQOuDsefDkowvBvFF8vPvf16CQiw6VW8W1xUlSFYNjwHW3y2B3e
YIdSPHogkYQIvn3/fpd9r+/XM+haOFaJwkpMXx5aOSdCz7XrAIr+Ykel55q6EGtX85Tm2SFPdqhA
DkXtJVORNJV8/kdpuH1D2k6g7QooAsyd6xSCFr5mMrxyz0trwZI/+gU93+eC/+qt5XGT9nh+l6oK
o5aYj8I11sTqrbOXUESv+F7i9KK1TiXWJZopr7uDd8yKBbLn5yzSti1pasgPuDEIvCxoUB1IpyCr
Q6qfpW4V+dtrHfUWXG1N+ZD6ZAW5jZb+JHWTXO8q79Y9fUfB/OR7YBUbv5U7WV8Ko97C/I7aeRN3
k02QJFawGwZRkTHXMQ8KAOj+p3ASHfYHYbZEn2d/Xg3tIJ6is4tGzynU1lnKWPcpHeRglqb1EaRz
c+lpj7TIrOiEqfj0VthwR8wlFA4vBHzMKywCFckdKUlA3f3mgrA0nXFP1l4GC5c89p4Xg6/4jmbi
dEc533dIMlBMnjfeS+L5R9V1WgWXZCABA26GLUGbYGCzMAHTpEWfTDDpxQrzHOn6GxkdvWCABnwE
w+oueWSGG6L9yqwi6/WF7uzs//+q+mj9a9aYcUEPbNJfBpjfkQKbxNgWqGvmwIq2zK71e3O6SukC
btmGQxCvUEz3ifEUGpjd4HBI5UR+u40q6VTyZbgpLdTwgzW7Zas5l6T2Qr3pIzzI8LwPX1H+A3gO
eK0Y2y0ys51MuKIS/V3X0jq4g+WDx6RzhAueA+mWKQrx+4TIVx+UsU29p/z2rSGXycSiQqEKeFZR
aGjhHvx2pyg71xfkL1bYib3Np1Q17pGBet7zZtz7YvGb81OTNeaHw63P/LJGyjTwzPEIjr6U7Rx3
JvegTvt+mcBxTjO8Mzmol+hX6oDM8b3NeIoZQbUtav7qXeR9zqJmbm1qqSAqP5/rGiF5n+BP1+KB
mY0fRGlj7wgpPDaAYXcRv4lUtRAgN7r0MW69DXbc78aJg6K2/cpIkxIa9ekz517rK9O455v4FMRy
UzBbuzPqlPXjHmKccgjAXyHUBpnXXC0SpDBn0s7BQzxbGF+D2Ta5ZGmFpi31lyNDTdAKzSVTh4U3
ge8o4lR0NvOrctq01qSHfCL87VQulMAUHsi+4zYjRcj6Ieg23OI4FLC50xkQKguIBDb98a8R4exy
40eacDpoZqYq/DDDWD6maZDVZ2nOr166uUxBj/vnUbyXwAA/UlO6y8SnJxcTQM05P3XjOkYVFEC/
dsSNum6ugNSAkQw90cnO9WpLtM+UNHZFCxaZa+HBFBBNSfiVYn4osFVzwH78SVTHpSAKijH9jKjg
W14I8Csq3CzQ7di2N1KlK2lewSBbg8FLOedfM5QOfFiL9ndxuN2RS85ZCcW5cc95rpIzbYrBXOaV
5N6uLj6oCnEwi2ZoFWdAZVX9DppPxBQcPbc8pDjunYXbq4WZty2BDqH0wC8R6CpApwx559yqzGy8
87VFsnKU2thKxjrVprlPA8ZJQIrwdaO+GS1kOBca4IJZL5so7iyFe/C8uBVdZsgAC6rAmM+nsU3H
sycXLQv4ZPzkDWLvSJf/rzpJnYYcFlTOZ52pdN/TYCNKy/P+JlAkaJ0XoA7nF3PlNHT07WoWWKOg
dmaMy5ZA+u8G3KpPEIpCi0QxOlL3AF7Vf2joCpVVgc4a3ds+o+7ekh4NRBiUeMdbHPZh9Qir6zgu
OIQjOxYIcfsJ4j3YQfbYqvEksAHF29v+NksIaKDx8YrNyqLu7ptyBKoquqXU2R5MGZGEGi26Jlab
gM35FJpGZ5qZ6McCzJ3Xofy5j9i3uY/MjdXUmdKD3/eslw1oS4qcOG8MVW4fpwycWztk7B6Vd9Jk
kQZTX8L8kpndWqt/zs7z8gw3bLPr07ps0eZNIotYNVnUTJq0Ud/0N67mJO1vYDSpmNCSqIEjFWp0
/DF2ZFQ+UFoLsjdLAbjc7YNnHysBdv0cVKPKBmPjnA3+gwU68t+B84b4szFTYLMj25L0yNRRop2I
uCB3N4is287cEbHYcxqkJAO6IanTUehYjArtnxQBvFoSvT4VLUn3h0n4QUqfNkm79/PCOWrurmkb
IMKo8yEBhuoAjQcmVirjgkd3QQmgbcxDPBpSzW/l+rllz5RCy5RuK/Ls53rbncTlZel2F0DM9Gat
8YUHHIl8N9TD4Avek1DL2VwT4o8T2S43n3YAR8F/zVZWsr1xllJ6aNIxORxK17H1wZfgXAxTCSkK
Jd3QwNeF8rpgs7HB22kXtvVoUbNWsFZBvcv0P7Zx4F4NFCcvSiXFk3hSU+MPdDSZKyCOnNelwkYn
7wxGNIGBm/np9yuiHl2kIigcd1CgB7IsrXpB7FQu1+fJxijsp4rzHvGaYiw3kXVPgLs0gzXudJQG
iPX+qeor6HTL3sZi9uWNyuew6xnkf9oimdTw1CQ+VfBY0pLli5iCvZSZbNCsBc/dmvEtL6X2xaX1
S+gavOmNU4T6hBSQPicBxXW25XO9k8awFRJ8pnTnAgk8tlWmdN6Y2jfzf2DWz8FbTKxLI1C4Rw9Q
5nCUcCvCh2MTTAt4gfkBWbYK3SkhufLruWCizbRBqvR6xj2eIVxd3R1XWQrQq7buzIi6NHVY5WYv
LSeTnyN5un5puxRhaK6OasnW7JgsTJdsxtVztC5xkWW6d1cyfnllXCI4LOMiNtlYvaFkEfGg3Pf0
j13x9eeVMYNWZW0NaGNZuJNCbJwxO4Kf2awMnGjuMIQovLHLS/MdYwEZIDguUY7lcIhwfgGsuQQh
TWMxXvEp6Erq04JrKufqKH4j274lluuQLwI1TqUuFth55r+3LsDM2cUlscN2BrBLzc00t68mOAmp
2UuvEsijzCjUt/OOjb49WDBCH8fGyYRq24XXeJaWxy0EYWhWHQy/uP92J2HI8EOzGJXnIbjt3rED
kM1fs2VXxQmyvw+K2HMIZzJIJCFXONGobnpRl6Wwew8YHA6o9Pke+FrN+UVPrwdMx2cQdBLnccFf
Uz/Ojie74TjLDFfBB9pW4oOV08/NWIWCSI85vSh+NcXxJ3fi/azYuyk4sFW9iFPEObOmgMjjDGPT
VMyTVB37RypZ75/tkWsn1J6ZAVcA57rf2PG2mprT75E7ddefpVD3kzDXEAuk59qk2m+8xlTd9Rf1
fa6FD9dMoE1UtdJh3ydHID3JYuxT5hx0cy/HflY+Y5gTkB+o+d2zTp39A4+0u7PnfasDBiknFc7K
zwRXDGdPsLYkgTPkvF7ejqAI/orgwlYvp5ClXN/DFYnsKgW4Uq2aVOtgn8whzrWewyyaJCEsFYbG
CP3kKjF9KnW8QRvLDflyEBssiv2WrVvs9+zQ2Ef72BXn/CYRb9d9+P4eAyX6C58/BjqVPuam9nbf
6asYqb73McUNPoH/tsmySWnj9Xg6BXOZ19Oid8KJEXMbB/I5xsum/FrWj2x/+hDopqbf9nM+dfgv
+bOssaoY5rhz80co49CNI2Oe2Ubs5ekjqb4HwehsUXTF/0IWJupDmQTFqYUAe7b6dMcYm205nwbd
HHmMsvz0X6Z1QtmBlK/IN5ggRGTGpbTa2Oc7Ce4XxRXluMUnBXra2gzw5xcdiROuDa3d6UpYu0sI
ALc+CPtI+cfkSlRyysfvQO4cD2MScZ7+TNvikfW87FDdlLgxGe9DI1QmUTsRoz81PQAYNXD35G1L
emYtneuq0Ke8/v//neypk1jMiCwsYznzjVhZ6VCXFbmpiVX4RKZ4MeE2K+1Hv+b6xj+144Mjj9UH
AM99e7+m5NOkTUc4lBLH7JMMZYbrIIvIZ0zfH7HSJfHsqlDLC7E3PH7d2BQ92hWZh1z2c0vpNqq2
wvd+bpjRKrt9pVNe1H/4rp7Rw6WLb5oAOjXp8xcRDLb7XlihaMi6KrOILR6XG/VKRt6A3LWuKS/d
oH6d4x4YB9nHRzwW3QF64puqJKzWDSSsSWhorLmbX3RFbutM8cy97uwaZL/T5ZYDobWoqrgw1ZcA
UcXhPlETG9WxElW+HaeE4WqXsm4IppMLZssJIG7GwjzxGK4Sx9WpJXRK5Hr/IELpPSzr73Y0aJ4/
xuPE59Mxv2tul357uFHZVKJcubul88Ys9R/a387k94mxnmBDcP2aC4kpDWrL+HjNbxS1uBtJpiyG
Jr2oXwttzNVEKNodbZrQasihKNXqWopMPtrcj3wKB5p7x1y0m4iJjuXY8eB6C/G4nuQLQeay294J
CH//6zMUeRT9ngZhVnSzujhOfTmceW3Zv0s5iYm3tDjdOKnqYZ97HKsH2uNldWMmz1zuMRmy0drz
aUo5gC/kb2CUyhtEIXE76Awspv6SA/if2gdgKrKom1ohL8ouY1fcgD0NCIR0a54p0b19W18mr3Cp
R2whStZjLMcUPwe6WRj24EHiI7ZR3wzvTdxWvIvQRXm89TcXjWMrYPrV53BejsoXSW1JQUh0PMm7
xrrkKjZi6Iti+ydBY+SF82s47hvW/VZzjAFqLsW6ahq/Si+75scmzk6gD0+WpKdYqcf86fV1+Blv
f+Rfunm6gG7ju4ocgPmJGASAMLQ/6Hj5NcF3CrolPhDHRUnI1kdh+gyKpPOQKNQLryqkkni6DaUF
U5Gsi1EO3dyGAIf6aJKaGqqjnsZzoEnHYdL5HvDCCMDDPbqhg95Iu55pfvxCRjUfKoBHxklnzTmn
1mxAC56+whj9ebNQ5p/ZjJoxN5WSvO0Ynt9O+VnvlJfFcfMfduYDQicmdjxLkAtMid/gJ2Fe1lxt
ix9zuoICvUTG0VBFx07p7FXSb9+S2YS7yE//1rowiTkkl+c0IqbwP9LULa622maP1AHYjro6pjoo
FZ5HUDXxJfQJYLd8D1QhY7TQHkciIdO/C/HDwJAOy0nVPSBorg3vTNz7D5pprdoSq2sNXZ+YhWLt
pd37hfZu7Xt8UO0JrCDNlxzprIx2ZxQKCqp1NtBJNOmkGeVi3Ntep1BnuWuL4YBFxr2sGsnBata0
GkzWIWdbZ4FWt7QxN0HZZNkQc8Psq3ZBewlhDVm1nm2vREma5QL8++p5nfJBvgnfe2TGlljL0n1P
N7SoUi29qI75Tql4mP13UYJTvvAGPZYxbI9weybLAFDisOlP7zH719lGwDCrI2Kp3Mi7SaOdxo1e
w4h9Hm6jmqLO4ZaNnsuCnltoISnE1iRRzmeqQCB0xDVgwYWIH0/820BBUlZLszn7xAZ/MCl0DWPb
wr3nNWZ7EL0un0E3PF9KQNo6FHOLjHo8fEY5Zi5Epnay7C4JuClB6/cz15FaPAoVzah9WQ6MMFXB
PMHwlkytiuSH7Ge14MVhRCJj5tzB6C2+2u5L0AUl+kXthuy3QffCNbC89AoIBkNUsByMc5HNYIz/
zqGOpMu20GYKLedHHaM5oH5rCvhMuU5X6wwUuYtHcyyXn6WegEaZsQIatKYs10J25OGEaubp8CH+
WWxx+0lGk1+Puj8fA8SNvuvraJ2ZBLA/q34Ihj48JmcF2TBusEDT/eQz560Iz+hJ9OoO8nlO0P/7
ma8udBW7ekL7DSE3S6if9DokgxO0iMLQZAHkDQGOnREBw1vZT6fD07fxHZDrpqof01kmb+eeUcwr
/Hu+kvjvEp/SVwyiSPHALBP9MwlTy8i7RJtzfDdOV+oMSI6Ax4PpkNJGnaJ0IrVnCggleuUOGIdb
2ahOAwQ3O2O6bjVCqOE1vIyGsXKESRAhUBnx6zFnvcsWhjWpjifs6+p/TGqWNDd213MnW8RYdGNh
M+v4APP3LWfw/CF/i8XtZze3h8Sr3ctdvPWZ704c2AvBS5Us5q1EpwKDsXq+88sv8d0cvGm94kX1
orPyrxsY3bsWSkjEbALe1wKAGIQHl9rWEkecx2xuh4T+Dz7NHvsD27teDwURA1uhx2eFb5faazex
vhhphogp7/7gH/L5eouw5Hq/Jsche08chf8YraH1dvkxcYrCT5P/C+rbto0lkD30bDXHx6BeWV/0
hLV83X0lBYfzLqMqu2RrOWs/7gqtultqkaofYVXGWJ8LLNN0yC/n0J38lXtCn3ZSvU9//rv0SbTt
of1seOifqRMAMQlRlPEdp0Hm9B4nGc//muV4s85rdM9O0wVlPk1b/zLhxkqO7Q8/awdD7EFATlxe
BpZQ6ByCXSi9Sh97k7XwHGb9SlJrokIMAgJRFqj7Rgo5RUnaEm+FJBqaBKZyAsdvvwBPiOUELE9Z
gwduqZJ+e8Dpw/WEZBvrJrppUQXTjHod8X6W11+8+FZJgIVuzYrZPDciLiATUWf5R3/fBJwdVQr+
Pgl06UPcxulmkBUoTKJCuxP+MZXS5E3Pv3WbtQ62bMTfqt7aB786/fsZLHAUkHXzOfhpBQc4BazJ
rTPLpGlhVNszq/+nP09DY9dhRP80Ls5Fc+VyDwS8bmyKmEBIYMIoz0yroelCiansHow2C+TDc3Jo
PxnTGdTu3IhIr9/eAUTij9mE5XGTboYG8Bfl82NP/+Tj53N4rU7opUfSHUcjsbt/6IgLEyL42lZ3
m+kOiNMoCd26aP3JzYZ/Js7asMUB0+HirZTbdrQ9FN+NtvNlERwwxXserw7xqKDAsuezYnDtA7wy
zmMIeIcupEtpO8wXTOMG3HkzT6rc9Qev/OmiJkvZzK4few3zvs+HDYht0z4GrCaJAg8udJXWQ0yM
sy68pMdvC/prfxXWPuJQS1j1xqpaXXKFje6HQvOV1Y3chKK3A3NTc1DcK6cDDeqwRQgYjr8ifo5h
kAVJvFzHQRXhQODsDSH4X2Mq9ieGYd4JWh5wrDw+Cg/lGbG4CMu2gY7uka5wqrdZJyiNKZkUh+Xq
LUHKv+VBlQLG/uaVVpn0+8fQIM/bl5+8+oxR7rMbahjJcvqkg68CsM6w2IsC+fbEWt7lTYO1ypai
TUi2ns1+LB935b/bADEXrEXZuKmfDSGZSYzLad3UD84LgCJ8tnTbep0y4tD6TLIfha5DmGVCUcsg
ZVVpprKnH5nvoH+VSLBXYqglfXDAW1bhGxjYwXWU2g1GKsToxMan6UYCHA6B0OxdXgOJzl44UGF2
y58Pz7N8sqJMkHRrmaDUKotcMsQfURJVa36hKILiDmMd0W/wB/URUhffvEksew8oKxmSA9Grooz7
mWmkP8icIahF/glo1+tjL1yRiwekkVLs53jZ3nVai6pm0HZC0WeMXzVFhVwECWRUoQSSc3nvfqW3
IwlePsVj68lKZylbv+Zyb17Sm6rHTaux9EmxGIbc17/LKCmw+AdwFTMtVBrK0Ix85LgWkDltuhzY
xjDlKeuqrtiez9Nj+5OrCxG9CRbP2McMxt2lDUqd7hz8SBS1ndDezMOF/Y+NMNx0ClZgEwUBgj4n
zEW8oVrjwaPwLQbQv7v7Bqa7YSj/jhTxCytjDzajE6yFSymlQpHrs+HM8+Aw/sYfKTcQx7UuBztU
XQ+uqo2uNOPikhz2ZNQkwWK69SNjkyRQuNGXotcabP6y1wRaJHzrovCdV4jWnUOjMaRBOncUtrmW
hrp2DCuePHhYDH7rXgt/urg+LsRaFgw0yWxqn0xe0tKuxuyF2z/4dNUbtKakPRfop3d6HgxkROrj
7GVPROBHQouHo6Ro/1Aqb8B27zSEx0dqnw0WVsTIZ/s/dcx1Cxd7NIMtlWfDd/GaAwT7PpbEPQFp
QkcabPIu3f0t2evbU343gOSBWiGlzvMDYU/6N5WadtbOon7FdwBO+4tGLAVWOw0dd0F5mgkJNAUE
bD0gRlDoF1vqIHkWGVrDTiKIih6xn39qub5EnNzyA/iBARfYVny7DNdRVn7NUAZsQvn+1IbmjPlm
9UlmJh+dEWKyBW12+CJSvcP408aLlosR2uqLsO0m1aQREwHjA9skvtJoUNngG08orPha3IaEzvi/
+VWI1MlbVPFu5tVgih/1uyXv9MYIuAvf7F93APf/ss2Dt1I3PMTt1/vcAxzCetCyUpwghz/3JGEn
X5YQZ1haIkv67ytrYaJWLcRCWiXHQa56K8UTh1ohcA8BKgk4ylvdWhXkJ1Tw5FErj3pdVcAI4yr8
cM+TIrSTCJVZpD5CzqLbWGCHF2odS+0ntBGxmhKSz4DGabDX1pgty0+yBOs4k6q54C/kWj+Tdtrk
LzQ16J9LOkN7f67zaX8te8o9WHeNJpmMo+BLULTnO4sj7hwPSvaZqpCaHOY/sqxyylnGyW0OVxGY
6+CWZRzmVeWac5I88K+5YvTJQW584OEdBGKxPuaVvFgvobNIA+EId3AkiAWsShAc54s0yYLgyJhS
r7B1plFU9d80wBD44lRxJxzOAZQenIr5+/tpT2MrASRdGjVv797mJGVbrh54Dn2LqseSntbBTg3M
ov427DHFgePvSpAzXhG5BOKCBkdBV9QUpXDqvi0TJIqWsHuuQoxYf+kb/HLQavFIvXjaw6JXS6cj
DLfGTzKX6ID7ywe4oJDGVK7JagQPR3zCZKN8gRz5B/Ilw8bB1X7ADf2KU3eB7WpPz80/O1ng1IzS
pthJpp2t4+bfw/OD0E8+xHvLIoatEN0PiKU1PW6XQqwlV858gJbz96SVK4/4ToJJcaIRsAhCiaGi
wTfJOgCb6j/ypGmT8vbWU4HpHfn2eX1LSX93fhOFN+HmQ5aqt5O5ydlmG5l1eq+zASbmjnplDsR+
BNjjiV8Lj40E8aIfjZLoz1J6wRrelGRw/V6LMJvb/EkwemwoMGmIamTcB+XI5QnAGNq8Kin9xEj+
phHoOsVNavROKuZEqikOciGVlJidogYhF0suA6aI7JQJFEYhjvDeVefIEDwrpVgl13Z3Yk4rEo8/
QE/HxZTFIbZHw4Iw0SPHYI9WiaE0MLyvWH/Mw90u+buDDJ6H3NVVnyBjI/unwTy5Yue4HZ0k5ZdP
i1enYWvoj0Yl1nBJePTYibdgMIm5yUWneyZ0PuuM3mPsz3+vEAP5tC3OpaKwnkwfsqmmcBjdg3hS
2dZb3n/b5FbX1+D17h4UBvfPS53F4lI229AWkTdtkj4HtuXkg3+N0BbGHf2ltVPt5JjkEIqtZmYb
my5wIewGH8HD9ce/1JNVzirg3zZXxoMHa5SfJ/niZHKw2F4cLAaPtv4YMcBsOHhqZ2QAdShuWjFq
miqXp8aA2tjkhIvPk+hYvtENEiqzAtp60I4wH0VpuFgOnHy1niCazgW/w2AJcPF2ApuxjAAVmZ/Y
VKhRBh1H/aiVxGyhFpAEX4aoCFCy1RqiHYfhw6+eOhS38iuoCpll+SOE2DKIGUtAV+2qdFmG8a35
SMZYUOqGzilQXgTuPEz0PKxWTmx5MNXfRHCyZ2DwATk0hF0FNKHa9t1ran12YgsosvrTrf739ajR
HGQt64WI8zFIjfqIx8C7SOoea0wQMOnsfLPX0zPoDlkFshlzfJezMGMv7Wgs02wKGjEV0BhFw8UY
qjh1ALZGKfXo5Jjy3E/rncMaSfloMoHdIv24X1T8+erhSZlLefOmeKhD/krD6B2l4zjrEk9+xU6c
L4UxaPXoA8XE984sVsDxlwTT11tWliovqnz06AMdLbKIodJmkw/7HT6iIAUV8X0pqwewybCwZs0m
2W4nueT6HrACvWMEEaR0WK8ynGQmF5kLcp7k4QXPeYSljkR6a9oD76V2ojvw/MoLg2OW6571LQiz
RdaL7R0z1/A98rPusuUQzgyJHduum1UrvaHt1sdb0BBnA52r8M2sqa2QkaPgXP5S3FgOE5WEbx2b
J8pb8dbHJrI1zj2anDTGEmXpBelKk4lBnxKfPyTq+60VXrl2D4509d/wdDfXI/zrrMeGbJE5rigf
VRnCuaGdayRiQIwPylPBnRJWwzOYQcjAl8dRWq539Zfojrw/wqag2pOskyGqbZ7mo8rPveXFHocv
gJEOOWATnHxtaDUGVz3dYwZEpx/m+CM8I8kXsl0ZwjmsK6yXXdUJERMgt/vJEgOJTtzBWpO7bkwh
BP3NMz0HLd1NSdAv450ov4Ur2VHyZBgIME4JA4z53Hdu/IUN1g4Y4sYaOtB93dVUA16q3wo1h3Sd
P94IUMeubZKfT3MoxdtONIlqWVWLJBoR/BcHOviMkndHkzxwWt+G97lAXD8f64Nv9wslhQWc5lUM
VGAPurOiQMmIYY0h4J9bw7ZFMyzNQni1rjFJcGO3iHH7N+cqeMj0evyTR+AopTcgI6HmKpeCAY5J
Yrb5HbvQ6qRNhx6nZePCJLn4eZhoR7aV7DCYAKwG9leN9qCAPZMyQHIrrUQMlDD9hKqSoJfgrrTK
BPVkPI/jZ8VUWPxMEWeSnQUurFv2wshLz/TmF5jSMgJk8ohPmgLaaJLPukrl8LAqHgYh2zzptbKp
/EjZf8wapPhCXBczz4WDfEDStcbu7JdnMvSnOeYkz8h1cugePoxyhjtZzJXc7YvAqxoJCZB028bu
U+IsEfu7faNahX2KneFWlzba+vwVYx6okuMUEqAKkNrMkNFC21OS90Sj4Kj5eKblmqY9JVK2XCqm
dJOk7eAmdwp9asV/qjNRvnIa+96f9CuUUIZX+jl/tsF+oLcVF41GzhJ8m98kYyW68VnByXHw0nT8
IQOe3MsGUoNdKHNQXxqFojLp9+LN4hJf2Zt2xroH+3pA4h6un9nXA025MMPOU0e2WVROlHBKCtXR
UWF6/Dt3Wp3/1jAl0KnGk9xbW6fev7KeICnrDa+XB1V/uO/QDx119yV8hoSFR7jGMwj7mB0TO4O5
2DFXx+TuzrHWvjIhRWczFRwjqnKTgLl989UUqEQsUM6xD/v99n5Hs2JPxH02dQqaz5cG+QmdGieO
U9AwhEUsA4VB46bhDMoTAhdBZ1vWaTGg7jVtV6ikmKWonMsaU30rq8NdeQtt9AB7Zhr42i8Tphbm
7F9TDPmXNpEWVBmEMGHgvmKA3nMN2f4Ajazs5T8PUiLWqEmHa4Nd4lH6hxAIbpnyZKssUgB/jvpT
FMvSW+Nplny6h83DGWE78Amz0RXMWjkNjvEePZF58/B96/h3bLhPAtMgTSRrayIyf7XULJX2ioBM
Vhg7BrPKx6IH4P0d/OTcC0g3bUxrzsyMt93XYwqR/Na6wEx9aUUJICSYNCX6Nale20JvQqam0tJz
jvyKgGQRdiKfVGBry3SmZGBbR8C0N14gJT28PPOClxMF7NStmHpWVJ7SkYSRt2pcolie2e7XbVmd
yTquDSFOY4/XXolQIO99Pb8xJtK9aseuuQt37OzhIFxmQDo5kHS0UeJZdIVpt3xptSCJQno5livT
pmWlzU9xFTdhL1afhx9JJU8KXEzrQpgcjgBHFHwcTewxpVmN8SpNSwPEO2wBNuife2Wlx+tn5I95
C5LGky1Aci8zT4A83Bc2z0kfI5R44JmB8EHhP56apB54kgbm1iALFBVdFEBT7XG4gkLVbmAF8bWl
V44W89eUzGuXP19Z39oaWp6f10Qlgq0R8PccI03MaaFl1POd5jxbbVYv5csHP8v2Yq16pjnRvkY0
BGq3QV5hsTC1DIhROVFHEu5Ep7T4HUGTc9PonhxkTs+xNh7asmzmj4L9wO20ul62su0tdnHdqO7H
bW5HHSK+ZNFkLkYEyrzQ+lDPx/GfKhiWuKXExRzUmtuRjVxJzNjFQ4TBX4I6MUtDVD0O2HJdq6he
Zx0sxSOIyY7vx2D+jB9XWVLzIw36MCfXcIQoOHDXLsJG+gpUry77GACRWm/J2nhY92VnjKiMj9q1
yALPU8d54qA4ZFOTwhONZcgZNYo16QqlQfTzJlZPMgo1SwoUHu1WLgzTafTYz3CgBoChWfjgW7Cm
my+2PoCoFTiiwt3W6sRLC8ohhw31PNIdAZxAXYdnaHigfgD8FEOwhuUgtUou9MWrUiQEUI6IAJei
aq2H4XqmSeDuIQjQ0wN74kNudbC6dH4P8NYdViJdhbOzYclFcSczKtguIKBHkPt5HjaV9iWfXh6Z
4PvovEGLD4Y0HUTqEClHKM7SeziPHJPsU0ZsKRLkodGok3SOflZKTPkIWKu7+/Vjkgp/W1XaNVGK
jquW5DbnSmNi1nxk2zihmZfFFV0n0Sxx7+nqDYwLAe5Y6C8jsDFmgsswaYQVHJhfA5UL6dG9gmGo
tqq25a7fGHqLpFSNRQwTokTD7UcDKLbv5z4/E2ZnvjCW4Fg02tgzdGuPfkU/lkLHifTmxYnikHu/
+1gDM027stpUZzXbri8nHXZwSNjjLnUcenZvNvjuJ7E78Q+39ptaBGgYtwN1vZNaMk0VDnCen4Ql
fotLqOfJuWdPtZ2rjpQkitQO4bYNUO6eQeWq2xyDiY9jpULudI/ejL+iErkxDxmTVbL/K6+exljW
3R8jsZSgV6HGruEIUyMgPCu3EEvHcQa+8vDdUOykAPta3Rgu2A1txig3Zm6puREncKDtBRqAlRuT
sMuzaHaAn/fiMV7BYzbJ1Zxs6hahWjVO8m86NQL6ZZ9SQatngr/iV99SvKnm9G243LIHMLUQ4AX4
fjerHj6E8x7CI25E3Pg/1vveM7MIU/0WEq4FEQ5m5or3Rlma5uOqLx77y2z8O4ItlAnbjmZYRQ0u
sy26lL1HpF6Zqwm8n1ACiu74/Tg6V68faf3eKlb8ObKyG9uUrfbYP1QGIyGd4lQ8m6jtJgrKgKqe
gfEuO36fWpFdLrnTOkCuI/uAOMqKc+5RTBzVV3dQpLBXAJoUgaQzi467z4nxc2E6g7fAXSZrKznY
uTaapPzf7NK0ohiezgOHTcT3htdS5IHdJADRhlTrs3Gqt8RQgYEUKn3twSqKlHGWECeicrYcdk/n
BZ4oxdPwDHNFnKn2TQRVNTm1iZHUWX4Om8REfIlwrZMWcUg+ALAIDvnXtomD8vegwLnrV5N2LhLI
5RC82/vr/nlabFN/fFKJPSLOfokReKMMgJz0iK1yQXEGc5L6+jZVhJG123yVP1woFZjhDpJ7Wpm7
915ZWYKy7D5y4nu3+u1hFEFFp6aOn8q3wK9YVzWknIyXI//Tap6gWS0NJtK8cTrZ2pg44ez8Ctd3
19EaQYeHuCCMGVCB0ZK2Yf8hCqXrvWKQI/MkqgD3Dmu8LVB1Z/rb9wyHojMgBdsFStZ5X0z4q20y
Asjblo3ZRxYVdoXSCTuq2eRVUIlVTOCgIQRiwWzWCeXRmp2G7UzPyvcqCExJYomR3MiJycEMNVMk
Pt7okE7qOzApaPycer0DaC9mm6NHXwwmELfwXhIsQAgu2KFzC7WZyIdjmkEphh5LRuZ3CMHz9uAw
QNsJRyf87Ru9/m4Yj0nZVogdrxpDDBrfGMSH/EiIcy51dHxXQ83wFe6RbKJg2zOyujCrJcBhUsG4
MjzmieVQ7aDqb4KHGi4ZUw5tiPDivBJd21JVhm7qUJsgfWIxqf9cCaNQqpZUWp2XojMrYX1FlwRU
1OEPwNrz7lEUthsDqKkq0bSu1JZvzPT6/ktw8B4UhBFHHSC+bF25g3ul9nEkSQPuKMPLKGHZjjF/
BGCHdv4qLeA6ahWtTxdjkSLOnzzR3oeH7UB+YDCHUz9XVo4YPBYmEZ97g6UP0fxUHJFjX1AQM9yT
/ez29TV+WTk7Cr7frDImk9Jz9UwoyVCVhUvm5z9kVFESVxAI0EYZ15La6RG/9Qlr4E4cVyCEYboO
EcxzVvO71XpNvCoHP/Tg7Ejsv1pzZYqxNhVf2h/kysAetKO5BIIhZLc/M6TkefmhUCZfwkdxAqC9
HgFO/GnNEagtEa6cDtRWzyJtfXycs9zH/Vl01tyZeMHaPYVUbUUDwj9tIun9KACz9+9auXgzfXwK
2aNGwD1zP5s+qQ4elnnQ5Ym0VJlO1iavKE9/QA77I8Mh8hB3FucWC8NnnfCJ9kZJSll/bMiE0w6m
/CiSFFGxQLWF6IL05wowCsrkvsEnATSjbrdTIwXd79sDfQ1rU3WGXQ77KCt/kOj71oD2MsztkVk5
W/pzM9/0EATaWgM8yYvqt31Pv84YuaxFfzwl5DtpczHPl/tZwbRejWuaAS34ujtXwPLhJ5h3s298
uZs9n5kLx2mjxWwkhSPSwUhrVDAKcuno+mpaSdTCTouJgCHUC925T2r005IufNmf1EK5oxrFwsTG
d0yB63iLGZwOFeMT9A+RQc8VvMDV1m7bT2StsxflaM3wu5KQ/HLae54k31vuMurqQogTqXSOmakw
OJFaKWwZW0gwS+nPfe/Us7NNBAWFpxL4ZIT1DRjr7CACtUuBzLyK5Zq1nuFeJ7uHo2ksw0wnafsL
GvCie62nxhtxbTmHQhbAUeeUUpJXnC2ajXih6jTGxZwYVaGNJtXNoKn6Cww6d/hwcq85ox+Xn6HM
qtflIEB+7JRVGu4AM5ahwK0/wDn7JETTGwNfA/SZ7aJ3UzHIGdb/LcZiXbvFHyNGdrfvHSdrzZxW
QA7qHFcK26tMB49Xr2mZPBp+5dn9DO7u8lis6CKlAJLEmdZoH88YQ5KskckmWEZD56j5GKkMQM8H
UXyCi7sVwFd0EI5Dl1X3Ly2aPpXbwTgFK6IDELA2/xfZBRv7H2gJ3yx/bPLeDXZ5tXTOeoGtxbEn
+X5xzeow/t6/n6gNVi2VmBKnP7vtVleXQ5t8wWy/ud7qBHPVrtozilItjDkxh39Rbu6fnKV2Gp3L
O+M7CamIVfQ/KOxuvp9adjtkZRWw34dasysx/kRJOn5NCfWnH8FvQ+STZ6ri8p+yT+pXMoAvoTtc
ag4VgQ8gXPW/2dcnassaPnKGZ37QOCBHJ0p3vHxRUO2Z8ARYgTKZ+BCIbKwE/Du+fZoJlL4ppA4X
9sQMsU+Ctu7Pqtl+a8ZB3WZDGl+sbqza1TcnQ14Wbzy8kEtG3g5yH8H7jiSecNtFExn2cv3BKASe
NUdEGhQ/cGIWqVJr4ip4wekAR6Of+z2n+l8HDkH8bRToEOhJnLPVXrblNsCDfvttULaqLk/zwU3t
JQw0ez3A2QXTJ1Z7e/2n0q6h7jp/DrvWQiVNPZRdSOOiqFK656x6ipc8HorNZJy+toLuD4MlDSip
GN7yUxI3J1T03UV+XYWkA47Lcj8atkW9Ho67m0LvzRl9fcb2vitgK0k+LTIAAafdZ2jXv+x8v7Rr
wMQ4KGMDc34Vrh4XrJVbA21jD/Eqy/8hLd20OkAFo1MghYJ04kGuwr+3e5Bh54bD+tqo3VKmxVkl
IHvZ2IxViRTRKaXewTDibIEoGsqs2PcHGqeU+VPRsQPAg8/tdZstQqZ8JKCMORJ/ISO7OC3MsOuh
VokPAYeXvUjJvNkKy2gs+HNieLw/F9ArM25MVVjx6eAXzEjNVr6RAxMQFoAFsdlGwnrWMDdjN5Mc
6myHU2+1h7x1Ne6Wf5XdzsKLCqJzw6gQp0tZ/HIqFyXASAA37k6D3/1rNSZKJju+r/n9XorHGXwQ
rCjqytvLSuqNxq7bRTgs64vJWw2dTjlwJeXnieOUj+1raw8gyLpIAsSq/AU5+oDRJu6AXZMG3+Aq
SriqdZdBkc324EXHQ9KHbGCRD76zwErwyWZgygXpJkH3nY1OcpgTwNzvubaab3eGI5y0ngXXlSfK
FyyGx7/s07iqAhJeWODnZVkm8dRh/QWvQbsPCUKTSc6/xhC8YeY9S7xFTlu86mgSNDBQTJNsImxw
UClJgElbalQ3JtulU5uOb7juBTiNxPEi2ZgYZZyKBIbPkApx3VuL5gyX3CUgk/fpPlWnE2g6Anze
1O9nnBrlQ72YB3xdBOIxlVlVbsfEGzUZYA4ovu0yTxuT1+Mcv4CeZ8YWBBYvLHLEnF6LVAJdEMC/
mOIx4U8p2hb6CBZeB4XGgeIZu2N5IaPA/7C5oRx68B3MRgSx5QqR2g4+F/+Loyf1JC2ER5G68M11
uJM0WJPPukeGGk++4PHgJCEFdYAK0F2w8xvCcQwti+P6dMuVQW28uBJOLcY99oRf0cC803hbGDQW
RzuMW32peIurOQloAqXbyqjK/hp+aFF8oskROd5gH4qlSOO9+m0k5qhW1GyXJzw/X3NlVgvkGO9L
llo+48WPkswILDUHpLMMgVNRRiJcSWVItYvL7qvIy431BPFmVMgf8jLYiAeH29Uz1smNbbf53lMK
+dSAY0GKyqmuZWzIxtrLIjCfE+mpTpgNtCJPEIl89SX9TAz0HS3LFYdTvdLrsWqQDORLe7snY+/i
ZXwOEBnmtRLWYCp52f760Nt9CqiBryQcoilJqjqFmfUSCaBua6Byh0yEkvT1EWjlPw2rog/Q3WC5
Kd3w5KJRY/hp+Ln4gVCbagMYk4su5n0LLXfR3nDu2m43GDBJ6Q95CMJHRqewjLG/WbwUwaCC/QHD
K6OC8d2chGttdEmgAHogYqtUYOi+8ihMO0XnNZTR3dxCPhR6ZvDAA5Mn69AtQfZZ8Z/+czkDKN1p
i/Mohdj8potiLgQyLnrNSMW+FFWGLRgfI5fuE/Fdw3VpxePPeJeLUBaRB7t3jfwO0nu7RNJfdlU0
2Hrwa2xVVTIi5DynUpfe75CMASyAzoegu86tj8uwH4HbvotskRPNoBBuls4MO3SNLdOy3MP86WGG
v+DkVLJviawpKWTsvB04xzkoxGf45R7O87WC12XGSGZu8+2lft1CNE7qmAt38dntJ55nTf5t8Fzy
Qe56h2MtSeWtbXN1JopfHZbf6KrHcZNHKQJqJk9gOBpesBzsabB/xpoe3l80L3R6339FMXDY13Ww
XwcV1HCEvySh2Y5uIVC9LCJPFfAp7fxkgcWLXBR5oyo7boHK/jOZaALLThhTPDv3Y8hXXgG+klP/
CiWJi9UJ6kMuvpyurJD3kchS44dXWdtRC6zDixCPGOVCvzkF80kBaAnoX+VTGvoVvN4VEbF9d5ZR
JMs4VAfnk9+a4DVnRULUhDOoVjTCW/c9QUWZl1tGbWU3e1N3GKrVnFT1dMBRR+qzxo25WMa/0lnV
k+7weHIlhaTZPEkjojFKlXpeKCBnb/rZ4eHleDiPTsGbr+G9jwHZSeq5SiRWCLJu6YTvMo4ZQwmd
syvwitw0E9Ip/XwykqtXaeZ7pl3iQyQ5Jt26HVAN6Y66+NpHv2q7C5+JVtXntrs6Q9nOkSBYQvdV
LDxTWPvBCxKuhOO2IlF9yVE1GoXwyZHuA5moAQDj8RtfJprkzQvzGVt2VibxpE32EdPH+F3JvcnL
ozBoV51K/45oM+h0ijn+a8rKb1TFYPbH8F5/AMGz+vH5jNu0UltnGGGd+DZVhADGXwCLNEWw73qe
/AzG9ZWt/oop0yS7BjeTJVmDmahyAa3XsD5XvhU7VDgegkjujZg0olriu33GtiuwBtmlZD18y87i
DKsWPGtlSthAdNJxDa9G1fVNCO0FnvF1svHhSNDB9DBnWQvRh97yveMZcbPR0Mh+Zjowb8kp9/TG
dAK3hnVx1vE+seT9cyTRDpLU7UqvnQKMgwrAAus33vdj4uinPsWTZsKXjtvMl7kmHPlFH1/q/SzU
8YATT9fbi7wmrxX9wSaFhDl4EC1n+FbSiF0W06XWOM+iU5IMQmQ9UMCLJw5ImQGxex2xqoo3Bb/p
RM2vQpI5cNPDE7DWv4ry/I81TkpkUKXV9Ru5eCn1fcEyZEG5B4UE7icqiNKUIbbnSnRbd2LueJ9k
IQlr8gSyM+5IorIRk+VXbKTOIjWEF5krj3JdFoN2cFRkfDPg6xEbHPCbcAXXwyKk4CTKuXQkd6dN
0Ktyxr2VKdcCRX4KH7d7kE9RphcLLXX4dix9nZuyNl/lCLVJDlpX9S7uEScsLyOyeF68FMIVW6qa
zKETsDrsyTjXowtaoDGqN6XiEEE9+PoFEKxw1TqHWuO6qtCe0GCyjopQ8xFQziKpvHXKJ1ADibM5
JrqQ3mcF1zSndfM3hKbl23WTBI27fdaIC5MVoRXFC9tfF/ERWUa9Y1q5bTPwUlvQCjtkrVe46dnJ
0RGvsntt3h54kSXv55e9vW9X1aQ/zHlclRyzUV6Er740dSuVbEQUUIWzUjr7NDJ01QKFd2dhDV8x
2NSaiLxsUeTpUowr/Uxq2qFafKX0plPUN64vGRK7nYTTX/sOD6p/jLwbfUNsRFm9oUfLzTZIYOsO
ZH2nY+91MyGGwYZPoNli31WLXGs0gbfj8eYOtvGGmLOCSz1how7aqY2Toe7p/nPIGzBFhuxGxIiw
CTg//3d0BJX0uN6BBPkhZr+k6J5Al4WE+hbQiufE2h5sF3LiMU9UPXI83J+cdrZrMkt+cI4iGmgS
n/xm1uFND+u2zN591zm3VjsCxLut4G3OakFTvut+8TnfWJMMiMRcBNTk7yKYjFM9r93udDdLuSYs
XJrt2tNezzWUTHWLDhbC+aWjEuUxoMZszJ/0YVkkL8rccCHkyTvOwEK8r5QT089FaL3Rmz75oyNI
KiAC15jKbtPER2CU3StoGTnWXxjvqSinRN3oG0+zJQsSSrY8JeTrHzHDgfLmdESGHzEoiCTm++3w
5hbb7SmnymomWs9JtCEaBCDmyrGUaeZX4TwYTGc1+K4NTASo9cOoMt2Gk2rDhw49ZnpF4AL0DaFP
o6/LxfAj5eRsu/C1A7KIxH8huseJvG//1HugLO8yJMcMS2GaEgMdTSL2uTQGgyikW1Usdfrn0cqF
Bl3xBOwdQmVFKIwqMGp64CFk7C5j6up0XfnNMlb3N7pX1eswy0ZeF+vjARp45R1q/tX7r/cfAlJB
MFIoro+ShrVkwbPY/VE/2VM8QRh7KIQ9kAzLZT7pgcPpkMrk7vSKmFKv0Hsa96KOsZ0KfWvzVwPN
tut6vT+Zt1/HxNNUuC/YEiWf7uosTxHMiVNrDz9nmXITPqvhQN1QPRalri2bYFLkZM4FWS1Fs1H9
7/aqh91pSlZADk1jv6FnSWWbYCd+TcRIG98quSzK8Y0MkrkkMtpEsUiYzpCK8WepLfIk+7H6F1/E
KVfQX59fgOyZr+cn4xXGt+4sI9NtvZtulY6C7TJqBYzGLWZP8SMqcdyJCwMx1SwYI6f94trl/KQi
T9kuBxGzTDTYKdfvK2nnmZ0zk2HfoGCelZsT5BNiqQS/CGoBxztel16ZVmlCptCEqDRVw78c4c7W
oLQ/dfN4p0UJAEgzbIC9uRBIWPKrXw8WfBM6EEZpeMEQPKiFal2MV82ENlENzPu+tcqENEdAcPqB
aueQANmHbisjHJEJZpdmiPKJw6Cbu/tDVPJTlkVSzNU7lhBykO11ch8FPnRvv6N2dpphK0rNhUtw
tJx2SmqMTT2X7UjP1/Ygs+uo7iZhAmNifM1t/348HxTQ6LlmaX3BDi7oWqsR6FIy0I7KaaWwNRP6
ihwggW+Lzd7AXu3K8aE53m72LW7b77eTsV4YFBPqyoUwK4IXCbG7DbDWI+MDa0qe5puXb/Q0im3W
/1ceXjo1xf9rM9Hk68MGjVO+1/artEpC49N7I29XAVbI5kTo0niaiENEc7w87m+fO+YYSWjuMavV
erbCuroASfSa3XdJTlACezhYF/zvILOqiGc8c3MwOqN2Gwz8djkNCBNfAKKYgn6Mz4HQV/4TGF70
bjd9MMXHg+qhvOdvKzifdmpsf0IjaKFT2Za4aVhsaxxk9itCcNWj+MsB5jW1NDCf5QbZxSfSfnDM
BOCvVCqf2BDqULKw/uGcDN2l/srKMnv8MDgVJ9s9vI8bKfgb60327bhU0SRbQ3Nhk7Z6KO4ND9bO
R1jvNkif4hNLa2wmzlJ1x4jfkAPoG32tCIUse0xVIgbdcqhMJsCJ00hqFrwHeJylpVgnhJsbrO4I
u40763PNHZJ+G2IhhVgqg98YB2pMckAKjKtbPN63vMQud8TegCNRXv+DVo30XvwT478Fmn2gNTCa
BbznRGKwTW4Af2reAQWgiyr5XKsKH7botP1klAIFWiPphpXAi/YlPNnetetx2B0SZVCsWP9wmu5P
jRuJyouAZ7PnQDklwg0tmqh/WYAeI5KC0aItB0q/h3k/xX2OfaYHNSXw2s20PxWOXwToFh9GRyAr
QsAg6+E64W7vk9zJpzPCJr2+bgmsFJ9kEBR5kNSzXP1f2GwkBQFzT/mQax66CcM7S7GKoUvvGR8q
KU89dsahy2RiM3qRPrioEePPBtltMecV9A42H9KDlZZT9XEQDXrrVv/nUVvjFRa5L1lf+C5bRHHt
KkLzfYyTlfcabyjd8O7Ek3ICN7QZ6vKnYswFiJlwGvk263D+65AIlHNrRnDVNrhQ7gkzciBdsNrD
qbyKZ/Hz6u0dp1cgdVd7QbY6K6Cjh6hgKUl68u1RqU9hTW4SLX2N4qiVMm8vlQtpBOAVi1paaE3R
sfr3sL6NagOM6EbswdtWmyMSL3JFF5/vKShv4MrMoIOJIXJVzF713OnWZQUPkWIhUTmnRLxLA06H
Atg3dxc2OnO9FZ1oyhSvu3SeoNRW4gcma8hP0xeeAALO8nAh7tYLOmy7P3oKyu4dxTmiG2oxHGQL
YA++QIEZOYXg11QlXEKYSPQOIi2lZMZbbL4hX3AJhh1WW9wkTENDe7+QhhToON8FW1y2DrRWd0qd
owJR/qUCQBIudI+BsiJkl/iPuUQAL3x/WzX07RP4p/AodikBxNuqDNpdkMyklto+kl2ZMW9Qg+B+
fEKimD+tO6YMWFMGLo+V97dbtsngeQW2bed2Ox41zvQYWiW/9RrV6vC1+s3hgMdR+naD/85vjrFH
+/9GDxg8DJDVcVdZGoitbWAsIAd+sgv/2mKJCbTVKbhesnjaMdnv6X9dJQHTTZ9wMJBCwyyodQZP
AAfXjxSE4dpw19lIIrhXvdJcn+fgAruRn0f09L3xTbdDAOeUeondz1QYbPUc8Un82qqQL2QhLJsY
ez5tl8tbCaIuhYEGd+/29DWNemzA8NYmkoWLYwJ42LV3tPFSI650JbdOvCiN0YIsJ6RJl1KOBZJA
mSpLsMafuFqoUbocidCDLdp4DmcBLicG3MQZJfJmhbdoFw21g88+pWjYTKkRq9PWJ5AIu9bVGEnW
WSq56uNHTV8LMGxOSthjOmWLg8rK/GThFBYBzd2NghpPu3G2Y7mz1fG8lKoFKCu4SRAOEPbJlAm3
ZAuvXJCg4VPR1cTFBNPK0ccGjstzWp03HG1zyDwrOgMYpHqmCbzVGUPukDQmNp8XlJPniO/pjmG0
orRLwIhLTcQ0cubAP4jaCSW3kKSY1djRzYIY6q8DfPRUxPAq4sLlbI0cmi2jZ/ZbLgC9S1eO88ru
UG3H2/kYmqgVUXEgYJ6VwU18VF54yLlBf4zgjEeI7vlY0qk+G6EIbERKk8GdLU0g3P3FdfGRtbmX
RrFp07h6OJAdcFnfUdJGYukeC6B1dPBCFs32Fp8cVdLTDwIwIJFaHTmNoL1HRorhaBBR0wWQrlOa
F+/BsR1AvAN8jdyO8ia1bnLrZUkd3SdFq0tdbKMUgnatyaKshP3jCXLxNe5QIEbEueS+FQHPl6e4
Kf/s7KPX98ipwnV8yLsg+ojoubYvfeSBkwVd5XzjlEV035MEJ3D1YPiLxYRDDSjyFT69oDP83uBt
C5/WZdCSA3AoDEsaDgk2mVna4TwZ+VBBqZRQY4bzyJAw+rS0LWjm6WPcYLA8qE+ryDXBrkUHhNE4
7Gi3jaQmityHW2bSFBwdyoroQgBvacjoTG6M1rA0EhetobouO4Swt9B4TvXMnX5g/ZGX1j9JGuGz
ohXVWFEcsOui5hry9W9qgm7NShWTf5t/ShiskpDn+zk0dLD0goIcVHUSPgwoiOAEN2+/tGEjvTzl
HndpoX4anl2A1ZrVQKSj8jq1oun02+ZIP1NRg2+JLLQwEslT29b+eZU9cRJzNtgU9dkZPqKBQFpj
/sRPxn1u83K6pYfetsE7dYb2rS6jRzZgksd9TeKAMRpHLav+CN7i2Q2Lpf+JTzKWDkNOW1dCGxZh
jUXI4x2cWEs9ga0TwCD3ofMNhoqCv5ow3+zaDs6HhhknHdnGZOSsC5OC5raz2ib//DFJroTJmiJ5
mUj34pkmGbunfARMkNjjapT2UwenA5xpBLYtSoY0NHglNF3/GnHJL0Y7lmUU59ISNg+1EEJj6L3h
70vQa3KLG3W/mzwoOJHbGs+K6gNn1AcBPPtyf4cv2n6NMfXamWqgFfm33iy8B4LoRJeZPK3WMjmc
NosH68/iYnxSFY29PoBWodkg9TzqZrqajwzdHFYxn2fPZ3TCugGgUSh+opoxb1JxJOrc/gUhTp7Q
gfNoJmibZAwX+duH4KWNqOXmUFZx+hXmfCizUrliLQime5ZtXUXpwhgvsdwzl6Q76eC8TULCWz0e
A/igWo50LxzYmfClxsFDV3Y/ffFngM0eWmlNqEMgRDXklcIuSHj1V+y/riGZ4NgzhYOWlGu8liun
Rm5RUkZFF6o3X5tISv3WY1VlOSxL6PSGRR6/PYrzsJMnV+q/XQ2hTuSQyTLY5OBU/reox6xexkiw
n+GqO2OXpuPX2rDAbjVrGo1s6up9eiR7iT2KOITParHObN2BGcmFsVtjk7Fiw2ZCiiaRGuudf/B0
Lemits0kQjSbcw4gnCAAiX/4Y4l7qn3DR46uNQ/u4Fawz/ZbrDdwSl3878fWuMYIeAzHfiFivpUL
Zs94SIsgHsEOSTJN4dprqJOUqNrD1hlmHajbHDLfBIk0SEfQJbTLduaUlWAGiHwJStqzZyR4MwiY
f4+8fu1bRHTq341oYA5nWGHMzP+TtZsBJDcFF69FdZ6MWtm27Cucp1iQUBGXBHgy0Y3YCHFFWxUk
DwQ/i/S9SMlW4tfL1F3pMpzPdytZ6ICNIY3nod067Kl+AKl0vq9AG2sUXQFewvf/X9NQ1z8PstVb
4KxgNkXJv5x2uK3uETWboRrUHyDXjmHOczV6B3zM4fsn+SKVTiyVMtgvk4dzWI7I3M2+20DQUD1J
xH+9o29ikQS/Ab6A5pHIRN5CkJjr7Vd3XDfr3SWjMsZIh43q2EKChFjYjKdZS0K6rots5fvJu6Wq
7X9F42MMa5P7083l/aGt1/4cQsPq0ZdTUQHqC+ShHAiUmXzsnPQqlLOGX0vIR4seRxapurTs95at
3MAp6A7vrTKGZfv0LduCF9I1kkCyEmPIxfrlzSkgKc9Fi7WB03Cr73+ctvvUh058KsNnD1/vRrGd
Lp1Yg+TsQfQdITZT1ZbX+NklXdffazRU0NG7g8uqu0ustppLB9SGYLzNiHBAkLlZRFPT+LHOBssk
UF7z0bvvV04+8/yYknsxO1N02HLclnv+ZEoltFWH5Iph0OyVYGta/PxRpRW60CPgD3RJuMhLJr2j
6QMXQas4nDMP9Qp/omdOSuKQyaMEI0hAjWr2sdsObtMbxgGgLPFLAzgNDDkoQyt2TmqOgRWfWcBa
p3ijlo3ZteteBssxnjnIZRpIPyAzth/e8rVb4a/e7QFteNb2ZR+lXKwxR66QKXRE+IlENVzUj24c
ZN5OPULMJQwHox4+6EY16o+1il2X8S1sKk0UhxyjlwBO7EKOwhaYMQfndr8rp8OJ/blDaeopJFWs
qkmbGhtrX+zzZfI8WVwuoLZRz5eZQh35t9hGbtQpkpbqruhdbFgUZ+4QIM30hf8z7dNf97OZ6Pte
Rfm7D3V8xh2oE9E+Hv1fyzAQfZcZroZIkGpBkfJ7dQfA47oZepfMeihYerSHBuzQ/ebW91rO6isc
XsPFJ5ANP4QoeOMNSMGXM1at33bPIOtuFcooDdAtCWY0BRvZzUqL/AWZhJt9xpjt6onxhiZ3J0mW
wEsNzVfcIx6ux0Jzc6cUYZRoIvE2rQkHsuq8QflUOwzSL4k/4BDxBIOrMAVLoebjn+2ibYygmerd
C9PyXgxMoN1dSD20ipHZ9lh7u7skX+XSW/HcS90ZG/+5c/TL6Fp1xE4FwvC7lAZRplEOdlFm94ZX
Ayxo6WkFjAlw1r+qNlSGjJcEf/TECMlfturz09o7elt83sjch1jrN6knsli2aquiOlICxAosJw7w
6h4wxgeET7e3yAnkeXe2ILMp7IYah8VSdcXisBB/P7R2WNVKzmnQOC6nC1ntBgRgH7ORM/JNg0Xi
Vqe9aaRoTSahwkveX183PoN+BRJ0eDlthv1gDqNl7lbS14WoqnbeKreXMTNhmCorsdDoJg48W2jY
S6aDLSZz1mcEWT8XSZjt9qXVbFEyqmlsYil0SZYw6l0uVny3aWI03CNsV7FftrS6setdGFQY7kpi
nWFTMpniKI3oWc22I/Wqq92aH6plAUvuxQFTTpJ32X2U6IVSSoNiGSteVa4ALgLQSLSdMPgGnwfD
8yCT3/g9SGvdyZQ3nJs778LVAWyrQzjfyLNocl5tGBRFEL13mxHuS4HJiZ4czoTNNX7hHGsz4X8h
h+me4sf3LWbuQoZdxJRNq/tGlT/MrDJYMrXcodm9MxlW/ynZiE7MPX+bJq+kxK2OLiZ9C9x9Zvap
KHDFauHsywksK/0U3jkT6o9zUywGsjF+XmzxFu5AoASObP1ZX/237oV2l+M/czdIowT6Sq5PDEzh
7pf9gdq1vJLZxINoFlN1Y50Ufb0BtXfJ/DM9txGRSQXZhoq6N9jfRw1LabsKLLPcAS2vPKnakrZV
fReL9i12Fiu9iijg752ROgG+Wd2eVcsBi0QampXAVjEOmgmL0ntcp8na3Oq7QmKZrI0g/2BhXryP
HvnyveLgItB8i+SS5duhs1EwW+FrF/nSWNK0RMUm050ATszOJIBGhqnpinZlprnB6G98fm80E2U4
Gq/UT/i5Pa/345Ze2w/9wAWbbW4CfrXRzVUDKbJ9M9OT0J0BJva7DJEaitIOyjnztayVsIK/cil7
OhqVoL+CIzxaHct+YBrui87TG0fLDm41hAcRd9XCXCEuLmQzlgNJcsBvXuxjDYVvxthQsHY3i/t0
cunA+rQ7fVyPGq8MXlU7z+VusdUcBeEHyzULqDMxhnA1RrZZREq3UBE3rXdE+uhQv0GMnvpDXLAi
qdyPk5yNiGuEBMKCB6bVfOylM6Z96Lg1qiiLXD3+mSNVm4Rd4B/2qLOH+fyi/IFHJsLWR9N/9KRw
qNnXsFXpx/tXl+HHH3UpGK9x7CK+ML99fh6N4VH0plWZkbNWZOIfFfs6QtYWEqdo6Cmy1yFfUUwl
6WbgWod6W2v/pKa5vDF+RR3Tzl7+4JcCRMOcuymaaBvK4SRj7XfTYPtMQIqWY9tHbpX7bv4ZIDs8
DS2FeSdoEzRnyNyJ70LPBeLX6FEZmU7H9/IMH8hleE574pTHlJ4LW4/Zv9t7fmVYybxwJtNtwFuI
0cPqARXETzVu/DhrJnh5GZKVxk23QK/xeiUZ8pQAA8y3EF0qHao+vFmUEnriuDtFMWpSeJPd0Mzc
3Xk40OBUhbVTtHmEWYfgLK+RKtcmss3IuW+st2Yqdvw7biTs42K7tobIVTa8r2xxqEk/sCYMa4aS
oBejhQCXmnEWv+Xq2a1aohrtXA/j5ZWswAvNCT5Uc505XinqMl91WpYyu9ymfDCBS8zEoie+2FTf
DmaQuEtbxDqmeWcSC9nBN0fmgUkSqHgp1NTilp9eUjkedPyqsjGvI4u1z/J2XTFb8gHBAOG1slqz
v/hy7jbZpjwOJKIansjBJ4cTFkD/+eQ1YJjCVj5YqUWta2T/YLWDDZVB6ZXXLqMUBBN6WQRuT4DV
IXSuUH0eNNz/9lzL/C1I1KKfPBXw7u/1IeHDT3ZLhx0Kt/tTkv4hsBZsJbgriIoMouDAHCjM09T0
URBGlAeEu8//r7W7gViXkYdq00Zvnl3NI6e7kUS5KSpXirstvRS3Pzlxrx/EMwudb/jJuQKc4n6X
rjaN5UJDUfOSwzjrTgVPCT+nJSY8muITlFNeT5L/gF6yFDrmrCSYT3ePnPHB4gi8Hwr6Zsh9o5YJ
AYN3ccZUWKR09HOqR+YtkCWiPnZjuPA2U2jZIgFvSMOEn+2rJl2pCZHOmFzoJS7yiSCrqYrlPPT0
Jl4zmqKD31ECLLw4zkpFu650U1icppJ0+gm8TI//Ut7S2cuLoeCtOG3ZxxGhWPEFxLU876UsLCPp
j0kEvDHl7qloItApyMQFffnhEVl7sZbyZ1/WkFg6qkr4dJwJholiOPP9XiTru1V2I4ZKTyCmQGkO
Xc7XKG8GmtTtRv2RAPUHjIAZFahim/+xiEi3yCh3ZAZgq0iF94BMkYNmZxDn1Pn9ePgAmOMvzi11
/zWW+W+BkQcsE35X9rv7+fUP2Lzr0s02JQ2hNR9YolBG5lcrX/wH92GccpDL+ly/yQ17dwhICYux
0xedPAthFxesqXluc0oDvWPs3a8q2VRPUENeK6jTRpJyRsRDs31yklmX/3fyKxQxXxRAMH5w2TSa
2fL2URCqqOyt6Huu361OtCDhPqruWZNkXabFFkim57wB37VsUUBZ3OGwvOiJKDhGCnAaA9PkNxhh
rgAxrcXMHL2+HfbO6GUAP0ZR3ArwHgWsrBKiPq5uMnQAbGDlMbcecE0023Pvwp6o4sJaBI9V94Nj
3nVIv5nZxbsxNMZ2TbzH5GNBdq7v/KJ/Nzb+sQv6kMXVBV9UDnuNl4v4vsBgO3LQj9AnS27mpu9Q
m4gYaX950OpjmCDWpNwygecdtmu6hUbABOonHtBUe7xOGYqPvNO9Ma1jJSTExWDYXDQh2xRl3SBM
1joUZvAnBCo2NrFzw9BZT1zJK6yhHC7dac9o7iWKiDlQlLKVGuE0aTG4yWn+ulOINIKHFloqFpVa
KNBNxZfBp+vh+T3eTeJPqZsY8ttx53Fmf6030k14kjU6igzkm0nQgcjgfflUBqFhfpeWF41pgsH6
YoQRJ5Sd+iBETAlw/m7NMScCtzmAEzXsmHVJAZEahY7sV5KicG6Ak+kqOjbmFxcEm/EUtzKSIGqx
jZzOzJEUJYPg8wQzD2YZ7G/xZaM2XGCl8vvIZVUhRhcJF738KtQl0Pe7M6nweUSWEOhWxB3pj8Xj
2HJ91/i6Fq6lkzYP0fRPhgdqWnO9EgC+sUt9MFqVG24n1HD/mYG9UOXJmp8+LoTkZ7PW1JTkJZVe
XRiDT+GB7So6fbRUbuU0SmA5xSxUaNcvrhMrQYdkN0IuOkf+i3du8/WI67CLspFE6gFtVVullNQJ
sUEm6W2OwTXyZQyonwiKip2ekZa3xEoMizsBSZDgVz+7jXHar5HtqO+DvgRyPXl/7/NWmB9ViniF
IXQ5sYCQ1ZEUTd9wNzTUHNB1LNI4VelZsl6TV0q/2GusypqB9418crUurEbsYg8QVakScnVCn7K/
o+4h/Cd2HxgaoO+3SK5djfWZDB7+GiG6XtuyZfph2O4a2Kf9BR6nCSyE2Af9/56IpQLwjZ8N9Lpr
0ZpzlPIrIyxMomMZVeIepuutPFGp9uob6Ls2JSjWAWzyLvJKBZ7SjOd92TLv2Qi42XiSkXt5ca9d
ePSebm19RI0t3eBQvBwt6O9gO0NDkls7Ww/6yBV8+jeQuClKXO5Wqh8Txt+fShRX9We32G3f54MB
aeGoqUB3oBoMtAHFxhgU7JoFGSMn1QjG+hoRLPi5InIS/IJD77UZod1FejvnqUtvGN/PL4PCN9jY
G5DgAURVQ+tFCliHOtiqkzq3di358muerVz0/LMc65l9e+bdCqjMCaAZBuyyZJ9AZB/Em6AtI2TY
SFrDzXvhmnZXBs6QJ7MdAExaXX6a8PKLCnfvW6bF9MqNOxG+Amr6LvLy9pfOpP3E1l1D32If98It
eUrM7nm+jxL4OHobungECVlPYy18ElUFtd+DLRM3R8MWp8RCdKqF2lOgze+eP1C26pDm0S4gcUWO
vbXAbAfpwy8zQJskSYxOzNiE+AP2ehMs3+n6FYOdVNwC4s2eTnpMPPgt6wKKFyyuQ5mzZlzk+TwV
mtloLMayMXybfi1jkeuihwqJnTBLZDGZgPwjMj78qBGWgseInCk+tkjxse0U/+gUA/uF2zScgWMF
YThSZw8A7fyyY7Jkbd9b6GOYIbTeCP7JlkGf6lkmeA4vMZY/gXUEceOxJ+TIAMn8pK8qE4mTI1c7
FQJWzKu53c6YE5swoeWBxMBbm0WT8yXkBQ4E0tySFtBmNvjroDjeAkIY6zlKsrMutmvvRNvG1KtI
NSQTqk3GckkeY6Denkj1YE7tEUa7Bxd0ZeUNhSGfNqm5xkmnpojM8quj4zS9jr5vuC+B9h4TfuCl
fhF5VtagMIiVfwGRVQ6EYFv3w9pFdYidH1HE+ZpYIoozlIuOfRJaT9bvAiv98rG0ZqCC8yxnOV7N
+A+tooEdkgjkVEIP3srB59JesxoV/vFQ/SHfY4jNLcG4mZu7fb2einivzN6z7vy6yJcJUHwAc6wt
8RGtaL2tL9PQLiEvAvQu2wcRsCQ4zOtle0CyWw3KqeCVQD2mOOIv561dNhnjmlOnNL485l0s1A1P
7P1gcNAG1g1KgcRNsfPrUjX0sg3ydnoF26LXLt4KkIf8e/31oGy566xICWb71ivPPYXaUrq7jnP5
4/tNcFu4136C531l2UdKyr/tZo9BE1Qqgb+lm49D67VI1GsNTANyyDi+gIFu0jwxymxfjd8YU2K6
O7TtfPUakhLnum/flX25GReFn3RfDJhFmg6DeYSwp9AZHnpY4uDr32RxJcd2fRWOSXSsolC4xvk7
RYxvmT03yzESyK1aDrEx7udygn+UslpTAnt9Dr7Rp7w9tlQd0o3NnK8p0yRT3eeb66oZhb6qp9xS
Rb9i6+I+9Rpric9QzrECbuiHaLq8P3wR9JeSRgi5J9bttVW3Qso1+CLP8ZlC/cwjrs1aPW9Ec+ml
jh3+dDu4MYVvVz+5q6gy02d0xSAVaPh7o+uORFYJPIq7bWyy2lndDNp/8eMY5DsUEYcA1OS/c4lY
QbcDaqa5JA3T9Fz7htaIKLQLz9eBxFy45sgau3JtMQ0nELRst7QeJMsmjxHjYSeMPW6KkNVeJKs8
mjzuIkLm2QM+/M+h0BbhwgckFNLWkgKFjSVZciakVEzVQG0v4ERZqtPMfbK7dwGZ9Ivjs48498FL
xR3SkOA4qK51NPJFM8RWYWBtH1QShzS3wrPKgUb3JcpIlVZJm5LP8gD9VroZYL1uJ+06B7/3s0z7
ziQzJSMLIEfixLHfnwuvlJH12O7ZI1Axs6IKrFdlhIgMvWoIIf14v+T2z5s5946DVpLSYXZ6NMwf
5ou1ZdNuP8OdC269kxUMDRfDemlFksKRUpGhcOC/vmjrGMljb9QBzImS+sqbUy4PBCqshCzB9OAC
fXNCZoX/c7XoBNJiSzN9z1r9uorPjJ7B46kXLIDmKEW/hye1a94Vc3YFSuhUyEoA22Lb8y7qlI6T
P5G8k92W+phFIoLU4YhSuKEdCi9vLktruH6X/K0upOp4WFVHr/b1Rawvh+3Lv69dMruNIlrnIxze
9uQbObdoS/eCz7mvD8wqEeYbPqRoCj2vb/UvMlAaehT3KbPjFiQrrEcJsiD3NcM8JNngZ2oL8sC/
0iBxMkI6ZLRQ4HPmMzvGaNbbodNGU2oGLyQM5lj4XECv3JRWCt/ESU++0MJglZ2GoAn2uxiSvq1i
EWGR7KVNHWYl8ennq9Ko6skjXX8BGEXbXK12zfkFjCu+xpiSNvCNJtCxKQE+aHZ1Ay1KV9dVt/XF
E6CfWxODNma3AGhAMo2//qbYeGLyPikK7JtMinNbuRZtTLIJhCeOYGLJxToKasE1gucj1otc7EOv
E3ad5+pqkfUL9EfiXkS5AR4ACjV6zAuesMb1EsHrTPJAtMxuVCqar8kz8OKW0J9UIRqfMRf6sFox
ZRqevHHG3es4mbAuZyT0Q5NbForsdT0IsgFnJA7IFW230pbr9gVgt9cJbhKqIjjyKzgtPtoIV8LK
GAwNuzUjej+7lUo49OB2HGYM/ad7kTbfoYrvV2cwIim/fmhAEbz0lrsgJOTXKYDG4LHEIDUd8cAK
p/3J8bEJQld6EKOF0J0S+a3JUIO3qxkHEbx5U/x1eOHuFgxEpKqAQlkgbeqQeQ62kqas1tqQcdHk
SNUMribJEM6stHdCIxliQFnMliu+WxYdGZctqxGzojpqw/U8b9CCIWIWgnVZE2d2pb6SsLsGiu8j
Y52R17DodzPwJ3eq0t87i71wp6hjylu07Ua/D5hizzP2i5LijQQ9CPryAklGHVcPZ8BBy+1SmKhO
t400UeFf0I6f3lx/z/Ovcl3HO4J/HGCDrSs0a9C2uoeX6VCqPLiXQoIHHecn0Xb3+c+Vb5KtfQdf
b2SXFNaQKy0rpnP+AN0RKQ+zTLr5YHlwMV2xdhi0rA4U5MeXAFw40NJJvJhO6L77IdTBiKJbBhbB
uiIGpAl28IcAeqPjF+SiKpbp5wDvqmLeowgMhO7IeevbIDoElhABAmABnJFg1vn6KhE0j5353Le9
LG451ZSdxgfndqL+1mYT3hnHqAotU/xYecEMDbHigIjeZUrwZY5MOXwatv61E8CyglXjQ/EWK1k5
O/M6ms8aFXrC7xflhPtR0o1f1zDWfqI7RKKXAWKzW+yYDrZOKsuottqQ3jEc8iAKPCFjPg6rbBK/
djkWJyKodO9tZOwKy/K4KsNKGm6ZLQmu2DVJHV/jGdlHEGfM6rjebXR4r5Y88Vu1I8cblblP543k
8VLUMUT5sLMI+356FnFQnS9npsS0pfSClweL6YLxO/hsgW315TeXCUOP6CcHgpGgOR6TM7WHXKWi
STYlE+f0Fk0CVuhzVQKmlVngf0f5z6eoMX+U/z15LNTEaQDj3y5AR6Us98AC6vHj0h0+efv2Unc3
umBb0U0karRCw2t7ADpXyhOYDiaFwwXzgwAfxs2fq2vuTBuTfNi02oVNv8iB4y2bseF70anTVK7X
t0AodSmlX7PH0LVrOCNM/pQwKcUKiUwtELF9KbKtj1RXK/4VoqAgH8fY5F1kpMjFWIFGmzdSBbaq
sL7DmR+zWUwQgdnzGuHeGZFeN3VqlQ1zaTUFB+mc7DhUp048LCvrEXP8z1Z2Rig4Bm1NLwUXxdkV
BzmiuBQS4RN6OJn5hXC+Ei9VxY/5t2DgKJETgtHjlJvDr/PF6iYJH9+HSM62US/4onoXwckQliSL
DtR3oQnNRxR0yqF6aXTJPFvvlv7/4pkuSws6MopSrCfgcdUFQ5TJEkwb+PZeJw+4ufBUaYk0LmEl
X4mdyMODedGMQHCNLt0uPEB0RdSs/bb9KtkIxaIGZ4G9CoVo5p7WKTc4lyFtwT1uN/ldoSl/DrPN
407lsJTC5yyNC5oPpolZXj/QnLUoOqziLJY21JC/s9xy+/g3SuVC+0M0KdFVtvWy9N/1QZLWa0s9
jXS7xvCjSuUyg4QZDH4MW17zJxHnr7Q1jo+sjVj0nu1TOUCeqW5MX4gZ38vuClMNQtCf74H8EvkU
+ViuFfm3hZGCLIRjNOJyP68fjnftmG1/4D6gkCOJ5IrO0CxXulv5rQSHkCLbq5BsTsM3R1IbPeJE
rms0VaORz9YWFmTIJsewwR2UdblzPIwKKWWgpXrR4EvBu13GHuhUfU+0+U5222T1BEefXBGg3eA2
3BBemjVLU3fny9Icm6UjpgMyM9pXBVVvk5LxkfUsiLr20Y+wOzbA/ep0FEnYMiOzUuI8stKNLtSh
WKSdholFl9utOfI6rJHQaPwh3Bp5G2naehilTV8AWcLWFnTjn0+eJcQLKgJt2phOwvN6Bp5Hmt81
2t8g4pAkBg1awWzR4ommIj8QurSds1XFINv8kn0OWF2Hn61raQ5Y87Zt/eHqIdWEDu3f50kl1x4H
A6lJ2emeVhiWPQammg3PMRvQ5xFystyY373eMZUpq980nuYjjfrQenzjRN0UQYIBtQfdrEHP2P9f
ndUflQ1VBm69eKoX9/2klHbenFYKN7vw6ta/hR8MyAVjAl6I/22H+xF4sT/2PjVjEHKrXIDTKAYI
J6kKkuzzWl6ie4gqHKj5roUWFeTUuo1XlGSyKinjaSETHcxs171YDGu1kbQXz5VnV/8WUWxxeZdr
8SH+/oYFQmBmCo8zKAzBOPvHQPdobKH2Gunb/3F4JnYkPPlgP8YowZBMktPi+4uLfpJ3bbe+lsSp
JHaqmS/5WfGOkkKf2mziwZUuRmWGbqhD8DKv7f8ZqK3msKaKi3AEbI9rXA0gDYpdmhorF9+Nf/TR
teHF+CXePHrIdnzO/HKmlwQndmjJ+f519WALD4rpUP6o5+5CDg7ZWYKgdppOJ0K6gmWcNb8+cs7x
IPRzYRwvyc8CY2wB5ZFd6K6xzOoUn2fStK9hwIcGAaqUJMZulN5b+qtuT+K3H9dVHhW3S3UShuO7
TGGiC7kL4V0wS116xxty8fyx/a4Tcl7JJnAasN8e3LjSMIXm9J3D2VIEGID7aLOKa1D0zbtnOWu4
q3+aXSe0EVMzzBMSob3FCXbqtu2TP75Bb8gWqlP7jLodo+Fgog+ZLElt/fioc6FfuML1J1xKD6bl
e19ir676H+AajJoqkWMwSypeINSG9icxKdW4Y618AS+APqj4wTaQJIB+lzydySnNx5zaEnttEGZ8
kJe6uoE7mtmvMRKdWIcE+eeuXrUuL2+m1YVha6pX1FxMIADt/yDfNvexFdUidjItWnw1LBVXQ0ZC
nVLEanl+5V9EpqxevQOoEqs/AcULtXRVyTrxe/ZXtDUNW4/UkZa2Yf2myCkFFFrM0ZpumlIMs23b
byYBiHmw/CsDUyXBMF5Sr7Wqth4IAYSjNdZgDHc5ietAypjdvuuuUnVK8hdMNcRO9yBAzPWP1PJq
LIjxDiOVAEP5bSIR0ouiF+ygvitMUn5nQOGbg35ALSUzAXfVtsvk2Cloxq6YYpOvNFr38XDJTFjQ
NdhDyfi4qZOfDIDucc9gj8Kcp7IiSyhBonYFWzal9pEJTUAI+DKQBKKcGwK75sUlUjWi/YW841s8
pEkGkkfAwIGDXxjxr5zVxAVp5OWOdiqXCHdAOj/lLjQeLyjvmsWXFnYjZi6TWA/wwaS6lEV6Xscg
Wv6lsPeu+Kh8j0YEXsN6I9jVz03InndZteLqZCErDjcNoxYGPnrgL5D+sEvZ6ToXu6Qv2ejVyB5h
lGNXC8aJGH6RUp3EmfPuPprOVSFXIK+/6zltyu15eFu2+QojdNNaBclRtmWQ9SZEu3TA0cU2BvHv
cjeMDVMnARq7wJ/0BtN6E5Hwn5jyZC0b0wFNt4LEXP3mHv3Hzi4snxEKa5I2RJpQX2+H4rEmVj6K
EzJO/ewcOm9NYoa8yp86PiVVmJy/fTgs7n79Iy7jNdJsiQ420mGIcfog7/urxPN/Yt5/nXI3k+JR
cEdMjGJM4xW1C5NMn1Kf04cZ5+4YTjTa2FHfmEv1upERylWkoseicAe3UOmPkO77AgSpVpYSpW8C
GrSEQeDgQdbLTQM/AI7cBRUc6aNtWyvByrvd+WUwDPE0PhO1mPf73lBXlq7Ug2ixIrDLAIB4pGWE
a36Ec/o65dCXmB7c+mhqihPcyPNQW1gFMH4b9BvpADSQmhqhYvVzb1tK1VORwUKL+/1/KNY7ZAIz
i1Wp0Dj5GoBF/5phOvIRaLyGBmWp7giwtnOG6rhlG4VPa+lw0iL77qUFM605M/GYw9tuqRja2eVt
5+Rjz5SXPwjUT/k/sxipZcIDdvOlNvvz9k8MR+l3VzfDojwyZLATAsvgjyzo/VKbMLnZRAXAebSX
2RsHiXlmGj9cBrJCokAKXgJ3W5kBGkSwLZSkR7mST2pN6aUEnmwIO9OIYssi0SY5j7LDrGaStfJC
kQUo3Lsx1UNLo0fAyN6JAW+Z0DDk74qESLxAntP0iq7msu5PAC3vOz3A3AAqBq6jRs3POswv769A
hmutWwEkXLaYoy9jqx06vWnO4ntpThzd6KMjGyWHgG49p9y9z3os55w30RM/DxXVdZzwP4ELFbPU
tqHjohq0gOassMaJBDyYd6a7eBdB4rHxDh4LLNNCJ5/A8rnI3JRK7JMUhVE6vA5/4eMDzNY0mKib
foWSDb4FpO5MKlvQizYdz+7+M8N7zwm1Ws7n/AcIH8Ezvllc6KkWiNylvVIRl1jzHEUth/MCUhbb
QtVf1C9Pd801Mlf+YJo6NVBaqiObrRLJ6+eEpWvlfMVYBhV8bFrHssVHUgVQ5Dgq5xHtp+JIqUXd
Tp8hA25x4AMO7/UYInl8rg9caEEfvzARtUvssN0q6Dodt5IiveLXhGeM3roBGFA+zSnP1qXJkSuI
cEMkamLr73cLXRLV/JGYVqOFBY5NAjk+uTpQxJOZ1+K0aDXK3F8JB7B4usIHReuxRMbPvxckcWio
3UoyFlbGpoI25m76ln5xcw3mgb4nbVizfGe4PbWtpGbpSK+S7h4fwQkQ6qgg4zmEUtTg+eUI64KF
CZSXQ2kvcT+japRhJ9n+adb9UixeaqhhM+qH+WivxnCHH60dM3cqj1tvha/PQYuAmDC1nXIRvDcn
12h25xB/G7hYeJ78TO71/yAxweV+g0Zxon/XWqP0cY5696pSkN2WEjNMTSlPXpkn2FrqX2UylL9q
XvfsqQnlp2nYUdSDCFnXq8vivjk9nXhOnM9QI6pQY4vXc643dujURXs5WF1Mh/IwsJApbRjiuVWk
N2124K3W2XSPB0d86uUhqwb1cUDP0U+/JFQu9KOVfYOqzAUZbu100k2ukOF/ZZ/eqAMX3Y52ms3W
zp+e1GQHrX+DQEPPPIPzVSOOq32aEBP+nY8Y4rQc2BfFMPTw1mzE2xEeEt8oW8rInHo3KjB9gCzC
v52u62KaBt1xFhEk2yT//u/S/u7UfS0zMgf5JWSCNoF0+QEWktpaxdgAY0YbftlPTi9Wf26hP+mR
Il7saFETXsNh6CF+9j7Wh2FG0Pm2NgPXaqFN9tQS/lvIpCfVmPiCuRM2/VwHfI7aWWCLFGG1CQYh
90oTRXq0OsHhERc3/1VYDoGEYzZXC1fM/hqc+io7KbA/TnQjINJ0mFRY1jF5wW+EGD8+U3juGaLL
vWWS0GbLrKNlAk/DJKb9AgZFXugrrbeOJPtVFlcZdmzb/8c12O9f2/OLZPmYcfVXC9DHdHHvh4f+
FrjaGuCE/j92WmSr1EpUYI+8v7b/c/ThDXdF3wSzn6FwOYwr1fX+Cc1vvRJMZNo+9si3+1/OjxHg
vQSvjg24fXw9Yw2eDwmGWwo3nCEKBhNadfahHulCTkIqxNSTHmiTLP5IHBKmVDE+bc3tTZmmS9rh
1EHgmy1+geaFAIaFF9QrBp85wg7RwfqzzngzEAYT5TNFoj21aye550ESyGYWWwLtXXNT2MXOs16F
h4rA/Lp4+cYMH6UKEcM/MDQttqKgjYeQK4tC5lSOLuuzCrDIa6BEuQTRrxGf35Gn0pgwHVMhna9p
gxLRI/x3D9/fPeNgc3nIsZGbUXP3dAfC92798Jd3rM11csC/smwQQGJs6M0MV93aPj7CsfY4jHfy
XJoog0WyYLGKIB2jjHDKuSMV8FpESkyjWMcrH4o1pASshVftU0o7WrrGQWMQu9N7D6t/amCdDzug
YGv9zVO3F+XYM5S3d5KdAh31p1f2GK2NpmCPbwbx+UxckIfZ0im1urrmRcRdLG9/AIUMxqIJu2fd
YRcDConuIGKCYW2EyhtIjszs7t80vPFkOiWxfRMFqnYG2Qb6BlAJqDfaTFmtQgqQBXp5gcTNJi/k
4HsJSsYltwuzZOMV772p2kGJv8GnEH9Zvj0hRMOjY5TsEWYMX6X/zZtYOPcgAukWGFLEu0TPCFBl
Ae7STpMch3vSkvjSVCz/AOt2G8Mepya4nBqDZFnTn3+8coKb/wA98GrmBkuE0q4k3UGnkTDJr17x
PacFwOcJzQtdIcuZ9KjeotzRELRdZ7hwZmWM5Oev3K24ONTp5c1CfC2Tp741w7K5WMZ95h5ZcS4e
oylwVV7qqgKUT0xNk9jIpfOF5n7JYCHBZ+0yqt4/os3aRyYZkpgqI0FSiHg6NLE6sryzmMC1qDV5
2RDrD6lxtHnmpu9rVyU12iq7XMwGyCwnVaIWspG2P9aHxF+gCL4MaWQrISVOESTA4ED732izFNw/
iVagUJC809ADijuJWahI33igaQCSeD6z4WI0rtUaRHJ58sZSiuz09GjZ4KppU6QOaXKvCc3B/brp
DbuNB9UnYa2yBiumMEguvq5IjF4eLMFGMcgRp8C/Ym4R6Rdn+uVcByjH/A2pAobN0tCBxhAF+rsS
FByVEAhAObj9iP3Bav54CZN9+8VozEs3Zwg6Uo2pQ0Ix1Da1U9Dp3mjQDw6fqC155VbxcAw0X3Qk
1dgKuvswaJq7V1JDaiE2bvdhpcBGrYcQddmT/2hZ4RPoYSJG2NSMJkuJDTkEv+bfgxU7wuVLKgGe
BPGTaeSG+427CA4HbgG7iPgt3kyXmgWr/AIbvOwdiIwoHXG+EhiNSEcMj9clg4xrnOa9BQl9ICBP
LlvugLV+g81kZLNGZ426V/UWEcydpR7I0rzWQcO/W+AvwsylL62FJzsoOd7YMBoOHppnkmuyV/Tf
jOI4hCTWC0Suly1PEH8WowYQ3ieDVCPKejH2vha56R4/ZJiPtTFokIlKTCnHYRC3+/OYUbFjES57
pFgMAFjKfw+D2aVbmhzbUsyqxDRFasKZX3ZO7a1ht1Oy1OJSr3mYPGTKlXHjEtcXPV92tdepiVMw
4AALTexsyg1LK6LeHWUZD3KbNpIxdmfxY3E3w7qG1ar8CsRuPjr6UUWXV2YWyU4AYXCfey/eVm6v
PmHYIKGuL1b4t0TcnFLECL0xyfos/8dD2HfF+lzKKo/5kkWsFu2IcguY4amG/Q0rykBCTyuCVPP1
3NJSl8PonhS6mdTrczS0QvL07FzXCPp/QlNCIzyjKjWtYY72Iz/SenoCzUgip2r9zj8EigM0PWBe
loP+84klt8LalJTH3ZdVHOry9E807jRnfuy3QNxzS+O16DNT2+VBBq4rucRPvuVpQHQC798lE4wr
A/zsnuczyPYApx8treeA7RN01MkB5xUyfz628Jzre3TxstZaJtL3OurnX+OodVxWpTbovsd9uLgs
x3AaZy8JaOV0KwJvaHNVjONFl3NeZ/4pLoWBSWkJXFH3EERxCNkloXefxR3vCE61FP6QI/xhT+gk
5xKd8eRWepvI29lF+bwxC/tplAP3effZhBhNyeNclSuYPj7MaKFNTmWX1Z702HR/0jnGDtwE5HA7
1FtJakkZZpzsUzR5xiafl9kICrSRSeFB2QTJkBXfrbbLjqibLx32W7Eoj7BFH6JFRoqYk3d6YS5r
u4tkL/AnFb1c7feFyxfyDoFOfNvHSHtRt6Z06AFPCjw9YJbmNmvJ3Z7m3mUCKqg+4LIjYVyi+mxf
GT9B+56T2bZ0iACV94N7ihrSQUL5ZHHHfe9bHg1Oa6sWtNKO8wl2QQ4nYeza6JpZMBwtHRer5kpO
UhbkcuGnEBcDXuDEQEN7onJQgd3B2zG1PnIEgSChwFgumgCDIDy/uGv4nLPhd+m7QygeT4mn4ADy
AhkQPh3371AXWb+CHtaaH0MyjfwqsWdMdh7r4RfdUoph3+mz1qcUKA7CDwenjcu3CY6KD5duGrBX
nz5WLwZstO0OAn5UaceibJOGfrRL4q5JCdXmDY8P8tG7hc7kIYnBUwzEp7u8xgOXbaC5W3bsNbcG
AX1HMrczQ7PHZ+P07XwD25yQr4aa99O6VqAfZOFkwkXJ2voXhl9mCjcdywhO8OC22Okd9QdS05h6
E1fAudhFJG8o9+ZM2Aas6D4UsyE6W6L+HiIu3ezIpTo1rJamCzQMFAikyWLSqhWp5CqAIyGj8ZQw
cXko59CETPj2umcoe9zAiRUOKV0DwxrZI5//wEr21Juj+8JuvrEIEgCsfUiFhZDGKPVepHd6PIGJ
xdFQmk9kqeXQkHdmlMjR7QP74vRLffMstLCxn5useosvgtukP3nXm/Mfz1foCQDCzmO5Cr/xjAyA
2iFj6sMxXIDtphbjGcloerNLq+d3hJcsaq+FSLh/RuX/fQ30e6+rkR0qtEOoi8SpR6LREUfFaMPW
xFTHJM8K2b9dgW3AGmxctDb5NBbLPTtMMR5pazA5gsGYRLhWzpES7ZvtzAo4ohvEedVFH+jDS3X+
FeMfeX1i0F2R04wA8DxnMo3rccaEaQ0QPXE4+4Jdbgbz5/vWg6q+KeHnLhawkhojVDnhFWECqfT+
4FJfyQHlJHuDh8fseVb9tKo52/z5sTSpXyLcSmoEtbkq3ivlJ41gif39UmLZGdotrMxCLtASiOgX
VGjJvsKLtym4G3FZ9Wy93dqm4cyDdm3InvJ2ynIbRhXuzg2byzmRCIRRedjifQVe/qEZ6oKB116b
Ms6fQMYlotMxSwi/MxSkByLcZtpSvv+AMcYDZCYBfB9+I0qztAwePSqTRp4DrZxl3mGvifexG7BV
hcB3tMtbwLggKu+Z5WuwoOPBv6l5ZCDVxOxxTcGLL9vW03IkiR1LlFu6NJqSk1oyy6P7i9AgMqxw
jBoYWpkWxO7MiSKT/p2Fvdo1ANuTJ3xK10kikumVTKW5Ev5gBOZ7ynxFB0TRrSGOQwJPQTd/ZW55
ReuAZjlQK2dpbsPr/xM2n6zIMKGwaoWSgcVnIfPcsHgC56x/Tj3oQ1M8/G78n35nxdZQ3sRxDvvL
w1J80feKr05F6oc/hv8Z35qSqPvs7TXmiYQtgRmBS1EDvGwLGgM+TxUyGRX8NSCvaDDdkW2XNbZ3
H0VQsTiwvPxnJWnRoxtwblXq5GnBIqqWe/89ha4/tb+7f/Is8Oto4vjEQdEImLoYbYdb9etUuqnm
EEnSJ7YiM/ybhYBllGeBkGPdeCR6Re7CuPLbAbbf5zhxEXTVaIAVOswA3axGmmAbmCtKY4mcIXue
JKHes7ywVXAG2U5Z+K5wRU6FtN6Z9hIC+khOTgDbydTVXWIY4or7HvD394SU2My5b/ck8UJieppN
7tj/vb2i4O8vnk8vrDLsXttq8oFkE0tUIJJEPqMpCyCEW8a6gdEFIDMBF+RV7NdT+iwvLEyuV9Bm
+RSEXgvYKYNShfubZ5pM+QitgDU5wObMKhvcSYV/pbQqppYj5Q9ilV1w53ajowREy418UTOWDqGX
snbMjidtEOBkUpLvw2kHWtzAYtjmUv5ru3oQUlJZOP/OSRn+/hfGeB5CIWSRblJ8B8KT5NYqAEW3
BmQPO8nzF117ZDgP6zsvAgLQdAyqC3eaDJq9y/QcCElnictVuU/YkMX9cFe9LjwdquLBR9bgP+oa
h6/aFDiNBZCh89+WmFl2J8qOLJfPBCtegwrs4ZcU6LKzj1WJCTjtGI8XWsQNc7ss46F3GIKJAg9K
tkjc9TXKBosRdyby0v8bsjxZ0Chei8t8gsvtB2Lygdq5xb7nBaR1sVD1tshs4Yo7NfSdybMc1XXl
DIt9KpjT2QbTMdA74myb9eAIhZgX1Babj0gKipWwrgHF72FoTGHVVMJ22FjHk0MU14UiuhnEtV5O
8QyPZK6o6iOJxTHugUyoTW2VQOGYt/3iLfWcz5HdQwqxCwhZj3Q2MpgQf+oXrFne0RTwgIL+DRfN
n0QzAd1+YIyjnagHwX3DY3jWjfjslZuETqby6syrR1Gj7wszqvo1ToO2l2DTiQu7IKchquWsolk9
KXzz+lDrbZuFns7Do0tv+IXaJBKz7N9hWewh/wxsDTVMgivrQTaEc3+uS6M6TsZfinTbmqjGuRVt
EaDo5dezOKXVZPDsm2GDIxo6Eqf/UkrMP53VzzBaiX6b+CsygNQSWZ0Xa6GbP5MmVZI/ol7xyCMd
9JBVomwPYFY0Kaz2U1dRb7le5bCAZkj3aXU6OiSpDKW3Wf3MdiHXN+UneosVD5x0vhR2K8qiFUK4
xdo6foFPBBzQNr1UfEiUNSLEPqNyY3CwOiK9Cqwf4NIEE9q976F42O9FGmcPm2+EsL6YGKEBNy9L
ls0byZ5QdZodFbx5Bj6OCs28edJlwg556Y7r2w2hhLky+nyp94Ukcw0m5qPZPSlfwh5rfzMMbj1n
46to5DIPNiwrD37s6NA3mHSJJxah5ogaM968DESwjpBaj9ZnMK81CqpvWz5ZLzAg0iBwuidA2KKb
U8OeYCJsUOVQJrx9AqUERuOYenPLa9nPDrwnYWFUoCA/xYussrcIJGjBYouy8JYomTdP+l2CVW+K
sn5JrzH+b+gETptR8LeTkTGqqRa40jBey6v4uz23ZqGoaVeTzLs933YTBf+1HoMlJqsVAiu2VdFZ
iXXenCmTHpu9EhozZvwjFJufoLQaVmisFWglu6D9U8QgR+LRssbKAwkqcW9tm78vM5lxWQMojv6D
wHcdv1TKjstMVySdSCCPdLaek+he3xKawyPP6izrxMZTsDWoeEeUFTUOZ4BWwhpRqohoGnqe1clJ
j4mY25xrnB8hAF3ZJkushg6qrEfcFiempJNhCBMzsUSwAqUwEJjW5WIfMkNWaJbhEJzEv7I5I0oE
koQtzX7d5NGZwlXaXpkiywokUESZmQ8+UYfcGkAVRoyPQnkcl+t79Zf9vhgVdJwH0T1vQCuIa6DO
3LLoKV33heVeXxOQ73UH9txesp6hjDP83B0BT3+gY5/czOrTsaqRs8cSyszuEWjr3pV7517aoKQ2
MWHPYelJfU903IV+EFDyXEXJQqM5kmLU15a4fNoOw5auF6AfqUVmjsimAn0dOvh4sib+6XmWwzyn
hJDrgYU+qfG/iKzk6SGb8qT5o6m0tecD5zDrLERu5DuUtWsQGfh0OV4G68bWBYEgDYeIcdMUtzk6
JaeKBLQu28s/0uzkDE3JGANiMFyg5P5I0DMe18Eu8vLcgXgNzTgj0GlKiqllSYpwYD1B70WJ5YH5
ZWp9H4YEzjxu87kPFO8nwo4LjInL84+C6p8Z41k8AfZ1yfA5m35FPCfbQOmhPk7bugSDuFveIGJa
c9gSVEfSWZtViDUBKvdpOTEdDp3bXrJemfn/IpsC0IvifJ/4wJHbAaqUveXMEOsbU4j3YJDIYmdn
+ZPBijHZ/lAkj6Ti2Jbks/lF7hl+s6xHXcO/EzVGr+e9NLyX1k64wktKwgIbGTCQKGgiBfwnCI5S
kGgbgBAP/2apSLJdFyMjDmMucXJyVTzzzmDRmg06dqz6H9tPHItKhckRj8qdbuO6wxAAAOnvlIfk
0qMh5N6mHeEHEjTL3i040YfswLJLW0Vg6IDocpakliylARHqywaKRoFLp8nWNShfRyOfwOCO+n7P
PHWL9UhfHV0A4oYtKXXGB8noEr+ymKVsl6LzYd1Yqfs8J/oBHbEnCNmhTnDD0Wt9GSOC3FFjMelr
lK49yIaBqQD9gu+HEsEoiDrxJI8BLOMqkCy1R09WY7BAHZ6CijgHI78kmuCs1NiOrVz+FA6eeNLd
crrYDf9OZOg66D3bax8i1XKF+l6A48nWSYXkuYhjfSfx+AN+pmUjSgOkBktzZlScmnaBRZJzF2j3
rgBjWRzdseLyO05x8uvvJ2zRBATEX7KLFlU7v04NFUcg17UZayBJXhyHN7/wE8Em99SPSY4qx4sx
g1n3x8ExP+dcQuGcnE4nvDzCgimOwsE/D3+cZdUxJ13bdjtjVfs18PkCHbhAL7KDu65IlwnuRihT
uw2/17mdIbvZ7dcP+iKnpeX668zy5qEj7/amoYsfinyz9e1c0OBjnGq66O8NwlbY34xPqk8I+hvB
zimKdNpRL9x9X8BCWGBsnewHUGQzvRZXxLSGpqzz6l2QvmbysXbLejlYA7Gtr1tGc3LGD99K/Nwf
xkGvDBBCbmCLnPOYe2CB/uIYLXcxhR54EKltCsX/vo6omIeOtSYtrJzoIXERPOxZ1s9GB1uaM4tr
zjVWaKoaIMm3smsRR2CjtY06Shca4s+MAGJXSkNBnuUda6b/UpiJvJgADeIdzNlezpnxXrR4891a
T6f1+DzY4vpZycYlQ+Gd9uqwx8UR91kbMHhBn8n9wLkL9+Udj5j9Rqkp7rewJecZyv8Q2Gea5DNR
hpDf7KMpDW+KsNH1qGrALOWch0luy6pbKtvVMxUCv2IMMrcS3h3U8Av4F5VD7ppNOSZsDQZs1p7b
jppcUVx6pPPwOGYodR8AHPI5hgSYgHY9ZWsKM9dyekH1wC8+92XmP+0qtscATe8upCM6HcPf6zL/
dWi48O+bITxgpmVxVaCaRtP1aA4vbOHms+fDbllzx9aNGw5KRxwPcSF/gtL1NOpRSIKHskijDyXN
KctCq6J9dxrMrVf3cu/4wP+uh1hvsTR54Ms3SK66oI1huyYQF27FLKIe3Wt01vmqRqKllV3OpwHo
6nU6zAcNHMH0m+RDWhr31HyGfo1R3LnQ05lJ3+1WDGzrY0NtrtoNTOEgLG7DtgkW6tvSucQG0Jfr
bTXWkMChiUY/HkjfaqJu+OFJbCWlFe4ljmrgH6nJwI8x34+OSclcTcgeSapfCMRynABowLi9i6sp
BxtSK115THBLDHgUGEw5JxlfFOuCJfEhBxtiWM7w2LMyoMjfNB+jRD2R5IQBWJ8ENRbenfpyziTN
Sbq2rH2QfIS0+pMIB7TtEp+AX/yP2d4zzhMsmQVlJYN7qz5t6/DuKF77nvP+O7Wd3BOZ3qBeCA4h
0I+SPRteENDmrWQslwvPMTI3DQbaDhXGHjPsgzIDlX/SfgAfr/6ycO/ABAKDgfcgH4WI9zDkU3Rz
sMf0YklPU8wZkv32TxwEaPjjFppgcS+g7UOlvHQpRFMXCAYQXlr5XqCsto8LtvMA34oLaHGxv8VP
Zbaod15wTI5a/cPwDMkPz9Ziem7iemTap6vPNZMXK7qLKvseB+diLbPdT13dukw428B2bk3kHLOd
FWrCz2wk5nbnEKT4jMywg8riCSS6DjaN4KRGEck55tHUiyQIKI2lWvLlx/T913orLswt/sx/VoGO
FOxtKQuIZ+EFUQvghowTJZAmTNTxLk+XVvjaebR5Xtft3OcHOTap91ja8jyvZy0QKyvP4au7E7uy
O2GEoDzkOXPIAQih0aivupmG/j05yC1uAx082yznNgUuCXuELa/7IS3loiEeb7BGCeJQcb4FOgAT
0s8WmG0pdY9jlgfQLW8Uk3whDi+9st/C4CufiyEhhwyysma4n2MS2L7MNNfPJ3UKBR81R45PZ4Va
l41VRqmijIjRrzWIJoo8Dh4BGSdUq9fpsdCEJJWu4iLQZzUnl3l0R3peOIqTmb6RljtRqXYygFA4
0tPnMJMAN+j5r4mTcQQmTBYzy0kM3OMHXAawIlsLASX/Sk1D3aOYEhjO1purwCpwT6zas0cHi6vE
FaA7NdZCIDlNlPbM7ECIHGvdyobU3AY+qTIkCGZZM20oUp0amkODmOFoAzVvMT9fTF0MnfHPkEr3
n0Df6raaPYzTY7uMRfGRwcfNSo/fQtWQGEUWknLhfVIh9QpMatrJCexw8jhW3WO70RrJ+HpnI1hW
pIBrxt+gB/d9kIon5+6pO6McwvFY8mCwMhGQlWx1hefoko6dF6zN4HBOGeecNTgtpkchCS0T8pDw
jHuM7hdBmFoN36a/j5rypkc0zkjK67c7wc8uaFBs+niQw5GjYMM057GIXT0epHr9S6Vl3c5FK2h9
audhX8bWDTv0FOJaeDRsx6a0exfvSKZH87BslwWrq6ADmqXqYisU3ukh5N4GkznB5vUgxjZGQXzE
+1xePajVNl8FytWx3+Mj78Nwp1rp8CN0ld72toU/p1KNUgLqxBB6cm6nu9SCXN13+TgCGKGgnm2Q
inYQdRAKeJc8r83G3U4yYVAVo/iU1Qp6+JKh44nfA3bbMSS2Yqshjgo+tUboeHv6m/FVUari75V7
CPIFI/KD2fmypwZUIeL/D5BgxHtL4Wt3OA8EllfOl0az4VrPyJ3GxVg/GXVvQJ+XvribTqb33/fh
wJT1WNTsf1dEyT68IbmxA5dS1hHcWuMcrmxCJkcCrdVFj9b0oucN3K/qkQ9iSloLy4PXKF1d8vRM
dGCCA2RV6wcjT6aOL/wuVunmFH7E8e0i/t6w21BpNzCqJrS1sWj9yZvlnnw6iwJBFHH4dd4xjG1t
6obZy7UnFykFG2swClVGnF+DfT+4VAxtq6giOdm27bPiYyAWl0j8aiA7NbD7IP/Yxf1wUAVDiZeh
wiQl4XeqBt9x5Aubr0+7qsoo0oj3gOXSd3thxh+8s1vRoXV8KdOswg/8fXOqa0WM9XkJ7jVA+qUZ
ntizyxFhnN8OXStrAOhz4mgwrlTYEcwBzgzkyL5d8h0oJCHrFyoo8Lgw2+kjggV0f/9H+ETyxN9d
wG+Jy3sUiLsmv4qW7jCoKv9A0up51zFFGdJ/eIZshgD2bPBQIK82svwAyC9zJS/15pthkdWBG1xG
a3oOJbQ0U/9EqUPCIpmLwT1QbKTjYb+ewESZZJl2pI9WpMpUMbrnwibne19pXV7AEkuFVyKQN0RM
9kN+lziuuFRePk+HswLTl+CqBTDBlYTiQNOZ8ENWR18tc7dV9XknYAhmZ+5sEdvTTtz36qejwarx
fnV1URxa71Z+zXRPuw61i0wmGM0GXCcdxysmEZfpJo4ronqwVhHfP3Kzcyr5yDrNKd341FWMSoo+
DlR6cTET2NakjHUP5lrjy1DdGB9oimYGzCPTtZ5X1j7FnSPyRjgMAr+i9QVXKg2sT35DEbWT0Nev
KbBjBNjOT8ugXD6AGvShXYkv2NamPJw9c7SWi/NOXJQU22N/2j7oGyxtX/Wkh2YVC84b/DxdNQcy
JcquJUmDSiKTTU14wyEmpBE0VSNvK1erlrjOtW8Th8bCMDKZJIMoqydr4jSiCHdFqRQ34za3OBgT
aXZnsFvkRRfSzLE+a4varkjcq8NDSpC8mUsKLGfconNWrUdrTOxat5J0rN4sQwp/G7LaCDCkEr/X
i/o9L/NW664p54dNVaQoMGhQ9nIvW3HKtTaj6OFB+HxemRQ7fHPBLwtyuLUbtEtNtlGNizofGTaO
ssUZ2cdnUJ8rPsRHUMWl5re88qCaQlNx89azEIx4V5F5Pc7GoY5O0LKZMW5XeqKzSf43PVBd9rNP
gsXaoNG5fxLKUu3Ds04TXqtAWVQiQL+kNqigMHgIkwC803MPk40zHPL5Ys6/zR+OidIXSW4G4UG0
y3uUVvwafSeQ36Vyol28Ld10xt2dfMGCJRM47bGBKmp4CEc0kJGpPvwexqDDVvp3zI3lr6uc88Ey
bjWAck6niMHShVumQmfqpS9I5wFDmnCpP33XjbV09CtFMiu9D5ydjBQ40A4m5V9ImT9Rk00OuO+C
HCGdW16EN5szI+K5XLK+jT+YZgYigQWUIPAj/1SjP9i4LhPTwi+pt0wyv8ZFgBh7GH3BrYrdJ8iC
W7TaKfiTW3zjs5UzCRA8XW4elOvF2GJ88kh9TgyVwDy0172Mohvo8rj97Y5tsDuECixhlTRqp5cw
2KrutJtxRAdYfkTd+ZCZopeuDlmqVDsXpnjlUkqMsudzDngTvdUmCaPWk7Bd2TV2QySMzgFArYS7
CdM2WUa8+jTiK68VW4yu6YyZe6c5AuIytmGVR/QhxDAg6VInn4JFF2ElY5MzxOA8DY9hDWE030Wy
B8gXhyEkVERBNBVXI47q/ZEb7PW/LQXCgvsTbiC/6AfbFk6Q5SrSBbBWGOGTgaKtOAmOY8YtZ8wF
/mHcHARKuv6RPgfgZi6YqNa9gI3dAY6gJVbbU3XcbzzGGnIOIK9wEdbBxMgoMusQa0eUt2ET2HWi
K0YbozQ8ZHfcqZic3u+LLRNSTwskAuGScZz6G6SpXb402KSwhk3EQ3RnYGYCxRPAG4T//5t/lnKY
WyZxSHokesxdbX4xtPGwYROEpCec31mDZGstw0n5z9F0KKDEQjRx6Y0JZlDX3IpfiXvhFX4hsy4z
x1QeI6qsbsxMbCrISqIlv08O3mfPfZ1DZl1xGNONQxrOGGCAXxBELE2sIRw7VTAIkYJf9bsTbXQO
o1vKtaqIipo0s9yvL3+JkWu1sZ+9nI4gdyg9cfnvv4aJrpxGZrXtXfPUdQ6GIFpX5z6tS/FEhrI7
/iLRRv2PdEfqG5VfHxAmRJLjsp08C+vkduE4l+j5PNS6x5Q7yZqkH/KPrs/1zqX27aabPiBn+1z7
wdHmfBuPO4B+b6obdkJLFjuQ4MFja+Ua0vSB1jIRNAbGHSjw+xOTmZ/S3YIhssHIUWSrMZXbvTlF
FVJ3baC6fEzsG7CuZsJUOS3F7Ns3pqBm3u7dB2344SY5H+L46IVanSkEnOTZLvSa5ZIQN4yB8L0U
V5eWLuOF9aXZGgexxKEwQdcXOtuMY9w6fCBO3WAzcKbYcIteffvBkLK80oYlhRwgGX5O8mYio5Ix
qGXgMO+Ljwye3m0szcd8jLdGslpbrmgCytz+eLkt+8weXFPnGgcFpOh+hsRi/5bgnLNqCoQZU1fK
apB+vz0fwF5ZdugTWMc7NP7F0kLXN4sDQpE0tDfferC+XDIhApc3PUNFspri0pNrEMo0v+rcjRy5
1L4YiFqRTLWslCJfP7PSUoj+o+dPK7oE7dTY/VsWjrBHRWPHrCw3yNNNt8/nInFlcycTWXCEIqaZ
kfn20s8DCJgR4I/dunnucVaXace2pKC+UtDGETU/Q9KPxQHKEqO1rRwjAsMfXpz3pPTmsUy7SywH
L7jIK552/ZwBkbWd8vz95t6LNnmTFswEGNoQiRJIzupftugM5oPsydT9ALuBYClt69vDH571Ehj7
BbmKg9J+aFsJpShFiA2O/4EUMJqNBp7f75JViyjtN+bPwg19oCYXiutc2lbF2CSw4/0l4SL/LRQ5
nkrKbRXOwfYimgD09fXrWEkqoMIxHaYBgGgFm3O15jKapgdyZbfTp1j0f3hSII01fJZkzKxWkbF0
PeinoHHH/GzyUPRbIRxoPQTUwkN8CJy+89Irsz6FPukoijpABXjulC7FDXrWiKPVIBfMRmKi21rg
h3PSKWZUxr5rtisANL9jd/HB/Ex6ckZAm7QTCTJK+DQqZ9vqgm6MEq58MzP6HS6vSRka9bOKtXHX
RYiKxHpAKYR/xNFbQ+YM6E+RMDMI9zIkCo8qBLzZY5QX5AOMfL/jHLFaTrxR3Et5eQUkRgqA8R+e
LvmauaOxElgP6c7kbUdjael8J2PnMy47DkkpbaWDPuVGexrcqSRGjrccP/PW7Fbpt2PcS816B29t
kCj/JqSEWX9rb8BDvzwCWLiHm8iNiLOIPdX9LFJAZqoPeald/Sw8s/DNry4qmF3iaTnHoJIlBTov
S7EZ+Ig0hwMfzYiPOWBiurV81c5govVY3q5SHPRgirXB36tns0Gtt30uKiUsnpFsnnuTOD5TDwCz
Rmsdp6ww7XzglvMQLI1kn3lQ7nsn7RSbxTRBZHA94fr1x6bp59Qt70fhR0tYJzdnci//eW4OkLMs
9oJznwGR9zwdxlJ3FZWf8wx0KqyphzGfzOR96+2UvRJy3ZXxxpWoXM3lmH6mKoYJrkzhih5Kl/IB
EeJ46vzypvjMPz9MUZNPLiFEHGmPrYd60T0MZC4Cy4mTV2dHr5gMPJYIrqEdFqX4KRK0Lg+8YO7A
aVn696zrB0vQOvxhdffawHvkv9SPMYibFuROFsy6zUw4goeWv6BpuRmNcfWmEMGu3jvtra0uGB/Q
fRMOCsRcGKK1wNEho2ibRq/NhvGQoR+eeIXOit2pu6gsx6VKNQjfd2/KZ50oCazTky/64Z2+H/WT
dRz+46V+BkC7/Wo+sRu39C6FkthqudWfNfQLmxIAC32tPCQnYfwLLAgvd38pQzzs967+F5wIrDea
79/D9K0Kbvjc/LmLco/hW67C+6bOc+Z8Jo5YfW17xL3C63E27Ib0E1++P3MHTeYLZSX5T1LxbBuW
CdGcqdn9I5gHz1sah7MI0+DhTmVW4vZBoHhAoBePbvq64ey2LqMcfJYL0O7Ms9IeHsADvMHGiep2
Tqr4moTqWl01QUq0XaBLpxWE0RjkFZ2CH5GAMY0MEe4WYR6h41e40McX4I+7ZhmEONCi9/e0A2//
y3rjpzZNiV9ceXk4aVd3gonQDF/wEzWQhRwiWKCmNMxXPMiMqAeyt4Y+BMp3Tly2osnG00KKxK8x
wi+NFnZOzaMo+UuZojrcRx1CRZOhXy0w4Cr6DTjL2OJRUVWQ83wlLaZaq2f8cS+S3McvVUWCUIIk
lU/z1MSJaUTKoVIi0SzMWmwxXLjAGf/YqBJnkKG6jcCAWbRaHhP3gRM7BvFRRd+kvapX/p2Lp77s
wG3HwlFc3C7R5mVqDrD3hC4Ii5O41CBqOHYfIdx3scUxkzv+o2RTCTMfxABmMRxCGIkVmnoivB2y
ZSjBKfjxHq78a04xdA1UFdHbPC0Ch6jXW/ihU3dIWo8DBsPtEphEnMPZXPZcapO/DWg985X2WW3w
rg7zMNgsGgBDxnOUrhKdFtJG/aFPUG5zfChSqQ223zIz7ainh8oYo0Tr1CbXl+jQxrEgtuK71AMl
joLHzccFaYTLMFy/7kdT/39XDBPmDpgtIysdmFZadocgRWoDltZXKWsouyA7uInxJyn+4ojCEjan
9Ia69TVch6A7ChF7ePf1AaCmYWpv1vmeHCKL++DIX+vi4jRCXnmKfeSpNgYTXLGB/UvWiiTVXHG/
dHXWTlJVu+sQ3+mVYBPmgEBC5h5KwlNY5QBT8wioPqBcw5tyy8u8dlW7Do+wpjO2INbILI4kzyEL
g04+M2fCeo1mlOmZytXA2dd3ieFDDVsAt6VG8XrIHABm/x7qnYckgaf2Z7Jy5TDm19TFpLfoVcEo
IW5VhRPD8ihtKVNcudgjEBhJ5X5JShEESuKH8BhGqWWQZbmOlFoiidI/h68uIUO32hC2T6kBmbI3
l2jmjk2VroDsOU8lpmJ0ZkZ5zb2TVuxU8PE3DA6HmL15pkqo1zm6AwF+PdWlGUh9agvqOKVRnwAc
CFtZsdiISSATfDpJEegngROwAIvkBPwcHKCjXMPr/yYmBMbH8sig0GSF1cIRep/jtlb0VyQS3sT8
IKkHpyuYe9mGQ0ZVPwRk4lWm+VK0DG8jmAQQfkDkzKm3L2FSLKT0A9ZhFyKrxK37LguugJaM/h3W
aFBK9W88emSiTukiLnu6d2YR/WCUtSppxS350A0oTaL+JW1HGoBBjSX+u76fNztkkPAPad7LihBm
ZkHc3y1FpJrIvaA9hCMoiY6xHZQa0ZcWYPb0+vu5Nx1nDb7A2UTEFrZw9+0J/a8RrQfb7QYHnwGO
DjinKycCXqMQxNJJmSv3UPCt0P+GaVc7TOl45xh7UFZQyiY2aMHPJB6fMsbn0Kbgt40r7W4eBDDW
+UYAz+dtM2xvhWDLqziQ90G9CKJHDBVAO7W2ZhdgsUXieHeHB7Ya3sr6h2nGy1zTQzm0cmFOIkAL
XZGUIoi14dIRCEftRAQekZZS4ctmE+y+o+5AI8ef0JcB1laF1A0aG/vwnUxZwUqh7hrOP3tZf17X
hnQJ5wKIBlfSRM/aOnuo0sM+3MmN7/P3Z6/5fqCQJhVhNkaUmbNWJyTn90K6x7f24cbSV74HYMRp
fzHBjlJQA5JLUT8F2pd/qX8HASwMQXsgzY3rsl9La0N1iybpEXWrDtg4MhFgHHAgXpJ0m3LTFmnS
TBTsB+usyuaAgy8Wu1YYit/EHI7po/nj7B6Wmw+XBgVp4lh85+KGytEhZVJlmaxL+10J3hRWU49o
NMZRqR3Z23ecj1kbTnIdsAz0uAO5EIIuhcqRryY0bFOFtB9oK2zR8jV8ehn+1FH/GhT8kYQ2ugwV
MNaU8mM7+wlcSA+xM6R9WXxBYexFG93fIhfPqF6Fwr6BiwxgulgtCbuT0NJ1AWFus3kjRYHCgHz1
H4GBvPWdghNkREPL68MWERD8bzeIJ1War/lKX/hRsWbzU52gQKuFqm47a6R2T9pr/rbZYsaZazbw
z8sR2tPRIPCk1GO6GIYaYAmGinXWmIldffGEQVwkhGqPYM4zxi0d6YrMYbeQW6hstH2hyrJfAgxA
JAzywSJVh6Ii2bfpcbri327w1zByjAHFCbEEOGPduc4DaBszqOLquSnSKY/emaST131jPvgB/oUK
dnHVfu1uEQFyYa3CfyCb5oQw56pzGCk92Ovdp7/jisyifADLlS11Kop//CxZWT2/LTvwcVpCec5G
pGqMPJqqxV19pHooB67p5sBwYrKQFWgLryiJHN/xo9ECgxgQhDyf0JMZISu3B//zDvnMgGta6KT2
u/cdTABBTiGVry0+LREvu5sObi9sjE5GBathuLcXqLLeqI0EebCz55LM0qM8grI8I/mtyKyLljdq
z72HNAGzvpwS9SlqHfcVY/2WyGleAJwjKZVpFvmVNjSwp+wzKUxE6ndOUSw73ADSixk8nO8CnKJ8
rA5yHVT+AE7KhrcBnGhGLkwtc96GRIgPO+Qj/eHVSQCiMieiFBPylhYDnZrs1JB+TQ5F+4DlCi3R
s5XqEwGKUH7eYsysUKMm6yF1wqrY/4upuyiIUsNDn596QD5/q1HQ+YCcHfgqoUTfVvKNJZdTphWI
nlgPKKwU0EOT830typDM2ZH5XoqaD9YDVl6OZ0hm1UQdQrWxRFqMo0P9wlrguWR4pXmQUOXpvVNL
ZVUtP7IYL2IsOpwUzj9lLVidQOrinEc4sUhkaqkLEG/vW0aP/Le4DldL/8zkufCvaiiAldn83KjO
3LZyUQE3icSJfLNEJUaNR05zhoXmSCJSkgni/0EJpsQ0jMljVPj9HNDjrE+5mQQf+Tb9J3xlKoew
0fr23hst//s9adSMPjdqg4foCcHqq+l0LmomAwp0+TT1bN0+9nrcGOBWNHtsLnbuhVzWnIzkkO06
2XxbFfMa39dmjZWyTa4niYHwxYSmTK5MpXEjcj96YCg3HLmU36ZCNzpfqfEdpOpYL3t9iMXuuLa3
J+no7RGRtc4a1TuVaTGbOOVIdj6dpOcSnrhSUK9PB44SpjmW2n66JV7Y/izNyNf6+Zf14hKtvSNy
SZMWU+5VhXSoz9WS6Rw07fBa1riLoBbzMyOafrPZgkiZmk5LXE572p8GU6elXtTzXVIyDWTFTvhL
gS3jPPhuWjCR21u0iuwQLuxKimJ8DkvZiGr8WUPdxHgjUtR+pxWdC+Tj2Lmt9Ga2Zrjcd5WAuJcA
isy47Ac9HO6L/WL3INE4B53rJ/KQFR5g3DQb2vNZUZ+IP17uJTsEoVCrTB2RVq+2vu42UHTbhLnX
S1q/avFv/U+rJuAsoUSuUiTlE0dxgKcptAAbRgYZVHm/i+DX40h+alUKcl4+PrBnlBK0DF9IPYqH
41rGEQU4gTpEZxsFNpJkEw7ijVisyi/4Griuv5KHh0/fuVxzqFnkIhRUGQrYHjB8/I1pWOOTsnlI
jDcauUGAd8MJJiM09p2bhh4Uwyw0XU9UmbidKhpNG7n3egunQFu1Oj6OmSAyS6LRF8Xo3LlZns06
6QYKNM3AFUxA6hNXRakTTIIMWo2OXE+mlg9+hSjEu8NG6cD03qrHEvfwzKwughKTjZF5GsKoq8CM
td3VjvLwr9yqR7naBS8Yt37MChDFgpMIx98uccPL66z7ssimn2yHXrunbomsgzMNtsh3vUJtwFfe
m0RO9O6v0pMLRFw1/FKn/Tr583Uh1+b04FSuO5vYkcT7103e459FSL6VO3kdtK+5GXEd714XlRGd
Bk8YaMTIiG9USAlF6o0PcD9LBEF3ibPVOBHDvPoeulsBPoujbu7lNdXfKkfjntC4VRpB0YlNZX1b
8vMCFGT++4pF5Fr1Dxp0YhNdQVkz3mxDwRwM2eNl2tRaB9+iYxwdxX5rBiv0cnpsBM1ejscVrhLE
GFI884IHBeOywFzg0fsPr5DztK/mO9216orlZp31WUX8Ak0IseN6Ddj0tPjFisQYLQ7X3ghJNk/0
dFDHjh/T0g+GeLIo1MR0WfIXp8JadUulthOA1ieb2c7svZ5p1+nd0C74MZOcd6nRnAmlr3RoxRHm
FDqitjfxp10juO9c4uHw0XoNdwhiKfSF9xsqmGJsszP8wCdsS8A+AuRvsZ2OTtsPWM+ZjZ7vziW3
t9uRQoqu49ubRW/s2Rifb8ani1YiCJPB2QfKR+v8VgpWqxapygpZSvmh6AWfoduVbu34dQGi+T4e
zC+TzyY5i+idHI4Ig91ppxN35gqwTTbxWAHPhHH7hmUsY337u8BTmK6RUq7HqhvQncaA1N+0XEc5
cb9XqTcbYCii2I6ZNdBKxYp0lhCopDPsnn+9oUM3OvlXo2Tq5HmrX7V6lyROc2lAG6Bh9dtGDM3y
zb5i6B+Dtddq1USb1k8cWdDnlb7WeckSrUT/3hvKvmM+X0GIOp/uT3MvTATZGnU24uC6R0UELgKG
TvuMRtd/7NTKRGHIJMtRmH+D/O9bPV/rFcpjojc0xyKVclZyYAgQ/KgSkmD757dUcorV4x4z2hCi
kNDiyubYqhgaKxvmqscmO1Uwq6OoFKOF2Py9P8DZV1yeINQ/63ZEhM6LVDbB982n4kqMRnB+SdLS
uUjvW3CvkGBYgQmh6dGRMsmwVueFev2u3KOvAj0qnjQX4Nf4s6AoMUPakY7C1XFOZJgd6ZMVbEuN
dPiIsjDMC/bpfh5sGh9CJyUnEzt7NqzyQE5YrmFiQYgmSZMSd1hK/h89xNhrLRjYASKapeD91j6I
+IbsXaBWYU9ZN04WMG0DKiKdzZgXhq233FGsGe2gQDRrws4ZVrkDThVYAjoxiuJtOMxX3/yxbuKM
9Kt/+bNVVcXtHqxFtCcvQM1ELjxdN8Jqxpg8+irOo7DkTPUOHyYUiifHxUDWiemuDOFrR5pOGl+6
wCCvhxRmfaQGAPtsGEw5XphI/bJ3mjzhhZsK1LlRk7znFwkKjoszuwRT1DsiKJZVmmt1rMk8k2DZ
8e+LcgIjCQ83sZ8+Dcvw4vNRPPbk2oB8AGrsKm0GqCqoLMnEOexlnSPJBeIZI/MmtV2M0Rui/BYs
OSPPxAH7fwrB8ADg+L7weSXDFCXIaKvtW8+6bT7XzNrc18SoU2LAVOQ1+bwm7mpWxcUpRzo72Ydg
wICGpcbVpKlMuj0B7f89ORVFruu2L6SZBGnfIrj2EL6gAGzXTQv1q362to76o8ibGpLOXRH4zWe+
jqaC+aM0boyNpbUnU+GkFBDXiWhq8QXALb0RpoXHf1OXizQjo1py5GA120JnUt70Rjl7voc/8GtJ
PHFi4isgdkQ6xoDMogry7zdR1QxIMNNhvQVJw2n6+nywJ4/kE7/HwKTQLVluGQjDkUXtLNjvztb+
52GpcgTJS6l93bQxo7qAEv5ZNc5nuG8hRXmRW7MCRsj+193MgxLLb7Qe2HACqOuMsmA7hM+c3nSC
O9xicefHuGS3/V/0hX0a7iu+k1k6Oid23Of4iIfnegfxpuJ3hH+LNJOoyQCxv+rWiQtVOvyMcBLT
wuRiIySqBHmQ2nY4HnKDUOFZZxGH0DOanhMRLcaWBk3wJ9DcU71lZCKKzjuYnsRxHZCoE3vkZXOb
A2P9rbIWkDc7Wy5AbnUYTNQj44a25YU2N9qE71N83Ef2Rk+LoHV72Wo2qzCxUCsVr6eOS1p1k5tD
9oR6VinqWElZoankAt/TBNSGHicMrKu69VGqssqwzWsVHLE+9l2JQ+emG/uVlgedBvwA48CkJx7g
9WepbtLch4VIZcOxcdlDlxEekEBS+H1wMNohOH2mvzjEO2wLwV4OPDPEmb97Xg03HwVH/kdyRB+w
3iBdnmGYgZoGJhlyJyHFEzbXxgqB/AWMYuPHE8wPAZ16874kHoNYD7adwHbk16CP5Uld7R0HAQMV
El5Kj/iAkZDRm6bz3Hn8XrzrtVppqmOwHbV6bVDyfOiBGsbrcul0e2lzZtDZ+nun7lIEttME5irx
ZMz7wPo8OhNoKXoLpOAzq3yqFcM4lmCMkOIAdmI9M76WkaykxeheBFGesfVRMkUNXZ4J0kYRTtiv
TFx7Wi10hQLMl99ur1gM2ym3j8lVfh7VMf9ek6Z3LgQCExYW3A31INmY2e6opa+r0EORBvLAUy40
5xFeuKxtXfF6+dTAgA5kEBHvfCPjfH+ds2Kba25FKgUqCdf1+K/Bx1uCI6oC17y/0jZB7WoCcKnm
U69ptWEoAIrUvWG0I9hbXyAolJSabmmyDZubhnS5UHlUQeMu2ZVASB163/l77G89BIjDmH2pqpR1
tNquF5n8n4C5OF9XZkvGs12uHp1/p0Y2Jr7wBjoQlspVNx+21UcojNiW6N/GftQkHJqU/NyuHy0L
wlr8n+tSf5eva4p1dSP+egyACfwar4SZwl0vmwKTlVoKPGR5DStt7cOeEywWmKiXxhnbzEeIfxW/
rryYCStTBrRHy8zSN9MLFa3LBbq+1VX5b8qcGb10M+PGYXnU2G5wW0jFz2bWHrbBC2OcpDsdW+Ot
covXQgTfVVEZuThiXQqBlcVnmZI3N5zpOP4UL8bxE0ezJCDW5Yuxd9XKKEem7Lm/74CkgWMRwGX1
/IseohrEO1O1WGn/RiqT26wKjAzt67OyH3hqjlcPYwxwXjpASJMO10D+ksOoldVF5ZJFAiIyquRT
RSMDSZeCkX0TmTloVUV+EBkrtjYRPA6djJGkoSEARFifRIJOUZ4vlP1DSzLOmZrU9/7cEj6Vwci0
+jDp7l0b9lpzWAOiWFFWNz5OXd80Bqqg+9wEIme6IcI7sH2n4rjsjajAc0DC7DyPa+8R6+IDJ7bN
okExZa40naIlSMX3GXgxkBEpwUA6nWrE2WZyJQTz93ftB4OXyJMy/p8nhbKYojiL2pHJs0iJGeOP
NMuV8m7Wc984iICopEmkUwJM8LLa0/lllu8qQqosDqFaUP7RRZSC/3ZYkTNtLWnQeAkxP4xxFuOO
Bh+85+kLl92amCTY3ap7Ygnazf4U1sn1sxhtI5gmgkysIt2X6BrrJKHmAEsX+BRyu3IgL9LDQjIf
4WnN89zISKwXe4jZNxCgOqaZV+RrwIzAALEaDa7kcDiI0IMAaF5ee7VYxvmOmlmCj4s2MzVmmkzR
HSm7zmYpYYpIV7qjyUY5TsfbLH+WS/19X5S508CvuksdQkPBw0UhJKEj7QvzpXe4H2CvqDHbmQKH
yjmXABxmPNgQPIXuxAytms9hFyzvKLmQ6JVen2eEwH/ZpC+5+oez2kltLYu+FX/odSx+cZarGQwI
rmATPOddQsaP0t9nP2M6MSWu5taTF19n6PigYUvviNHF22mdN8Cxz6IFzCKTp4yAoBRR1jNtpqJi
RyvQwrDyjptJb0wWytpYQXd2BZvsLUL3bVUKfVN2JWdhcWTZ0YJdms0vAWYFqEzz+ibsIInY3qrI
RtA/hMEby8qfPEN+IFtjd77sAKTRLjFG5z3niKRu+R073qTjo/CbUm4DaU1kZbWiYkzMyJf70t9U
olED2/oEAQRRoQ604rp7heztgw3WkA65Z6GrxUSv2/5i/64Y1s6H2U5DL1cvLCAX5htYEHNbS+O9
HGh0CVZExU9lZKLcB/FGX5IuR8MwB8liKTqF9bU41V585QNlPsBq3CxhA+9ozsbd5gcC3x4Ne8B6
rE0WzNeHolfRdQpiXaSbP5Vnv0pX/pItX5kM5IfowkAEWo3gw803NNH5CrSQeg6jeGPndH4BSka0
w4sEYfTnyvePyPSKmemYBfSqSvXZbcyiZTiWHtgrRWzgaTUcESVEIZCbtlm6EhpybG+1c8mrFu0n
q5GxR7z3U7LOMMx9wOi4Qgl4AjYdoQ7dh9lQgHEXpVP2MyMqHOyQHCutzZj+C5t7OhK4ZlMVjQrn
kSYeVhPNWE/oRmGKqXb0VfW8t+vIYMipdFSyZodS0yLQM1CwSgwFQzJbtHDhJD7LLOkxBeX84ZE4
MjmsGJQaPSs7myBqUS8ISO9HR2k8Hq8epG7X3JV+EPU5ii0DDoin9N2honIVZVzCPaovZRvsZmsZ
i+ZmDXFlsu6rkCTSTh67utsN0EUqObqO/NcnP56gkWFb8RBXHsgePsARec8oo21DdcyMRYQ8e7br
yuOAzYmaTQofKEj9x+8HwPMTCVGSv7xi7fkm5dpzyIK89OfgTKC+yac9XZyKgIWCNW2GiWJqkneV
++BruwaGp++fy1S7mu9HAcCyt8QIOUZ3F1gNiwrsjB9Yd9Bjuwcp1goobVQ6DIJzkCbtmsHubDGE
+hVJejYoDz5PsQoQU+rTyROK/f4fU34kDlrpmYK+P7ZQBKAnDMn0JG1GdtGJJhX7IIJ0uW2lAwy0
H6eBdV54g2mj9w9Xtf4NvSRVJ41HoxtVmXHFHRz+4EThuiJSSqC27ZfbUrsy+ujr8epep36UT7cm
ZnrTVeFgOpGY7zSNzU2UoR3MZb02LxTK5HVM3R0KMgkacZNKkE4I2oT0plcvUnJ5A4GosCPFnMa/
FRitKlemrLeAxWU1TIbfh3AJLMpXfdnywLRLpOlYS/bOWVgC8+Ik/hLlkQOYcdWyg3WTy8VtUjcF
kAP2hsV5GXXavyapyXDydprn1xPJmggG56VNHb9parGQdPBXHEahaCazALcIfumY42NuXfY0B7hl
ybadC7ZyAge9G47QxXF+49+Q6ZfMQnKIcx1aBEIfFZ2IytseP7jiOgAtgozEeRQFnj5aPg8fS+KF
wJaWCWVowNN91m+sfDHoqiulp2DIzaLUgXSisXNN4lq/FpD05i78LvaZpw0nXYpFjx3CEcZvFof1
bAFznjLpi1RG4JfL6036m87HbE4m6qedW9Sn50/DZ8Iz+veMOKET/PYc30uFKsJCxhlpdRdQKoxj
+TS4u3Fqpb7Rmg1xxuA+HzsEiRLwcOQQqzZYKP5ct3vPB/+p/7Tccy0cWRx0IH5VM2V0qOy2EI+V
55IL+j9gNTPY4U3htxvhc4k2h7l7P+gZy1CU43LClyYD9oaRF6tpcwgCFvSHtop6098B26dPUTh7
Ev4TqTAnyrIUrELCx57IJQt4sdihDJd3OFPrWcM0YAXuu3esqztc/w+GTO9j8gFXIFF/hSu1hsfa
UtM4lg0EJvyVL26rHWBLghxSCosBJU2DyJC5DAkHzIhtKruy094PG2XnHMe5HOsSobtJVFLdMxCV
+eylmd/cX+53Fazrz3yi4ouBEKTZsgXP6qhKtRB2iG8vDOcYe7dU+6nRQodgx6Bk0NoR1nsCr5tO
1m4W2h6rqDVK73wxKVCVrl3tyot+6fPvhcqxPXvEdH1RAgdUndLar4HE75g0W9nRBiS7I06Q/3b9
HPgPPl9CHDOPf/EY2n61/SQhG47oFgIJE2gOYU2+ffVK4NeKPVGYDYBGopo5GUmmO2QMWZZRBrkX
+GNJV1+mVlcJDFi8w9YzAfjcj6+/BhqLdzxJ9Ei8pt/JQ+Db80b4Fl1AYfGj3lRVNP7jTxetKW8Y
NUgseABTuwIFtTrzs8YxcD9LodXOcTh1WFsL4ZYyjS3FPCDGl1nMgv0dg87phyQ0GhZpkbLaqj5T
PJmsl3gGzZKSI6kuvcWq9zW9DjnQaWm3Q6OL/6EOlljX1kcquJ6d7VzPz1z7G9xtzeo3/b6wBQvl
F8sz/x/gB1IKzfnjqdhoyb+Bnfx7nWzmfXM11+XRvhX7cpt2MfIkHS3r31u8Sd7vDiWaPxyT6Nhj
e/vJGlc5eb70oPZt1SjEoUm4nVN4IIwvyiVYIpKmaLNgci7eQf0HJhTV5bvFhnHRWeGwNavaoFnf
qSozO7y4FA/ndf2/vF5qjPpEBYxDXnQhezEa0yK7DOGtvZgQSxMIRmQE8psd5lEbhxjECHXQwSUj
kpEoSD4VxpFF0j/Fsud68SfBgQKAO4rw+riXUHRW+vii0bGoqoTK3p3OoiTI+TSdva23vwDDRs3W
2y6BNGacm4WdHxpMVjJCBh6cET4emh8fCSKnvsyzQ9DQwNitLVMFeegZI9MM/5aX5GW+rQLOi+hj
qm2yQvP1FMoRgMej98MnDHcFwCk0F3/1CWpXe8RHnRlV0VLAgTAMmKZ4Hov5IuN84aZqekNFpamo
0Sm+Ax/JJ3+sY6TfF6xHQb2IIX+Ynj/ld6iiGy26xxdLHHh2IF9zfCZEXa5XFPPWgGYrNhM9WuNi
cD6vIDn3CaXnzhfd9ShC3ADY61AcjovvoDT0MDQW1dCHp/tPyX+gIgSKswGyg48xhYmBC6sD1TZV
QkmFHbQDPRyMVO6BMbVi5BGQ9cFfybxmMdnYSXGhi4kyMDx7YpcjI7YvR2qXCoRIlMTIYEs0PrP8
hYZLXbTnAO6L2q8bwryWqFxKW2dkghKPo1FtIUgcVf4nMSq7dUkOSTCtWqhLHoJN+fMbbKs5vycj
iHHdQidB2n4oI07heXk0eqIRYkZlpCsVSvuG9+eDGh6jDESBwf7Lqm1IhgCmVV9TRIA+8OMIF8GF
7pdE0IA/qpWXixwZU6+kiUbqxocz9ISHXwmpROFnIifXFkweAvAJXlqN5tok+IOrsiu7q/OzbhqO
/UbJqB54HR1QbdGXDy786DxVQMrlv+K0z0lYeipVIIsH3AhoIZaOb/dof5gVngyhBC2UqEK9/NWk
ZcAphcN/KRicDnqMYbDm0qfiX8j5qIMs/i6aYMVz5FdZxoFUHf17NJ4xJNdNUV5HLyprMDO1JHJb
jywc4c/qbIuqGZfCgwz47qEZxCDpRs4ndijCHeRwmS1oqj9UKPIfRqNdeJz2fzXH0kte5mxr/7kz
z9d1Td6KYbnipmoUm1k2A8k+mAZqQLkyEz2VLtVZ2Y8/59H5POzRf7GXOpfTC4nTgp98PtRK3JE9
0CXYmBxiiG/ipNjPaEQtM6M9ExzX/8eCiaN5lA39jgI9U414JO2x68Vxl3uX4MoIAMkWJ9jR86UP
ePK6FQkib1pn01ssBHNB7mN+clb2JJoYfHa11myNj3FwiMGTkzQbRE4mZIHScv/X1TP/lsgfgRLg
LtRAcZyU1eaHgohFavRkltk8cQZxsf9puKvs6tRrVUtBGB+HhYTf6zhfAqiODE7vvV9EBia+GZmf
6EaYEVbEGPZ16PxSGLyiOFaCM3gTz2TRrXRb1vQ7GA0oBAODd+1nB5xlPpTMieFgWiLmlsAISvJP
1DcD29PyML+5TRbBh0VqZ4DRx2emiUSnBDhC1AgtzCtVTjxSXpaCK22g2WnPVIPXH1CdymYsP7Eq
z8gzxuDkPJuPQNU82fdvfrkxtgL3aEydJklNo1LEAbKaigTuUnaXbq0Wr92SRBJvHXh68Dq8GhKv
mPWCo+EBpAOJ4gT9RwDJ/bPWoOpVoyrHSqzqV8VtSX27lMrYdi10Y8ae6hnkc31HsmtKsiXONBQm
dFzboZB2magZdVcbID/zm1hmwtXEjOapoQFbl/vXIgsn+26fuM+iCAjdkfc/XI7rhTb7mHHiJAp+
OHvd76IbnlRfkaaubpTln85M3sdd6su43XluJ13UivEFIV6fr27Pgfkj6PtSbIhIQ2sWTz6oz7lL
TU0uY8O9KNEykd0FrBpHxcXAhg8lFdckbUE/8yVQHGHnIslDl89SFJzh62AcO4UhDp7rmjsr3ysX
hEyp7G2UZ6uBhee/7Hqgb9Ll/oD/MhBxVGrANqBIjaXnEUw81xocW3RL4hNbBCQoc06T8nz+ynvZ
/QYzn0+OP66/nIz9aMnqc4a7kWTf+1LR1tcfu5LeyOzi6D+uSoU5MZCrWlbPeltbMgbnmt4FMBDe
T01Ozq0KqnMcsUk4K3AVaKDG3+IhLt5guITTnHA2Dr/J5jOWLNl+Cp4U63fhKxxqUrsbL4cZlJAS
+o8OBv0Ogv32rg5cdWIjPgHnbaGWUmA2OujRQ9Ib3yWt3NFXJtiB7wlAPV+iDH+1bgxj5L9J+k5+
EPT4t06yOrrxFucXPlli0HwZvl5uvn3j6keRd6tRhDC3iiR2wfIz1sYp4KkaxKNCbBtleCQgSvPv
iqJj+PtZ8s6QlOv899JsQeuHfHKUbWDvJtSTQFbSLR+9MN3Y7Z42u+JZ0TPxVpw4yOTtmr3SjIP7
RwbqF/gipbzQQNsyAiWdvC3s5hZe/HJZlkf2lTdrRfYjcFvIo36KMM88TIxU0caeTU4NNukAhgEn
ySNYXMGQzjx6GZLoK4rO/cEJ+vpK4tSKHpoaz6Qb5PFEkWUoSGN1bIdPAno0FwiTPBykPx6hgdx2
UlHVSM/p3tYAu/XomrlbO8t+vkI3uTYhuJMxec5n6Kg66sAR1Hk6B1UA9eeo3zitiGjmzZktPrm4
gFhm0ISCIW54yMDxH4Mm0mNfp00G9FHq38UZQa22eKqDjEJ8zFwLcBom5M5aWkzDMQdpPI0GR+T7
drJu89v2NW4Rf3ZaO3FhywhjhAG7SgCM9bzHBWyU4E3lCXLBdIbj6hqDgrHsjSXzro6jDbFd3UUQ
bOo3Q+ozhvtATuSDhXI17WXt/4HT6OJ9NAdKIn1JF7dZSjPq1dDP3MNLRHRWT4LRfUyb8DSI2OxW
BAnSUchEgGRiIAsAbe5h/Kt2isCawtnyPQJ7VkkL2M2juk0wF56xT03eOJ743OxEMjXWR0azulKB
XLPnBaqIKYzDc/zEUwMAAOJrOZ8r/uRA59MaaH9rQjx2q9OKloZM6rI5nVk7cxIRR1HA8oJ6thlJ
GRSjsQjhoQTrZQQe5wHDrUmrphTjZGOaOiD8+OF23gLxu1hcX9QXz+d6qegC1kbn9TXGmpdMxIsM
rUVd+eqvSHitNPR1cFPkNr2iD3b2cU+fSPK42Vu+c+suLJslGKYArQA6v0h/o3dckUv2W5jYF/E7
87E4PL3eRlGeiz+1/5wW1HPPpwlu3bZQRumIRq/FqeAHExLr0SxVwKHbO1Hih7OgC3ZlBvxsDrA4
MCvSl9lzPpdLDSWd/AFNBJONHOeBclF/2IC3yAvXGaxwsRqNavm8jSG8o/ySPuv4lfc4doiSnAyg
FT0yECVs3HowxMLKjQK9XvQkMLUs0/lDFNXEED/jit/NIlLAZrym4FCv1Qhv3QNJwbRg9NltAcjZ
nObq7sCjCVfcGd87m/bfy2jb9ph2IasIw4LTJyEYPWeRq1mnW8z9pcDcjtQ8OqTSR3GO8SS8rTXr
e11jEtc7PCqhqEsvBi9OgMVfcpTo3NLfM+nE8VnKbZcBZw95hqf2ULZGIDNsJnPtcqnFGYDZY6fw
xlNTZqTn7ICByGKs5inaQWY6DuHrs1lxjSCjskmtxI3/s/7JgH+1RsK2rkx5lYqCPAjs9BMyXnL2
7Hx2zsPNscdFZCGAr+/r9+/6uvdO6oyroeIErUZLvpa/hhZttJ+TUymgZ6V4mvdopR9ax9N2ePyT
QyleVrHFS1x0KJtnVKNT8CtZ7Q6+qZtzvItotfcSVHGXmv1XEm8TysVXLbFhds4WTC5x+EcJff+z
qDjb8Vakhv5qDn3Dq4pj0nLsJ9Yt05+RTpxW1vpFP2XpMMmnT0P4LGY7o3ra/pEDdXsJ8A3t72Jv
68XORPj3HFsgZ2/GzjrOwiw2kKfIDZ/Jjd7IpNZ7mXlyhmDPAwFekY5aQP2tjaIDxziSpEmsdKG0
HnVfIKMqgm0KRb/CtlhdFPb/lST5ffd6P4YhlXZwN98kzGcYbeIVc3fvX+ffhFitzCin7cW/Sh3N
lfhIqMI8Xux8nK6f3SZVFDpeiPKZZgQ4UAQCeO0ASyVgy4Np4CKtgMD7wJXIw1nWhPJ7WWwy62GL
LywLORN61ohYM8Gx4DOKhXgCvavsGFskStrIPA73ILEkXJTnKtUEFuaGakgcBvQHn5NmoDcKm7fe
4loTyncRaNVHWAZ+S3VjX+A7fsGIEU+mDcKG3XW6S5J0N1HoeaAJpESVIzx3PIWcPri737N1N8sk
1tjlPnRh8yH+EARE/kbxnzLVQKdK2hqTpnG0/A/nPdmRsMJGHc7iuj3X5eCZm1kVueUtzAR9excE
KJNLlPm8zT/SlJhX7JOed09E2fNqWTLtAEX6eA6Z9FeosnVVHKfGEfL2jLpgFq89/cyMJkCb63PE
C6ez7klG8XUhHBO4yUIAe0FW4t0cmGeyy6SdMeog6HK9GEMOgR3Hg2bXxTOZ06UXHdhzr2nyCTRt
fYpArj6HZjjEnUBXGfnrotL/ikEZIsZ6hK8yaEe5D31Sn+Z2pY1blR4kzQQiGtOtCgX7x1O2KEZl
6A4Jp/Dm7XkDKmBz9ROfq/BoDSqYEdbPdYSuBv46xvZZ2gUx62r/C5S40sqV47laalaipFDN9dSu
pi/hz6Pv92OAjqpc8nf+LElrdLMkZlsYGLZjBPj6s452w4pSCPsXIHmsgwxtF7WdXfqLes3ue96s
x3rtkRqZlcRQqh+A+O8NBOVFB4+3/wW2r9ACLr4WzoKQ/lii5Bt4hNLQOUMqfeGfLY9tY6zTjlmd
8gswc/XtgSblpHfj+54XxzJpxgvPoj2qxZ3O/YpxKMlpnsiy+IpTZlHjPi5ZWJ1jUK2/yEtvralo
vioXkIIcnHXKDqOsdKvWQ83Q6Ji4/FObmHaep43SK+7GLixMgHD/wncM/tvR2eBHlgsN0Zaft/6p
KQkaVabyi6Zg4yn2YHPS2oGcOeYtnNTdJpdT0XDKzmlRkXrXaKM0trk55sOq3WTQWynWkMc1Vz8T
4ERWlol94VizdVqowx29YiwNoOAltxbWbWDeEMcd0yJjIuxZ4vmjqm2D/Mi90bbNBy/E1qM12onz
74+8zHUJyO1WoiluXo4Cve+kNTONAUiijtpqjv/ViuFTxpULrcL3uLgbJKNve70zkHwNTI+GeBE5
jqviejDrBFMkmhkEUmY5/I1w43FKOc8/g50deLCLuytmqF6etxvSsl6zH+t6CqDt0p9GRaLfVT4V
L5xnfdmbmrzggtOdRvwBzV0w+8yLDLD7ixaTsIkAKlmwgYDup1S5K9PWS+Pqh5z3FQLerY3wmSVT
ORlFA9FlYYJ4hQ1EhISfSAMf6RRkY1y6djxPqjpOQX1glwlfSoWRme4CgvsRrhNvmoZG0UqK4di9
LP3n0YbTvvN9k1ScYlnARCi7qzNZ+9dqrAK3vclyi4xwuBMW8NrB1QVoGd7CJZfVD/GkFGImMFil
TnA82vMfHeh/2B9SP2gy2BB8x/pCRDsg5gDa2zG4Taxp6Go49Gq/2VSyUnZmZsiVLwYJx2Ad+fp7
459X7cii0M513hdQIKwegFjpGCtHR/3AekYIn7iJJivxoSIcTuIMCPMYTkGWdDgmjx3tEU8T5n1L
dl0VfzAzjZrhYiDfXyy8xnmTzRUZyLDSCoEaBg8El1/zhI3axNltitmjk2O/AgxrhVhvPhrc40A0
35UuzWDXjZfE+HwIaqS1PzsKgsc0ybWp3h1cb3uqRmQhbdwWKQNY4FakK9wijrUJ4/aXI1Z2eELq
6+aiEhyEtp93IVGbGPzOeR26lTKBVcnjktIICor0lE9D+W4aa3rSs9DQSI9G/uH+sVjm0xdL++sX
RSuDnxDzx7CxPRpa2cLTqWJkqmP7+lNfyM+GtdoieGWGJfrjcfsMcJ+/xuVczfRyIUMP7iiepl6g
x2txCX2ArngEMLBGLDNMSzrKYXapRdcCpDfbMNH58I5x3b0l2Lq5ANT+OSTOAn4bRzHyevUxkmfj
fpU4NoULJR56ZDPtXDLXZ8YU1soL4yMOmVnYaMSkjMiFx+ckPSSpmRwLJbIw5TlZaTcZ4mYDa61q
Slw0ooe4DcqWXJG12q5JB2Rd+ciTchpbR58VnMcU49jkOT4Ll857PApGeXPHLpoGie57mrZGtldv
pR2J/F9mTYG0jHU1y/qJl+blEoKMFoQ2dU9wZOGUSPKLDMBdd+S45VnR1iiDJTZei0TcC0yGdreH
fKM6/FDo0qK24jQN85cdMheW7HkHE1n5VxU83lDqpvpZDifFLtGbKTEzKOTvU02IdjWrfCWsN51a
kAqFjz68PWc6xCG7pLaW77BDX1STM6W7nzlKbVpRGpX5NYRvBvGg8OvIgI+CYixykHgphLSJ80ca
6QfS3AxWGm/nbJ9zAAQ48sGrFJtBWVLKdOeaghnXGbcEqUfwXyh3CvZtHuEXlxjdhxkm71LerIeL
SqjxEhiq855jZTJmdqSmRkZGCJnov3GjeXjF3Tg4Dr28XMWTg7romLncagJdHedVCszWN9TE8x+M
84HSwr9RPqJhxCcfuHmJz+TVVrBVFgZ+UCn3SPxSVsCisub+D6ukux5awCkJIekl+ZbzCMH5xj13
4eBH+VhJ4TuU14YqBWfMcw1dcsHrtmPKyzTABSJjDf7i+n5+0WgLmGRv71Jsf1keSa520KdjEJuk
a7Pd7RUnixj8Lu2pck6LtwidnXGUMBhOO6aZj5b4UzhLfFzqkE3RRrmtXBJjOKwdbgPdD+0YC36Z
YEZqaaVWmdKfXvWhe6B8QewnMOMti1R7KlXXnxEPNMor//sDIsXyzx/rVPinLWBSdGhmKw3rluEy
bVOGOyD6yCg2ZfaMMGLraz6lXDoGz3GxN/qA4yUH+YWHdgY913KsM+iz/jtSQWUdFPKUPpsTDGKS
YIsdjAaDmT+NxMYER5k/ViX1Awvz77HHw1ozeMTjLNjhbmGe/InyeTac0bBorQBI3hmtv8vLQnrm
9XRVhg3JvGCozdARqxe66jQj2pQpKDTyLiS1AR52G3+uart/R6LGQRFxwCQVbluN4z3MUj+nWkHN
d97AcRWOYU1L1PVBQJsKPYNwtT3IoZ/QSHyL11ISDsBcV9zEZKuNVBVImLAlWDMrWxZbc09n8Gt8
LdspAH5ye7VvlTeU39sj/e5FGvmLp6lDPv4ff5UMSPTFo4a9VYS7K6YVzK+BQNg54l0E6v1gtQVo
GZS8XRc0XWUhMJM+HlmUj+d+6ORAQZZpjCWgLRYJD6vZWFhOAJ2TGMm+JHmqH4WmahW8oE4e472k
0kiF58Ek6Mu4haRAkwqzlmujdpILy0/jRQnXVrxLbTGg5ayDGwiLXN23KgbJRlmZwefOD49QPQbO
kHP1fha+5qZWzaswG4+V/ILJpyMAFiNZP6L7eV5PL0NCKZmIhJgDD5o2TxAOl6naexDjgcoS839S
9BmaBs/bpMI+USJOjHt83Eh3HhgRvQYW3pxPOj2U162/zRtSXeS6H/fQTRlnyP4G/KygpTBe29cx
KKa2T5iPjgleRWDdyttp8yxEnq2PEwjF4vDlnek+oE8+ohIKFIR/5DSypt9YEDzjgLRlg0o1cTWL
gkw/18Ya0yz9ffrQGsOd4u/Y1HltPzAOv7wjBcAhtuU2fS0pMH/E/JKIY1VHccc5GzBjYMAPTQxK
ZhyXvrspSXhppO/LDkLPD6B0i9Z7nQebqUXPWoN73rkSNaksh/duYeOIQzbPi5Hnr5fLgWg6OSJj
AyMG1bN0jJYia3YuoF/Nbg64pio1yZh4REdVMqeXALrmXgjerVod/xkg8O+siZR4v+Q4e9Wvdkxi
bZ0+GSrBOGnP1HCk10kZFATLSHB7Skso93ZpHG+TSppYlfyd1btMcy7PSgpXE7IBNZsC1RqnKO1p
nux/W0kRPybKkS1SouRXuwkFPvQaBligbryLEGLek35B4Gs7OgKsUQl6YaYGa6h95QevgQGTsSS9
uHmJQIS6nNgamoNYz3AdP5cOpbihYQ8OA3swQD+MC3vxrxvm8iTJ+qTaY86dnL0w5+amVun8mkai
0h0CukjVrXCyausf7N7juECi+mCt4nzGGJY1F40jyJGGjKdKSiJ3xUkqG8gdboQpWofp16aqz/uH
UvOIzVdpL+Yp1kKw219e0LAO+Vkc2UoiZF7z2norhp9rBbZecXPwjEc/WTu/poNi2TW855d2QUJN
kVfzAmGoqhD62jHfZ9R+S1zBsAfhvsb6w9KwKNFjUF9U/8noyF783HxVRaEjns4ijQVNZagjrQlk
pMXCasntl13damII6lKuGCWIa+joSp3Zf/YinCrBGfvBt4omPJrJQUabkgbUTU4CeN0TIOaLdfJv
xR66f5A6wKGIyOwFSLt8EgBDYpgdWSt+adfUY19lBCQiVVVgdlJ3Wj7hkHJ9OdZOZsioPSK3wB1i
2cny44fFoxbx6ouveSEtxZyhC1WaAfSgW7TvaMMNIz4UZ1nA9xclBezY+aaUgZ7wsDo+W25ILvle
JGtVTbWggNhlgPGHS/O3KLPky+X33dD3J+p6XHCXD0QIg41/xtvC7zbRLu/YY6rVNFFHyOTqmGPR
7bFFMO7ojagoBhlCsZVmB+sXJbeVnNOzeP9umuxMLubiboSiPHzfT/RugTg85SzCTLmC8QtATb6V
AZ1EpjujPbH4FU1mkeoL8RSHjVWlCqtDUy0senve8RMLNAO268qya39qn8oEMXOrmBOkHitL+QKl
dZ9Z4bcVxUR2yhIVxYvr4rQUmwikm7nS2hF5x7uaHju0e7bu5E53EKBu6h45RfULHwrVAuQcEPTS
wff9VieErvJ8NmzDX5RwO0/BrE0jP2Fyp3bd/oN4c1PIieZQzu2DzsOyWBJisex4gGMplVw7KC7j
Bv44RtEbzjXVEy7XRZ3sPLuG+MxqEpBsgKL35NQAUMlUEpE8dG0msFemUvsgAMqM06MleAbvyf3O
JHe6hp2Oyp3myX39TdGA04ZiAMMG781lGW7k9pih++GIQ02uxrr3l5VjcozXUKSWgjbtXzlMi+3w
jJajDFppLmYoh8Tnph8WmoqXXAaqQLc92LSuo85H+v3j1bi2BsEmjmpmz+A0hTLxlFSDvFyo+K79
wEz7MwkqRvVXEZT5yn3b9/MJXOY1CfNbzE5toiVb3Va/ILrW6XUXtCC3Q8x4Y4QUxV/vp63w7NK1
6UZqZD4FjGOMq1BGaeb3QUKe2SGYkhXbHkUSc1DjQelht/L6bsDuTqQvc4mgmTroxigtD8UqBO5W
Pk02NEHV0mB0RHGgCk+/Pr3HePd5LGORcPkwIKPjY1P+qbNeSGBT7vgkne+JJ8BktXS8ssN2HGWg
/rn8X5g/URs6+VHvlXMo9ys662T/anaDIjkUSUQscLJxzTLg82XgufmDaFUNXhjZR7LX+Us9PaMW
3MKierGqr0HkZhjbYUsvIQMMHu7l1hxzSCznqjmjfeaCeFsHv/72L9/E0s4ZsedPgCB2ls2JYknF
GQqRIKOvHxPiWcdHURS4CfI78Vzja4v4gO7zvHHrE0lErH9wv6dnfgztCHUyG8NpgkRpCbtg8E0S
yGbFc3vsziBqXfZRopyQAyVxbYWmmq3xwh2O8M5sEyU8o+I6S15aJUxEdY5UM6zs/npfZhMOl6tK
EtKdbJTP90WVOjUCH7ldiCEUURelF7rVWV3uA3mPu0om8Bler9izODmOZEmMmsos/eOqbwHcF/Di
IV4s1WElVfoiHTFfTqz6ssrvWQHaBpD0LrvlnL0iIjM7H7Embx+9eKo+PPKsNjSDYNoPFOh3BjAw
axxFE5boU1t1jSKkROB17xbNRUEwjdHJp5wB3bgAykAh5Muz0h8JYhslEXlJkhDz+KaEtrzuhV3z
luSnRl/IGHq29HyXeT0Dq3BGNWDVGW7Rd5qES6+E2wrYehmGHSbe7f2CWhPECrRHUD5GDmB2lzXw
hzOH/oXcSmMwdhK/1jnJq6upiv0C8hp+/oL5yHQGtd4uzoXYcQn1KNXwihzL4qjfed6w/CaCgWdy
LbOcApIxvLEt+0s8vdjvdb1X2lEWYluQRQ5YltmtOld9MOEiL3+qFOgS1JjxfYgCz1B+IqAIox/A
T/n3CZqG4liVdJE22AhWGwbo9hZfddXrLTBg09R7rwcl9W0pEbCZ+d8Bn+tc/S8Nyf7GLR1jBEvX
MVRXwByhDRKXyum/Wtz+9QoOIeKGogyQumdSKLpsA2+Rud5gYIlwa1LCSSR5+vDnpYOh65xlbkvy
EhHWpLoPXwOAZd2A4lMS9vIC0suqZQ2dpHrRN9uhdgMIIfmbmtAECDdOdN252o7zNZEFvYwV6n7I
eRewTXnYjlv7BzECk+ZxT6OCMKzrB0ZAdPEkYkYZ1+pDNhpcZMdj5uSnkrpwk33SQ/kgGIJiJZMa
3gJLZ1mHcSPXfpFTTwtY79olJJ2VFPcWtOjkeu4A5sTqqJhLQDMVaMsUoswoEpKEMZt/At02zN/B
cne0GimP8EFGSfkXVf0JSbfbYeRZxms+oFjRKly00uSHXmz1kLRELDMz+l0h2liALSN/LC/xifcF
zfznrz8lKCLR/99m9WtVRqLFnGzdTKedTd7BMp1NEOB+3802QT61Tt+AwOMIBfxCIpATAlHvT3am
JHfqBDOsk/mQUxsj1ZrhsqPS8HEOSd0+B+CngDjnM7AJ4zHa4cpiZsjesqbnjjyrXcuOPe+3MGDu
XcyJ5xhdPCLsawNFmuStF5Xsz8qqJtWe/RhY+zvpkSamdNGcZvkhLBOiQCY/sxn58oHNl0pxg6/q
AIsJJUUv+dt7nBqUjR60FCe31/AMHMVgwAcnzAiG+DVqh0arC5+OZD68Vz3PhBvgodAi1jZj45nE
XjSJGV1saQDvfV5SRE1vTr3OkIYA3ppuElBxBQHnEZ/3AL7Vg8zVJBiqaRj1/zDqjKSyM1iXEpAT
TBtunHUfSTMpVq53KNuAbgDp6bXQNpqlc8UxD7pxU7IEDihI/OEukDOiqUWTfj1PAjb21BxjkBao
7newT7cYFUa1KOIgEnJ1e05z1TcY5kQzH6EoObQ9i4H8nhGwkCqUzDz4Drt4L56iAXiVjrA2SNF7
wGiK+XHrY8Jtb5Qcp85k+n+uorjeHBu3iO6R0et+kttFi6F7yzzCeIPlKwomKCHsIhyA/DUHV7DY
ymfvIrl3GYmom+G60foJfezRmGNs95PxsXRrMty9N/qnfV10hJ/LyqnVBnsx/dL6fUiwCXclhzs1
JhFlSEsn0KPT26X7woMhPb7DZ5sIeiC4YZ5CHwpw8/vOmzxlveNPSfWW4vAWTdPmf4plJmbrxOsg
Lks2rx9HVU57Hk+81PPm00vb0W5VdRaI3xiTdZLIDAMzplaF3C+QUFY2BCLyhzfd94ccY0UOjhw/
7C7Ek1jZKc1jPVRnZF0lxlxXyACgFcRWm3cQBIzp3HPcvV1I/QWrofeWC14Ic1lpX5QyytlS0okw
Lg3IP+8cFetkFqfZXDeZ956qFhGt6FYig+Kpf/HpC+u5v0jAfofyeBx+nNCEXVU3cqORMvJ632oE
9N3Wi+RokWmXEU1Q3f6qHMFwC+h8bkyZKuZRuA3hQGLFGAclCfhP1TowHWqB+DSmDKvqM0NWnHEq
FqkIAOZ2LERfLZTIwyKdcVMFFQUM5mS5G52j5bf9rcjerWn3/Py+DyAmqRGr10QTt1N3SVDfdf2p
spN84JycPwyk08LwgNCeK/xRlWUMbVXHOkhrPGY5lu1rheQZ3A0/HtNQThQL7U9pgr+vs8fi2/NS
GbGixTbnhLl1r4FOy1PvkWGexzXySJCkshpS5w7YsOCPduQgxil7ucnQ/1DTIBwmkKQ2/EPTTFBy
lj3byKVZFVPtFrVSuca7RcXcwm05xLg1KfhM3pyykDvg5R96dpK10Fhko6Vj5TqHFEUK4suE1PGP
6tiUs1hcIKO2HxQk7WCBz5E4ebp64AMmJBTwnnFSJBn/pyUQCKKoTPu7ZSqUC3hfHNb3MVEs2gUt
kBzZbA91Fi7BWPsuLjfxZx3Zpn39F3RBmd3EARksKFHJYhpgp+7tM2l0cc0/fC8EOrqPAiNtsmpj
Fo/iTMMA1XwCqlAi1U/J+aBvuhsKkFalum+jomK6hl0yJ+zhPc5gLqIepLKxdyaaOgnuW0v4aS2L
NCQoVKWdy6m/qcKFnAbN23t1xFaGc2UiEvPozNw6VUZMZVCzdd/6FcXrEcryvNTqNX/Z0QK56cGE
JxwujJX781xALwNO0etq50t1+kTieDbuZD2YhJBA+SA55wMy4YsApJLhcdzROSXeHYB2SJFYFfXh
Q+aHFt7Uw1Cy9u4b0nGi0GI69rr907MT61ehN7B2bnwZb03wKrzYtzA6OrWE14EVeISSeaTz+LAj
g/Omdri8ZZcIyOkPBh8CXGFeclnrL9jD5fTcq8ttyIqLLDPbFw7Prgtw1gU1ZB0d2ix694cfbzdV
gC4pOYtDNb1Sk0o+2uR2I2weBwqeGMD8wfEFZxs4af88EwiPTIIborx78YQxd5BJQf9DDT0sCoiZ
Jutw/BKwimgpxJkQ52IIVywSog6wOUdy0K7gKFYJxYin8sT2Tyi8qtl4jIdcJRxW+G+UVb63Sr+O
L67N0ooJnFIixlVRB26hVGL9oD89i9AR3JKjGxM0TYDuMUEEIZAodZWqmkRxP3XnCfm8F1mRkOxA
f0ncSkOkztQpnMhYca7B8hpwdcIvMXn9yqcu4ZuDEjSFwnPMXtQ0nXteEVd12xYrPGfgb8WpBc+V
71jxYTO7fIC4aHwcYG+4S+I1tpw3bB7X5esy+8EQnBI+kXbvbQF40c7e7UzAfwPLC7CMsYCW4jt8
fVgwYreVBxJuz25onPqLMw3K43Tg1pOW6rLnsv/b8IDQ9+C7nhhMibOsyvK7tTY0V1sTcGq1xcXe
UbmthUeXAUrjXSJVT5iPyH/ySs+2yyB77w4pwsSu8WOl8X2HehQeqzEBCnveZjcHo7yNKJl4M+dx
niUMTS95YlbrY1D5p/2IZFC0SnS0X4L8VXgSXFjVtNRliSC6tMqAYz+nfuplCcqrC9JGk4GHIBmH
rH9DwwYicZLt6sALcmLvg3I2nDfgYGL4MFxOHXDMhRoxAJtYwDGIoAD76BwMlPN8CKo/Y9hzEDOA
s9Q/O+8K1tpIVcPJGWQI9dO5kJ0CIFi/ooNbra+QOlUboCjK/b6yAy2W26wiBX8LJnm1zk/fLI5F
v4vDdnwBFDW1KAT/9QcknohaMkLOQTqyL4aADMyXIEldJoufQsPwyclAXAvgfj07KrUdlH5oUu08
Rl8lL/rn2YNNWO+q9XVCb1mKGD/in/5H1rGu2NBStlvUiGYGw256hnVfcCQbQaroHCm62Af2PHqp
l/WjDHHRJkC6HONcuW0mFMwafG/FQ1RgNmHK4C/DUaFgce+PcXqHW7XO0VQM5gK7a3szzCBrmSBw
pOYsjtzEcP9FYnHzU1i3Tt6o3GqesBdJvp4DEJnanyY5VRMvI679bBBJK/zic6dw372f/sIEA7wE
ZKYzhdODQBPPg6YYM5waABMFCaJ3ZjVhmrSZh3wg+HVHuxzNxr2nIJWFe496iMWwRYDagwBeL7OD
g4BIfbFV5wf23MySYIvj6RyVZjKfuiLZGVwLSioZUsGLgSFPIgHwF+ddhXKzHs+EJp5oy9etxIZh
ZcUuN3WkY3Oa/PXzWtFAeCD38KRKFbMNlkfNxisGKwpglV9CNDkcAxicyXniK29cymksDBApH/Xd
3TYrQKRs3+gcYKIx6Skpqua2G5i6ve2SNLSYk6MMBdz1x9W1uSHJPsHw51gFLnlKjMWFQCrgwCDg
ThRvl6zqPGf13EVnpxLrZYyvGRVdmWwdbSZ71/JubDq6RbopTEodrdlsZCY6bqkJTQ6mF9V8Ljxn
tvxVAHrQADC7YlW6Gfuf647l+Hphm2v/fkKzTe7MMP/sLlYmi0vmC10l9rL66vS6uAW/61yfyyl4
u1bjaDHUsLUWFu5ctufzOYZvAHiqGABtW0lMiGpzknCtJsBhtk0+PGbk1JRjupM0DDYvHXevj4Km
ZB9Hd1Nj2+aG4Pic58JAL4DtRDOd0i7DC0Abnpxgf37XxKT1nvKGXir86TTZaMG1vlRDIVpAs1OB
GSE5cMcFpxemG2WYxKCIySEFDRU3itDpxmBTgl+zSe+g+vwUzV+hVOeQ1zee6Ofoqe0P0UBofYQg
6cGcT/HviW/pnB4Ix+TpPmn4rFDBjJwEjR30qjEDbPz91R92rrert4cYKg5LAzxtOTBUVStaNMUU
k1n569jeezeQV8CGaHA79PqkEGR4N/c3uwLq1erCb9hvcUrWvBh41Zzhv2WJwaDBhQX3kR/BWsLx
4pg9YdhLBkxpDzBnuIojcgAkjY5x4DPnqyKJLVxQz+i0GFYdGl9qytXOmIbTdRGfW75uTTXvmHaZ
d/TNm/+tnmNctRCeeANB6izpgePFZ0C50r1kaepLyqO3SC3cvHNEPJCrW/RqKon5KaIXbFjLmebW
hGVdxPls0OaVXT8usXdo9RhbRvJFFLeH5Ao5UEHwbVJmixrVRuoBBv6ymA5qiDrNIOMIiwA0eLdy
Qo+ElEGpsQ4OWMCfdWOHxL2cCM04grxfTuVG3eFHgvDcBExjh22IqO7AWIXf+Ib+kopRRpHqw3lj
Gk8VUe66ikDa53bT9LnX9qXVK3FBqs/5xjcSrc4HvaStxNrR0PzOiUC1DnTO0e3lM53mKlKKobxJ
/PxgDifHARXOBpAxlj3mHSnfurWRk8IxderhkF01DBJ0tyEW9RB9bryZqneJCag8C7cmz0d4ixHT
4SFdGTj8EfGTthFUBC8ymZ/gJlC3Elto1ZyuYfdk1DMgsqEIfwVKvuslukv/mOdQ7pMcIPFfiYKc
BI/F/u6QaFUwYz0xLuK+MRppExh6SSqyo4z6k6R2g5mlUZCxQKPSGvHil6jU3bCaygR9RQ/9SAIr
BXdbu7aihZqwicXOWRckoMN9d+nG1E8cGatD664C7KOSdCx2/WHN1Ege2x7dpEH6Kr3OuioMy0cW
1cSh0ytX1A59VPylc80/CXX8eds81fr4KumDRoL4MX7/JQI8CMSJ2hlnliacw2bPxG41zkcS6emQ
0h0MCakjrLoNKCAp/cPfdsMbIJn+r7DjjQxnTfvsi2GGH64GCjikAuLKNyhWxtZ5Br5UaIMZqpgB
A65qIC7qJGwIw/ZxBFETJwqkGIC+X2IMUji0GW5tKg7jAmdfo7rJhcfPdlT+gUzX2ICQsH+B1mba
FOUo4ypYZjTTKPDHbndVqXp0om5ndmr83E7v6OW8F38tuS54FUFfstnivRndbiLDKVLduk272TIq
u+kY8hun8bgBoeIcXsbQT7NndII4fyCSZpMaV9WADcuFyJ/8i9+AC9sJ7ZVIvH/b4B83ilvSSJJN
uUrNXcxs/o3uRt8hIV98jlQJ/L8t9PK9xVcDVZFIOPobddlsbev3rPGOWH154Es4KTD9Os7AX6Bf
kOowA2KwN1b+sN10EMS1ht6Gf2v9+Zo2KDQ1fka3VtYYb+WA9qz9GqipH5s9scPJ/25NW9lGYPRj
vu+TBB6C+Fz8quBymxXud14dv8rBX4EDMsKZC08lyGHCbtce0YNe6jXRcgPW5hZ1XlvVAavu6K0O
1ePRG+A/6IO5hFb+WieC7QaFbngAAiv+K5l24kpsjs/l1pLqpZsWAzopfXnDtNlZUsRfedoQUDYt
pwzW5PHEn1PDH7RTz7K8AfRzOLXu49AJ50uj5PwBkpQunZq68iAV3x/RTziPiD5N5st1shBTMK+n
dSEc7tMU0WvXPTlfOvjfJDgCoNOkFp3EHj+mthIcCFh6BwdA+9nPX7OWLZzs1Wnj9U2rXGb4CSym
VceUAy2XPaV/lWktQcmvIDsc3zZRqO8hRJ0Hw6WxsSKBhX5L6XXdV2xvVpbzM7B5I8jWRcO4lN1Q
qg842/M2kIImYP0ex+AxHpCPXAR+HjwYemb4FB1T2SIHlreADwQdxK1LH71MFIb5a1Q7RDT3nUyn
cTHWKYlBbnopXhbu6wB6R5D66We4xRSM0oiUVJVRwljDmx5W/DyTBkVUmNEOTY7jGBRz6h+8QQ1w
i4FeoqtNjOC8aHzG2Wr3SfCdKw7M09orcLHCzHXcDN7Qy1Fir+97GizGij1+WpEH1B2MSFd+2/Zx
DyLD/dmnbRPLNtYIrLzdIsh5YNm8em2wp53B7RloNSWUlOk5g1Yp95pVy/7c7A4NMshw+G0S49I+
DsXQEyyGU7s29whD6s8wI/2e2+aMeX4cnxmAXZWgTPNHbqfS3T2uDXvUt1kokwHOKunqDPxWTyA9
pUkIJ/EGw6oHW32LYq/Dd67Ixz6muN4Xvi/XlrfsPLjLubZmZANJxWdLaosZz0KcfIuYQDjkeR+n
xcYWXj6G/KFCB4/b741a/0gH2RsmpjenATg94/Bh+v8PZRtAruO9gxjiP7b6JlhyVuwKhUFUATIi
29q0x/P0JGK3xP17reaa/48M4iZH4K+1JEyAJ07TgyY2AeWlUyyGAPAVgb1iPEjlbw6Db89yOpcS
40jcWUAA/eQzY1pFj47Hq3OwbLmvF9ZKaBLsiD9Lq+27yI75TR27pCVP2vqgv15TgkGavlPefnQP
of8QvYw+CIaoDkfQUIKeLacIQJwm/DTDIJIZJav94h7K65hl2HdrLY9h2PpltjCBdPYB/JEJgSWq
JIeAdkl2+lYCGmZdZ2W/PigJTD6amUq8ZdGJvS/3OCuGfawnKOkTxI6uXJGQoItCEN4YCmWIPu4q
vt+VeKkxszKB5/E19NXB9jd8vOVEKLRP0B1KkCAFSmbhapRj6xyeV9kpPmsESe8PRTICnjiqmjal
7Wc/RPxUtZsbFINX0zfzNLpUPD0uUTt3amWKJCESWyvO7Jpj0OuKqVU0WhaAgSm/16sQT+Fh05Uj
MSR4togMhv0H0k1sH/H8r4VpUDyayTLOwbGc7M401vxRqit7Zbttl8G1vq9hxNc7BJDhQUWtZ18k
p6O0eAxaF5Mq+g/yATuhcu+1zlN1gNbVXUozwBgqXLKwiv8MwQ7iy9FsWupWX74owbksvkvP8I+H
oAoOTw82irTwO+7cl8wzCitbX5/gz4NNqpBCZD0wF4+8fH8p2tMM0h5JILKRNx5Aj1QsMWKBJvBS
Z6YJFX9Uv3WU6yRvmEBgCFgLfJLO+5SgjEcx1lN2HhM8q4OFlZq/yQn899nGdk4KnRjAtCQ/utS8
29C2A0jEaw4qr/aw6CiQHjZEuGY34BrJrBQ6LH4xCF2TESJXDFWINN67BhlReUghrkMXmr0LMPcn
22D6FKYowQHZrGFHZzKGPNns9J3SrBIvlc0KrZMDVMh2M/FyB8vgL1CY/eXbWBO7wUnpCoUegfS4
lktzyFueS8dchou0kl8yVH3nR6W8vTqmlN+JQa8gIO4ot8ohEzGbFTjPmrOl/ah4SAO8t+34NK51
xPs4weLZ7ubeA7eAfWHENY4i6K/q84V6DzJvBJJyIMYgkQ2W9QywC9kjpgt1/Z0f7S5+z9iD88kk
fw7uMPsSkKJbjcYcbhzE4GfwADiHN+PrGb5h5H4Ld7trXQiHetVRYUGpQAv7CqvPWhslIgQCw1Kt
wyv8ywqpoixA2+7+jfYo3rs2sT/2P7i7O/AqqlaPke6RzTja6Ug6Jsy50JYoReI691r//HsYWXGd
B7w6cgxymOLMQ6SoVdv3MCndchGq9EOHC37v9YznES0ZShCYFdAnWWGCljTRedMt5TAaWWrw7zjX
SRI+q2Abv1FoIz4rhr3GSiJIUjPoO4JEcAljhOxI6Lxn8xQE8emo0zEyWYhxifSE+9Va0td8NDZ/
gVsaFyP+nBTklLnSLFl4bkhFYv6fKnBMJp0+MQATtSidY1T8vJM0YNsDdnhYO6Vzbf2ZRfJqfxMs
6uK5arxXAS15kk1aDICikedM8eskjuMxbFtIEc1N1ia41O47wPoI2D0ootNjG41NpIoYwSjhS+X+
DENT58xPG3+SN097z2+5fuEINcuVIofw/O1VvHwLYxu8XJ/c7F+sxmDeu9yGy9jqMO4CVzUv2SFm
GuxAmaCAGcS633qXXV7HYlASAVh0pI6CH7MmEi53rQ/0l8WHsdNOEPsgUbi/eCp7pytGD7csK84A
/UWPXO11erd1FVjGN1sm1tG2Df3Sv+r5W/brkNKINgllnU/81vyStPIo3TIJUoGeQD6tD+EwOG3y
E6Z3ig8QdfavlipB5dZXuLbe6Y8wJ38VKnMvXdJ0JZJw/ZRQxlnqk0E2t4ziufvv+Dpdd4Bg1Fw6
38p/J8Thynta1FovlvTjVdAa2jo2HOf367ZviLzk+iM9egAfn/YziuZzh9rq0chEaRkreB/vpwmW
DB6S3qits5O9YpVErFEdq5Rofps1qdI7dSWhqHt8/2KHkyBKylkJywN+VqasVhYvGYLAen62dnZO
Kh7hcW1sQ3gah0r0qinKdeHO+6W74rusqVnOxTajQGKZ71GdHQBm3hH6evDqOCgWi+bbvh0ZhZ9l
BOD8cZVZhg1qTZMSRl4E1N0MnMJy7eMGcce2yJR6ZMgThqGXk8Xqu8ehMesvqGgpkVZ/O4+63j+A
b+IsNJX4cafwOUagEkv3vOyQTUX8qt1Vnih6inURbRR09OQbPI34deS6nVyvJA4V/3hnVm97i5Gp
khdjhvlxWyzz8vZd0GPynXIDoJ7gAaXoF2Q2rT0kRCNHFFYcJHPVVlbEjruBn7JOs/RlESuzIg2l
aPJifLOKUptM63G9xvVgb+alf+YnpmO6iFc+qdiXsTYjp25Gx/DIYKDatF4fmTYgUnawO3PEP1E5
NBF2YhCtVTSemHNli/leTEIvfvz+hoBfPbN5iVhro8cLeO9ogVFYlNqGXzrf7ul3BZbb8nR9Fw2W
72mhvdKjiXH3eGa3z6J1kTnSyGOEPXhf62DQbMMnOM88RmFm3I+JJVfdN2QjYvZVaVwQfMy+eBBM
6VZUlYGAok4b9pOIdFkvBQMT1trmWrOPobkvQEDBrlYy8wt71xLoUAHntMQrvLfjxT+Lj4Hz94h4
549h8lhpHZfe2V18R/kYmQmvvAe4xj28aShTtM7gKHR4oJoQkUmSQcLGfdhBoJEOfGySIKW6zMe4
Q/zqSbqOjJ9jkHvSJgPBBeccvjj0IstQaHuchITZlOYW+USdgQYSVUgNGLQJmRgXKYggDK/1XgWP
3I9QJsUCKIl8bGWp4t9sSmV12eBMIuWxG73NnLh40QVxrRh7d/mw/D7ookxJZZEZnFfpomVWDLpf
QHGVbOgh9Gg6z0fiRJUOKbrL+FvwFi8/yuOnPKVc8VOFjQqb3zLngR3AHpITXpDgT8W+GwuTvAZd
dBqpcuZallOo5Ld6JfbexUHoBivkvbvgTdqeNtYEzXQfFb4w4KYfuzd4GvRQ7OtyvvPz889pHznl
IlUe+GOVLA7UGVlW6lfgbhpAGeZMmYHPob+MCodgD1n9ZWlxEuqriyHVsRe8dfna1CgfINLyjUUp
6+WZzCvRe/znS7lpCtBm9YuiDgfdDp8UKU/JAhWKdqfK+WXYoa+qs7lXXSp9ZpDb/SDtrhCLgIab
srwkUA5i6ah6I7DQ+nQHbBbEs36qiVk0TQmksVn19+Ya8nriPjo15BRlRSHRlJdkH6Ppx8y/BaJV
sj8FlZiZtyZk4TDqZUVx48s/IXspkQz8tkNhgDwfnALtcgB8VAPyIt8ZKEk57TUaHoW/B9/p0hN1
fWV4kyRHtb8g+ezEVHsc5bWUEV/gfCy2HTT+jK30aElk2YLa7Db2/HQTbTptLySYNzbvnO5XKDhg
Map5ONkr7vxof9XG8SEl38+rAHcfIpESNY6m2hSjv5VMeypnid3gFlgbenXYGTs12O9eyq7vUfJ+
E6aEqpOv8Ss4XnSZlP4v2VJ1rmlfRpqITdgMyMQS27dFScrrx/tir1FGZbd3TfuVx1b6ndzKuwyb
fzQC5xARKYnOfr5ViXVW3ZGDEA7hERfMajuJ5mGtz2lJNA7CrNU5Ye7XJ5AhUSz2T+OcIxaYNxjs
FblAQew3hH98M6sYQvKVJjCYnuZzdh4K8vNG8uSYryHcchhV4j4Enw5JstIatheFgF0PD3ZJ4zOV
iLzKUQD2Boxc/SLAGBaEEVjOHZ73weUuMx7bqzaLbKYtLeatK33tU1FYHEcj7hNYU7qBpU9xQw2p
NdLSftPzsjJjzR5UNaLnmqywjbfhZl1698ea5qiWkFcbAdtbvvVWfLXAFlzj7TwN/nq+376uG8kM
D795b83BmL1KbcYIbbaN/+SBtldlI9qqqXl1PflbgnE+i6Rk+WTreHkyVBAAcfCiXsEB2uRRYtPQ
pXxeaRmp74lXHgXlAwJE+XP5k0k/zh235N6ypjBgYUpM4fAUghO9HnojihBhBeUdMEoyznKCZ1hl
XkXAYgi8VafhDoLWQGgAfNuoSmv6oPr9etQBK4gQKfdZtKfz81aWykCASN2zw7b9izaUsYNqWDza
Irs/S1LNPB1AiLuLGB7yZ0vxCTZ2NSY8QLD5RiulIaSnPhnzIbJqJkcgd4GHP8MILT1K3Dj+6lLa
LVXNynyn1qKG+a4no+klx6DPpwTpetbpQNQaoM0uBcl/dAu29+ZhSD/i6y5hrdJPLJhAvX3ctsXm
p8jIaSsjfV0jBHiU8BixjUzykmRPCbgAr9ahdFKkFj7oNRhVUsxIdfmOMnFYcRMGM3xU041YcCz3
f65Hd1JfYjGOed0FRsy+149EbYY4y8H/Z8tQzjjieqaCYykfjD+QUtAnaeLCLiguqXwGwq9gCin6
G0iNRoOJM509cJrQEWJDDgIVJfioeyqFrvfzR9+agdScyNVYZi2+N8a70Olx0voPrSzQexT2V/Ae
rGpgo1Yh8R6buZX8ON/7sKBwMaMF/TDV+w234cJO0wwokqS3eHJFvX6bTIjiHNkxtzLrW3Y+RI6f
CsYJBMcU/DGlQpXwg+wyUsFnnc+7gcC0qptERpt65MlHcf7tCF0DuVI8PjqGkcgP5SnroI8Y8DLb
0Z4jOLkHyNc0YmyHtgIxYe1x5JkCNtjI7uBUHE0RolTBm0y5mHXPTH/aPAAZwaW07Ob78fOvfVbH
+xD4GXqS0bQCFH6i0MFIr31oSNFxRGK2WFaRbtthdbSS/v2VtD+R49/C06VKFXmwmvx6fEboZEJp
lOjrkbu5u3t5Uo/vzG/umhSLmNUl5C5Qob9QEv6lSvpNRufx2rU33jnLBOQUS9930sttIXDJXxwy
m5CtfQQJbqiGPCk8tJNTrt8/JSZ0ha39UzNWiD9B23CKev4UEyr18kqralms9Cweq8eGx/UK9VY0
JR7UURcKMEkwd2P77Ywo0FzxTcl2Gcm7EoUl0TccPFyc4XCPTNMbymBzZ54/xsLgZ2i2f9T8AMzX
k5nfb8ZLecszJHuZ0y4WPYYoWCrTIkRxZ3JuK2Ag0DiLxrTp8UhjhxOsnpIc1DNMpQJ7au8gxi7R
fUMPCeIhGgmVecHwAPb9SpsPaWwwYACxEGGu+GwdtoYxUW4qfb5SoXZwuj1AWKdN0dmRwkr710JE
4w/RSZdjKa1w7hIHxs18BXpncBTkrAFM+ZA2lU/Ftqzf4OMtxe20bZMf7FpO26ppasUnP+P4P/b8
ohWdnf0OubN0rGa4dePMPs0LFQBW/OjRnR5igECFdwW+ykEAPgsvAQuhMpEBzF1p4RCOsIPM9Aca
wSm69egmJu4k2K4NP+E2lyWQe21eNTwk1xsfehizo0+SgUTUfmy3ZXNaIWHV/ovJZJM6qsT9gDUg
31T8+KAqqKVKsd/NEQaW3e1fvBXCrIz+7qaD4WlyzLoz+vIGRUmHNWTCe6rqJfgdiaPzKLeUNa3B
NgrYlixM+J/hY1ySL+AZpxB9kuzsLq2bAQff6Fxa+VxcKstOXl6ClHC3USuSGj1CJhUb0CcPZ0n2
VHFdyHF6dYpIFUYDEO3G03MtL697lPKEQVj2kV1jljwJWmp2V5xFh7UFo2uF3eWuZ1VUDeyI2up4
F90YgtQulBK+GpE9mka3f8tBzROVBaYYQbG9OV/OeifDA8NyuUAq8BC6PUYJ82aerXDsRnap08BN
iNkEEPXih9EDM9rJH9Qs5nkBwHXMODUwbIlMVoklBBd0l90A2BP/kZAJ3QP63GjvhcE/r9UutvG4
h292sp0vVr7DQOLFe2B4+eZPDAqhiV2MmUDrLg8hSPaAYy7u4cgi5E+XdZ2pEq68eAZCLcQbTk0+
XIfcwtDxS1TpDmGJky66cp/p+Yx05Ho/vBGUl4LRg5wmVTmSsDqn07tCC7GRZyqtBdKODAvvTHCB
hNmDWmOQZTWbU4N+61SrajgsD5O8jTFv2+jR+nj4Ux35HJ/iyNYQpfcpGo6ILId/yYaPSYzoQxBp
ByuZ6VlL21GwRi8rIAWOakEjhFsjgkEi3OmGcKBJ/0J4UAHY/FX8oNBepj3gquE3TzTieK3jJm7a
eKQIRprljzzVxEHBSW2RwpADArqvMOJ4k4lSdKpY2cec9H0b/GBko2xLSyszIBkAxVyYeQq9i8me
m6XH1RAzFWGxqKWeFQCOJKQbcehxkMq4YzwQotjVUnlH3BvXag/WW1L/WcVkLyD2Dj6MGiJr10oQ
DjCosiDpGL79ESgS+VsxNz0/dtGhQ6fwj4YPOpCaZQ49G5y/TjTI13PaTjtAnc8og2iDmcPnAT9x
LmVv8AeGKzqzVkrRAfpcwm5JZzuRINbrj/w64f0ADpO3KK/uUDCV+/39izvZQ6mqnLnpdoqKq6bM
loyw5dJiRVx2ledkkBFSV3cDsyWzNfLNk+Q07Qan+n8V8wxwbLmCfHJn6n+9JWlsMh83RzZjSyoG
m2MPbIWxn+SedwdC3O5gi5G4Pz5qtslLBSLZAZLrgI4UpmVODMGxbs+J4DrVVj6+zsj1ekXakbkc
Syed56B0sDeYFWpkarSBQhmU1KQkVNAc7EsDTsTFIpPAEobSHjU5FIJzx1iDSjFdU+MaOpUmsFhR
d3NhAVTLGym4awqGKN8DA1ArwcBcdSxCMOf6zuFd/INiLNZa+lrtgZIM5/mCwOpLBK4CMQCFIhh6
xX6LoObHpfTUCTcPGPCx8xmu5OAtDyQXZXmYYAvenA209WE2QjvUIWBbBjZVEUz0qZswwgIt0Zdt
J28qnZBZ6/Q1cJrWhzy4JW4PnW1vYmApvBswajn0mv0inY43/x8phmyCepjWlKqalrVUvpfaA9Vd
KOnj+zZf18Pr3y7cC0dWu1MRNZP7JEQc5bdY1qwgMmwtm1u7uuNVF9HL84F3o/3/0TQmgbLDTCZA
Bb0irw6O5GJUqDdNZxql7ET8FXWYwKmZphWTEUAp7Ak8cGgnibi0pddIKEb4lmesT6w9yzEcWXAx
Sm9CgMuUrkymo9ThTvJGot1P1T2X+Jb91GyQo5vQhu+NsYPm8cvC+X0hA8NOl57I9iVK6bdMQcXs
17R9D9DD29I/2xe6W13NxKSWjqTInk9KEOJfM4pmXM49X2dnaPTim8vC1+SnPVlQ68Vomqku31+T
5Na9FrwTG7ksP/rhBxcpMYOptTiJdAF+dccXTGRFpPOMHcD6GKUgemWy6dFhQAtrG2TKE6FfLv3Y
7l47CL2JhvpkWq2QkTIashBapQnSom0Lei458MBP2W+0n3HoECDClDDUkMngljnWWEie95N02Nkr
uUQqLAKfrqTe61m80UcXCQgK5EisIb7HRikCxZIUhODcxQ2IVAJ8kUy7Rb+g9Vg8HGcpclx7c2Zy
eMyS+3lwEzj6KEXyfkHXmIdCxkTTfAxUPF8PQSILtQWyizD+hKIjOgOqzshEkiNU82BY4qURhIFO
+lwWYy2nBOPhcDxdnAQpDzyQ/HRutdjSD43Pd9LFxbEiQseMGivqSINZXaTqITzMwkRc7sntz9cH
zkpeAcotcS8Q8+v3ohJE3pvAt9sWkfdcaOACBpzl4u0bf6spKPuMcz0u8h9tXLI8AXT/u6kfikdj
1ETBkw+gMv8f7+rpCy0rf3UOLLt/jZFBCrYMfB8800rwQq2+1+j5fRPuGEDryU/MxuYc7qAUq1FN
LRvMn+IOjtncstEq1X5HqolQBac95ZR6+Ek6IywiIm0l2OJEWw+d4OgC3kiW+kU96X8/+Vnir74Z
6TosKcBeEDLzAsCDH+Vvqb2LBQqUJbCI7kmTRHRC3pPw/XGABYOVi+w/NZ1bloSwInJiPjwEyu+m
3sQE5Ut32K53Z1G4mvE8cmkryKwyOKBDEbktp7iRUBJyqUeLwaN2eof0/7YifaM+qsxthgW0NZYv
lCX0unar6gU6bfS5pi06/DpozV3GFzJKeAxvYeuzqMRdO292Q7FfvUlKPN2oMuazuhiDTzCMb9Vi
cehGOYneOFpWIyGVXxKwr5UAaOvErWW9PSb7yqs1QuQjSKomIgDPwSsXzfy7UgV9n9WeG52cNIwl
QDpMAVodimpRRyn2fNLLAtYwID7qaetr4M65SL8NmSAkBPRLg2wDw8oEb32d2lk0Lw3Vs31KWN6D
88Ef0+3MWM9mg5eck3MMDdlfZPM3wB14Xigv5P4j+hrlbffa30AayXHmTmVNaA3IzEgIrxIV4766
pvz0byvtODgx+7Dk1GJN5edQ1HqjmplNZjNlXBijV/YIPzkzNvgWKKVjsC0YkhiyHvQoGft7gtwj
rnbJT/VGnXFEOYPVFTGeoVqq6x/xoSO9WxXjEGX59QKJjq0F5V1RKzDrWJMhLslTPavUkMlHh6BI
L194PwcWSQeoOaGOIyZvYXgtjgG+EYuyfzJ2yNb5z5Iip74u+TalWQCCsawLwPpaoYueOBFa/yhE
QHsF41WuRCBg+v2QGuvXpDAI2Apzt2WKuj5UxW2v0bLP7gYQG/3sQ6uXQD9d0wkO9VQMRaGKy5B8
XTHFjRBwe6oWfVD+AHESpXEArS0+ZZNOt5lOwk+zhid/b/O6RihFK0WDbiZ4fr0KcD+f9TRT0DBo
Xd+CPmfsT/FzTLq+qG1slT9E5d05iSyujvftE3rBjDpTleil+iq7zILh5OhbVqB49XLXeQbecS8s
jXMJd/uZnmCDRjWVXxELewtbOeP3n3Xt7aoAIXZWqeJpWx41P6DSz1vvvuLajdmgkHWEnjnU53l8
ibokal3a/hN5QjVTA7O5V3dMmYwSmqG9avvNjZzwiurqXJwYog2CU9hcUzir7NevuF2cv08+vqkL
Yqueeee5Hl7hymA9snJcA+01gzdcxurace5DUXHxV/JLe3PJCIfCnZaXeCXCwdqw7gmaZrgldbsc
sOQ4hPn2UB8jf7Ko3Ec3y0Ii3XPk5C4OvGLCQy6+x1Mr9BVgEScVbxGngYwvjUbgqQxyCkYb4tDH
poq+A4zze2D/rCc71YZWHyH/Sh9mYrflJt9wFO99ucoOFf99lEz1UkXV1w2Wa4vN0z9JHspkTzaJ
K973UdEAWgVZBQorD6/wvEtReHwVGzUOc4+097xWHuZHdVjOs9m6ief34Cl0Dtdr4AUSZcPwcaFp
2W91VHPbs23jLjAe8ola22AOC0F1vP0fv2loErGPRpYQqOHJQtv5EPudZKrxlYznTiFlQIpL8Ge0
Q2NyC7rsCrGoFNDjTxn2xUXspHd3hDbo9q5BiIKMbIcoRa7fSMcpuk6ulbRsVjxdkBjxG208Yekh
NQXr/as2Hr+ClT8t9XEDwe9faRf6qsubVKM9oJV7X0Z4O2nE+Yf5oG0BJmgLpT/gSlBA9Pc1NH1/
vyRvMEYKOgId8s/Je6BAnEmfA1vqeV476fYI1OLxMdTWv0Os1BIE4ozwpReJfihArukT1h8MKC3/
qq/9/qKln7UymIpFuEwEAGJW/t5f2G7xkNbGYemzmb0ftzUeEqPEnZjNt4XtBowf31UwopqCwrwx
dMux0uRGwWAsytA6ZJyUcEIH22lH1lUJAhoY3FyWmKsY+4/c7oVTcE2n50AXH+SjvPHhKi8zYdsq
jtBwKzjD0Nj0UkOgnfkTYL2ESt6qFdJmtiIeZYmBDL42nP2+E37UODj5hLvFPe3+V4CMErveOxOS
b7jaTA9OhOWwjFQxw+upQ/MXPeHMc+FPPU4ldIOeZM5X+L9AMrAOUVVEEr2iC05+0ayBbXKGEVLf
6lZqnKmOl4JGk3qWfCgoVWzSKJv6unMxl1bfrvkhkys7+UOBD5Ffn+U32I+P+4u41wA+x20zvuiI
2otlJMyLiG8n7ysdV4ivZf5BWW3cxzMwKgMs2uWt4usToqp3HFZYFqf4a21kuGXzOdovyb0NfB0M
TpftHEao3E3RgbR+9+6lN2dPDPAy9bYMxl9EeXrnHVaFaXQeRqgtpXzie4hvZwXEc2Fsez6iBlAk
t7yLrC+n9Hhg191/OI8+eo/rBd5XgijYImGLARVv19vPwh3CKLRJPBZIBG9/SruWbFILwI5VHOfS
kOf06SAGnst2zhAodH+nZkjdkAUe6yiHoP2Z7DEETjPYURS7V0lmSQI4WXBFTVjEbI/rPgse5Fg4
wjU1vrKyoUNQcA6gHOimPuRaAD0XpsI+J/HNyioJC+WWhYK9iP8YuJ1r5OtXmyL7wnzVLnhUoiWe
hTfQqfGiTxThLy0j1pS6KJpBioTPVRnXeZYBFuIC6lpIHefVc0gqd+JXE8mjhMPtctxsO5bW0t27
Wd9OCUc5xr8dOePhV4NpaeMdBNrU+Rx0GPzwsjoIw4vEPQXUqhamQj0V2h8/48Ebl6XpkTZ09MR3
5/GdIbTbY1NWQLgCSFYj9DvNaVUOCt1uIJl8m7d5p7N7NuD/dUluSUFRsiVDnuQ9GCQg5keFv+43
PQSp0dZQ3atU6yrChVVdin930Q2+tsYa+h2vTtILcTmSfrOklDkBqF6OU7t064BU84SH6V4xdm2U
LM82c/gPj37oHMo6TivS08VEys7Lhol8UAW294dciAS0SDOooYoX1DPbmdR2Uf5kMZR9J8C2MiPP
ys3wy40VYhvOzB0UN7/YK7oea4FYxZVByV3dffore3xFAGZFB4T1AY5xVGM9qd52C/L6+YqTO8iM
LipbDl5uK1H11rkTZVCbABEuimP1k6Mwp0gfTMwZ5S+XxXW5Ttz5HcMmJX+3y+Cb6IWXUR8+zpf+
XRpDXCs54+R4KwikjA90Bdb8ptbAEdV3O5DcJfZI9XoO7jVYZGOQleBuAiOiWhAAtiSCAyx54pJQ
mEa+AYglgtSqin20iF/u3l+6hAFxXwZrIErkbL6rW+Ijjh13vVLB7FlZN5WVWo6MBkZuXzgahqcS
k/Cdvmz69k/uj1pvPcGej+U0004pnVu/GkUdVpBSzZeI6M2dWgbwG45dGd/jL3onrHjXfXLCgqgE
ezSrCiyeDDZPhLgmqL7HbcPRmECBVe+xxabeOUL4pGXKjg/g8eIoVsa6dwqcGemBhTDFdkzf3UhA
na2kFXmrlPqDVXZPGEWvqsgJLMUm3J4YiHTfDc1oEv3i0b6+70ycjXewHs4drtBrYyjZSy3HvqSj
kwli/JYVrYP2nN5s9D/J1ZRdDr7oym7gV1w2nldJpsgmG2Hooz4og3nrpCrIXM9zdKJWcUeyty1t
RJROCshHBiGr9EJtF4bx4G50qGqRTpOgZwfEMX5vTgSBLadkaC8gEVRT2ZqMHLMY9Vn3TWjsJONR
+LKZXduX3Ncw8exg2LGhLC84uCMRjznNn0ybo6YUj2fkf96dQ3QM9jGjXkLeVdOKRiPUFimXnVUv
LT/t6ZJp4n81wyFtY8tyIrxJCcJGZrWcCj/IiAB1HOmoF0PBiZe653vlTCVpGZkLt7EWrD81KdXJ
NW6Lbat2s2S4oGupTn3RHCtzFnOvjRCMA1F/B6R9Sg8FSSfCo+kO9Zmy0qNV7uUNnI/7/qoFunji
C5RDovTQEpLj/YyfoTfqnPjfLAK//ve1o1aI7JxbvnyKgnhQdwLlITvnN/V8/Bg1Vw0Cck0F5XuV
2mhw+HJNY+p3MR7zYWJjYcbgJx6/BEMSg4Q3XEaySBiKQOdobb+RF5Z8mEyOxAagSpKNKjiYf8Fn
cP+SjyZfIPxle/HOEwaTXIaoSfMNCNi21jfNBUgUjooBR8Z6yNQ4m98HlgVEN4BWGkXXYg2N5PXd
gTJeZevBWMa2IWbgNbKiSS8lTT8LGI7t2XNtk4Me1x3o4QsDPGH4yMWhl9bTFm48LPxKL6tO+8v8
uz7VXJAYXrTPqhIdc1ltNurDA6+n5UeHNvHcX1m9wNLpH3Tc5ugHLXPJCLzigOkgyDgPVEBUpYxJ
syd8MFlsYBVQQyRXua4g0dTjEfyeOOArK1LpK27AGKCZMDWcjqDzcAmTAvu5OrFqdOu4Vn3n6438
lbohxEeP07AQjvMFgbnc9Zp3wDWiMNWVx43QN5mWkLel1oacGlN4TFruBiC7qq88TQ825MgUsk65
iLVw0tu4X6fm/dLT3mULrxSx6/wv+2nEpal0GMIeykhITK3ldnK15Q7/3Y9dcN8qPN7+1FbxprNF
0Y5ESVvomJCBFhYz8dG2STTQhEaeMpScxptFCoJ/LjOHPomXiHs+e84G8jL21HWZSx8r7VAybkN8
6QACc6dm3KeAIJ3JkbVlFe3C7gy9olPJuywXzC39Aly1DI4/y/iQ0a4hIjP44qmnfk/RXswhpw4d
GBu52NTwzulmDbBsxsdzM+uOSEdm1dFyJbeBPSq10mk1pkV3w+A5cN3lUVeNSg21sdrxs7smtOlo
bgHgCmgKweoeQudEv0t7l6OvxLckFWsjLNzCnBFvkClM3pD2srcYyRH6aDNaM2qZdPt/9coHAdMl
XEXGdUL0RBjkMT5WaQBJLh/+BlVXfleK2E7jyw+D6PKlgP6x/C9/htjTtp/hEAL+9vTVc9/cGoET
cFy9O6HydCSaBiuYGM4xz3Gga5AhQwzZkZ9T7zUPGQj7haED+G0jWyPjx1Zl0c8Y3OQ9IIIhaURm
7Aw/Yi4k/TIe3qkZhY/3NzjEtC27wA5T9RbmMUy3grjyP096JioikFm9SBjhr/cF3jhCX1o8GpF7
IBJcbPirIZIYaufcMJEa9Vw/Qe9AucB3IVoXsvaOYPpyJ7oSBNyAk/pdemsGFP51srnZo1/gMFvX
NusJPxNnqNgAvF8sz539pAVz2A554kgaWqhLEy16PottsWaGWfjt9qHv1mCKLiSwX0V3hf3YLFUW
YEMXf6jqQ0n5DgJEYYIOb+5wm6sy4PZ7vE8B/Y2OQpCXukTyaWgjliIZlJ6xOT46wW0xvOsKx+PC
Z9q8MfnH+G7d4CpR3uWR8t7aoIexbpJ8vuwTG1XCeRCzTjh2M4VWhSEQ0DHIDZvpIlqYCiNylqCU
cBT7j303HvqxfQSumFUE9BGe2FSy9Or0et5lD8bBJ5zVhLkctWJDmuaozF1iGLcacH/2K+7O/FQq
zAdkSEvpshuNiFgdrFBfxjaadzpG9Y1a/j2RBWuOku+EJ3XLM0gYAbGIR8UshK85yE9vghfEAcLV
C9k+NT1qXYWXX4k9K1pLNag+jP3RhmcA76EAjhALP6/qgFHn158a2Z8Bm9EYGnxp9LCt94tkzEbE
2VbHvi2g/Xk4OOJtKv7WIZAEYsuorkHUt3ec0b4VNgO1aThysUoRImVET9XhAZ95dFa/QfGObx5H
eOXwfN7kWh8R3IjZInTfoZkNFkP7aZe6McQF67xdPuLrkXLM1JHInBg3h4xuDd0ggjyYOTU7jeZd
Qo+C2SQHKYiKRd6DQQJrBlbb7Bp1SSGXMtebcRa+kb6sbX0ZFdkgKy57mGXQaZ52KhC49FzgnJB/
GCJOGWtnInKcCqS2NzuMCqR/EF58vB4NuNAfkaM9kPBsyYesNHGpWxKMoqeoJIo51vhsLDjPzZbs
AY5DRiPmmT+cKLJfVyrGJa8GsQUrizcwN6y3CRqR32bjMsoJBzBoG7nWj5buDFTVvd0fldmMlSPE
Z6fs3IOaayWvZC5lY66WT/a2GQBFsFNiaFgEL5tvQZm9+VAADl6qedwPWl63AchYlRoFQ+e5sXeV
+kl+eB0jII07wpbkfniXmBpnAscViI2Zk03KxeSg1HovpWc+2h95GxlkTQQdVfN/HjRjtPckGKOO
FsuZHklSNPUBWo6Q04uNsSRXk4yj2F/mIwHejafEH2vks5kuNbDp9b6+541z1jeqqqldEX4gixGO
uwGvQh2RujBD5GiRZeT5bWHrGc2PxcKsb//Kbmm9GPN6dV+OUEp2kgI1+GNNuCTfVffQ1vcNM1eO
+TgqhraT5qpD2/J6hs4lTk3tiJyWJ59uX2rlhSgbSlv/EQdKpzAmDejkjqZXAdAgbo2tBbvNS5Gh
he4ih4qnEfzglXWdtOTZW3TVdRZ6hwe6urmyJlwdE8IAR/YZsJTfVhRaHb1ffnzFHQEnDM0MdK1J
DyaGvvCC7CnRLEZ3aewvEEqjkRTA0O1P9tufRu7pF1aqNJJOwpCVzkWvI5ibbqpNq7Cpp9sskcvn
kjNsNMnIFtXJ0rFojsF4s6VLrxRgs4KV7puiVTl9fAP0AqP9GTb/qJfqKnys/hL9dBeuIPNaVkpZ
DmYhVA7yuEfLNFo9wIU72PYNvvC7EIDFahCHFvEZN2XxWKyluZCMhGwcmLvnuaS3wblpn2Vyl0JI
mBwfiVK60r3XHzOSb8x2Lx+JuZfIhRleukrn1LQgmKOT6rsI+8jt59bvjd0VfN39+pbi0p4V1s+b
ogPt5WaM56XlV/Y742rrakLO/y+S9g/z+51bsw7pM3NdV9/RghH5I9yb2EBHQTp7dT8dbSdYMH6D
a8LNJ8dtgKJtQJh4z0VJxACyWBN3cCkfy1eScnHgxzSwlW6hsWN4bLfveEQSYXvtgHFf5hJnjoUt
4doSflRcZFXfqLBeIcnyLbaIi6I3y7iPpn8Jk0SQN0c8dmuiOejpQH2ExMD1iFp1TtyR+VQIepoj
uYoUVidtfhYeUpZlm6X3LZVdMn6iE36/sqn7CiFHNnzhaYtwL49vyrHhAPPV5TGRBNxDjzVkdo74
pNL6crCbfWqUPtmBxVeKCHVY/LVY0IYhg7hM6Cg7/klIK91JXBsazHQWXJglJXVnpmSudLwtTQ9s
p6H11LYBIsKfvKDcpa1sroqbc5WkvndteTfA2bjrhUKKY7RaiUmVfDIe/DUOge+YmNZBwH590mDh
d18fWuztvbSmCHIYGioK3xA+PNOUs/cuicsrquvpQ+sENcisNiUUuHvWWT4/zq3cFWME/WjgOeTx
d412ivBceZ8DaIrNFuuZnJLspAu31gUhz9zph/XB4+KIM8S0WwXjdeS8QmCadZGWLVnKtZJEEyn6
IAl69YWKpiUcrR1+EH4NTLaC5ENVxshdSG6dvFpkyKuHxGhc3jPsOYJDH94mEf9cNSJA6jbJI6bf
UwpdlUffeO0tWih5/t1IimFSAt/jriW+VvzAMxRnML9qKBhDDGKxzoR62cb5EoyUagD4+6ywB2/L
bQz4zF7JnQY+UrGEez0RQXLecoCk8bxXz40pLg69sFBIav5vbDFkf4X1TKXsWg1hhsHp+Cbh29Ln
Dc3h5YLzIhpzJVIuxPp/QKAkTZJD/hBeah4SgKJv3Y7xDiBHUCQv17wfOz1uh+zKPfhjbHGQTaUt
PFpRw5PTq/rkCqOnCoktEABwhdYbApon5gg8OvB+fWlM1J5uUMmb6ZZyq6qbIvqllsGrWgX39ztH
U4PK5jfnXdptjsc+F8QU+FpvA94UEhvv6JxImPAXnsdrGa1+Be4gfa+lj+utrR0oH5jx6gvnUkQe
POpcqkz6857gSVmnCMrkQ/sv4GNCLtvIpapqOAw2CKHMOtpyvHFxgdLYYP7RKTl58XLwO92AKQe1
RURq6iyQdxgJjfyGgZ63iwFiGYNoizSfxhZXn8YQ0nWVCqEU+UOHOBqyUQ5l5oKLxWrNMIx8/GyD
+7wBlllb/6L8wtrM74t93BcVXajZlBqnn55qzPlhS343+q14SWtaSiV3ntlWLTQg2d8pRHR9xNlM
QwwbxWtQfH84AWEQpHaXaRyItg6/DS647XQUgjAKx4HPwGOhR7tjGSsOkLE6ckbLLQBoNtIjWW0G
nF+Fr/dAzkLXoDycN/AhP1aDT3KpmQFgdrC+0h1ZREBPvjTTalX7v34SrOnF04yrRRC8W0Mekmzx
dMU/p9AAL93ixN+QGXw96IhaAvnU9WOV2eRhk/CKiSLAqMgtUa/eISeoPp3yiWDMv3QsBcd6zKMR
WEoVACKE5XZ6UJDZHSnR/PEsg93SRng6RFNucMnvqBuRzj9mbO7noAdxX749RG0Tx92c0iYtVpm1
0tqQYS4HO1knkN3xNL1F2CBqiSwWqIRJA+UCD20B+jtARQjsNU4V00DC21h/LCjDXRfZ4rlPK37y
W7bZKj/NCzR1NXJyaYg6IeEtEk8dzRJCX/X2tDuTQrZjWnlM5dhpR1O6USsEZhxvG1W5bP8qxHhb
1IqoPsCx0h8A7hH4r6twN+fRj+o6oaWJxAt0Fy98WWWVSMTKsJevcwECZ3dAc/u0SUHARonM9DWH
Uq1rruOhTGKKlK1B004tMs3SilLCt/Our+FIdNronuKbM2TWIndGJFfcGoMWGWdYmKKVU04BIWeL
/JQE5/ZKJfjDOQtniZRCCm7RPBwC1Wb9t4rHIOGFtw9Nyc2AIfPhXZbrFVIW1wjlCOT3WJi3mziZ
WFfVlzP5N3wC7sXKbbb+2rrshrix0kzkbuZbWEYyRI6YgLLIzS8DqtTPr76A/S2vQLwqP7ZvGrKd
6/YD5YTYFdEz1kA6oXoCw2TjGJwC0811VYzoewP4l6MwsabxQf2H+KyUfoBToHVKfGyzyA9PSdLq
VMUIXllB6UfxUAW4INSxju+44zNPBaXYZ18j2vUfe92Ij8u0kzfLRK76qIcLzvDdg/u5cOGAGgNj
M8JUIU1JUGppXWn7jQzAioeu3EQ0aAbweh/J3ypcRW95nnDnHnVjARbyPFPjYLbn+7uz61Y1mfA0
Z19MWj12bVe7wL6nA/euEUqJ8JlqX2d68PcL9RrYdKbD/ewCyKQczKTZET51uNp1RBF7GRCxskRZ
tQxuu9gc07AzZ43Bsy7p48GQXSx0aE2mCj0ci8s+P5wcMoxOVwyfp+u2S2dTRcsRpa7IYsZgzfJj
mPgLED4IVere0M/39ZxA1sDV0mz+3jjRWckh5uCSIb+MntBvwcDVczykJhdKc2VLErfTlJGuI7VW
2wRUA9dRHAymWpWCc1rvOjT5RrDtXtDhyRfJKAQ2tPTi6XczhWszj4gL0SzOmHnJlMGuUI3wNSyy
Y+vuQyEX8lYCbuThCvhFiPugwXxlCD7+fNUsE2BrUHovBOkOHSDSZaxG9Id/6j1jT72LH+J0/AZH
lpHHspX95BYDT4z4JlLCh0PensIluxT/6fWntZqZmN4HC3XaENVfikCtRydEx2A56rnWnDCwPT2q
J9eXQN5ofRrWdfnwlQ/Ae8whrhQiu+SFxxZVqVIWfFDmS3gPtkQLMKxV7PNHG6D8SPqZpv/hgIbC
dmvMyvYeb6IiENwW+/9LwAO7ANNdzSvmAUXm9Cwwxm9YJvNCjtNIUUFtzqnVvjXNk3p52xDN+35Q
4VZ8pvYhGGjj6PVZkzrfBFAJweC2UFC6fwDwAKX6nClevVzSaAGaGAvTAwE2FJG9fZRBvRs5RDJp
dDAHbcvPJypyig9z7v41buJnruzdOJpxxcg/XR6qlcCqOF74ID9UhGb2zXZth8GEiGbKOGrqEgZa
MDyvgo9KCnz3FedPF6D9iF5cW/+A1caKntXFMR1VrK8KdE2smzhCscoiiI4X+EtC6eUNhEjlhIyT
PHcBY5nbcSwx0+jNuhbg5suzsKtXPOuTiK3oWGQkXSTT1PUPYev+7c5U4h+UvnrA/cbURnW5K2tz
jtIxjQkAzlG5xAUVA2+P+Z6vyDv7oaPu0TvzwXGFDsYF4U8x0WKIWOmVsbPiivRAajtjVY7GOf5I
nhFogrR3G1CVQTEUFEtNYcI6EOc+1DmMgU/SeBbqxPgP7LGHIWR4KQZ+OWvde4h7IGEmIJU54DZ+
b1jzo4CBmC6+iW5AalZX51L7K6DqTtzJRwOI7LEmtESt+uMCzkh6cMZYMvSWOT5Dm5M2fELjBMyB
qyuVGOtOPDYT8yuCgvgTit4PciWQCNdOr9+KTUpeYJKgDBEnmY/JCs4EUbd+JIpvI2jfzFWiWVw6
+o5pdPdYcj1WPcLR7CD/rd+IsgzJLrroktIUTe9uq7GZml/yzRvaBa+7jgRezl0AVvK+J/O8bMeE
wRDc4Vn7FyhLJH9xeWZmImXlUEeT2CMa3VqEX2Kz8rRnYUx29SR6BWmdwc2nOk/9D+6DFX2FZBwW
dNNfhsf67eQp5L+S5dLtg0/76Rab8X1fSxc6wngKvRwecGqgCfIUBGzejb5YiDGBMdlkdU/VkChC
Sq6BzPM4BMdhGAFZpraWpJBGeFiXxSPhWK3ihlwwvi5zPwL4vDqaWJIEnWffbNcYDKlTlSCRkyTZ
QCBtogcSzg/3TRv58RlQBB6C7h1I7IYogZOsrL+v3xMJCWTaY9SlBaz1bV4lDDK57ln0i7eiducq
gdK8J3iY+kjGA/j2uzH3+D8/eSZqUAP8XxypOEvVzjxmW+zBe6wmrCitKHrY+aoCAdCLb/72qnpr
vdQ3EosJokvIjK2dS1uM6vS90cbpBq9mR20OC4tf7BKTIEE9+0XuOkD7H9KFWbZgfRohcPGF6y2C
Frv3ra9stfLVS1bCLdfZ8JRX3lZo+YEsd9+CF1zXXng+gUqcD73Yo1kOuUj3JfemgnPo9WMgCqZt
OT4N0aMtzH7uulB0zDDVVtrDDuj5KR/M/Eds1Nba3YL/ipo5oAnN8qUzeg6nB7x593utjhAYvNi6
/ndqBAy0Q3hN4HjWtD2dnIw6blE9EkeC8xm4Wbglc3iwNzP5CSsueeOMbc9zeIQGMdxqSLJQXsGZ
bIqGs+Ci7rudz3Dpo6TGHNOjoNO21Kt7XEjF4bOnB798NPsmbqVZUl5a4RSQSu8AWp3YvhVQYEW4
vbl7mKIG39NRZuTl00NI5wB9euSUs3OpKR/C+GhC27w9iOr3MVaykgEsu6ulalsbXKuqgi3K91SV
lb5/NhhmsjxqIEui6KEHkth4PmFDm4X454QeJoMqHBchx9rza48QGzJzgGHOWYlaaiG9Vi4tWcys
Ab16AWibX6zfWvn2aeky/1yT6UelLvTrDOv6xQhW+iK5iJyxx89MsU2M8iNzR4Rb2RdHmLFg4rvF
XJna7dqQO8u7PhJXaS442obZG6HfFgubQvszuFyGwD6bAeKulkNkWoXRj5UYEMFPlsP40uLZ+gcP
5usbBIFJ1w5SEY8mUR9JZ3MixucnIXWRoiB1KInhS3VlIfBFYLp72LQ29A6hg6ZzJ9H0HhPJQ35s
59ysg++gSqvD0WYkwkak455+OuM2UxPD8czfwUSndNkI0B6kbUGX1zEGz2P0rFOVqEG4K1I3dE01
3pibDxdVs8h2XuMKHrqfZS+dKgJ5xPK9LH3qxHhe9wdCDFFPSV4fAkCnGZD/XpzFtftUy/Qy60C5
dDUqPgpTNpvuLaPi02eFJnxmKlteOMeVGiRniqvsd28k15ZUWbZNAl9C17LuqA6MWPGkF9AT8toP
xaYX02ZNPE84+5lW091bTyiNgO+ggEGJHHR8GJhmY0NWurV9UerasTTiKSEFXgXetMegcx0mbKKq
1c6i9nIv2a1HS+XSrCxgszBVPfclNgqyTeidhjcPAL3llexMQFeE05XO9x4GXK1MuZ7iyNU0YmCV
6nNu5CLqv5KE8YZvg5Rz5bFnc6fWrk+aYibLPYtzeBqA38hDHdSCAU5GXPm7V5eKHb1i4pWdvEZK
eot1jPzDssifKHOiF3wglC1pLwRDEvr1K9PSFE4WP79MFegOGeUJykLfcRpRY8wny29YUcrzc6wP
t9fqbfzLN7K9I782Qe6UQRS6c68DXaWWe6v4IECMLSN83RGp72KbDeYogW3Dr0o3g+2g5nxruV4I
pGKPF8lkfy2vKs/+LxnPkZTkrxLcXNNJod1F6/jxvjuRWlOWLDXpubF3Ke57LKK0eQzJcZZHMkoj
oZTIi/KsKY1+PuSZN/haXNNN2o64Z8QdjxvMiAGK0jNMxiGDvT880v7L6DGnT4v2sjuoxLXN+KlO
aFq4pnNOV8aX2omcWUVGRNvHEcG7BYgi6Km2VfWmOMEFrhEVmIM5dMbKRfBOzXi6ruKo/9ypOtEu
ZsFUBjC4GR1Cvro2hpDw7cbWHZ69B2y6TgQqNx7w81X65Q1zTlQjOnN9XKPR+MZvJexftQHJ3bl8
OD+AI3acI020h9vSlv7ImqUahN5dFzuVJJiGoQzGPXwEhND15mOh4BrM7GiHmijhSW6PtQZjiyQy
al7MijCMiQyc4Pk1CL52BWjjgSXu/LtSrJcDsUAhpKyBZtdupwy8jBD2/UFSU8G3QNS+ybLJ4apP
TMRxAJKd+YVFexQkjgbkmKoMELfFJxO79P0Zf5nwQ14HrhUEnee9PqunuIlZDTBhMRTB9EZsDaBD
fnclpabCBNYMrdquoYx3NWL4YTc/i2+A9VFNKlzZbmuYPakkNUd1El8EOPalRnzPv3+yvOI7gorq
m+kR5ErOFcjH1XfdMgoXOef/NhouPxduAc9LTL7cFH9QLElLSTciOYtz58/stQRCUaepMKDrDcpY
dixfjoiGYb7mpi+cT0cyMQ6k/lezmf5o3yho2ITMsCBWNyVeQTYP6uVxugbv/mdB8uo7GwwQIV9D
b5n/KFsnamxzH3vmY4FhZH1Ls4hLgONZYSfBPxdrw0TsEzQ2WgwSkoqeZlOgcOG0gOJ9gisYnFYV
TpZBmODEK1xoXe5G8indBNArkC7sPfAtFnzNJC6xdARA7wLLg3CHavjzMrUtIRlVnStmy5zF0WJz
8nPe4SPT8VkdxVcIu11MTkH9EJhbEsMRKBOWkNvvPiFzPxM6AVmhaLm+xIOYyUBBv7NRGUjwoHS0
0REFeo1cl7yWFMKlLL5hp5/GvyeyY5zehlYCy1QKLu4mubqrBG8G3JpOpXbKNrP+MoOWqIr37fZQ
/yJ/kRSOwL3z4eoKQBSArBh5KV3EBKw0ixcv1IJWShJMf+IhhxM8cPsNhgt0h+wUIUUAVwQsSVoZ
Rm0RrO9QjFhUhCJQOaAHf5qzX/vX77bZLYUcr9v91L8JxUB4LZxgCBoMNjisDxT09Uv+5JP81YBi
G2TDayu6MUaPNw7o3k9+pJelqufwEEQycQHwI+nyxuwJMmfYe5GTWmT9tDPqVkc3sP9Ac0Xg7aDu
gpSjeom/heRgV0jeqfvTlKPfiyIfmRkEnfB4z5DZe1Fv/cA+65z0PCbhUDojE+cQWPgT1NRuUxPU
kTzSBPItpB9JC48WbmBw4F6FBJ+XSY3HalVL+snWw/SH3Lx0jdJmDRtZJO4cE73TGiRxw34f4Ets
+SZZ+ZYnrVVWcqcVkwUsJJ3PoIN1N5zUbzibS/eulUzN6b9W/yYU+0DAdtfzlgiqDA483zK8tlUs
dkcpafWV6d01Ns1iXXUWr7lPfGLFDNAhzzS2LDIjsPqOlOrXNNqMdtBpWKQ0gyvE6zEL5QNE8kzT
flD15B6Fy8dHXHnoQmzJxbVLL4eA84OXWuBN/5AsIdNLG1cnfQ3yE/3jigUZOVjdhBQfrr9qmxix
WkTmgBgtFbXuam4kGoPzWqy+CG70Bz1NVHgKHWHHxGlW+acVJEhBr+k5jibfv52O0KE/czL5ZYUZ
2+TCrjdVL4W9+zTBE9vnaVYCZoBaAjB8yb+Gal/m8C8lk326KqT1ecWeSV/p7SplT4+LtqLkQVYe
wDyIktFVNYyTX9p7wKXWESjESq3KVfPVVt3YIe9SJ9WM+uNiS3MNN5o8x2JN1GIZXwMN4CHnGxwS
WVMYkpOg+JMIMMac7xM+moeLL5mzK3B/4HOFw1CTUiXGvUSDhAq3Rd8nr71QJi+8j1tmBKt8duNz
p6pUZgQY74ExWccpd4phRWClmCoEYujYv4wmzCMtfjcTXJSLWd4LKHtRsITquwkSwC5Vegf80Tfa
DGv8xRsM1PNOj5OkrU/O5TnoseCJ9zIy9depH+4KMj2j/xzDyIC2NH+wR6mU9w2mpz10o1QP8pi4
FOMGQtfqDXRPufOzKO6M1rEMU5ZwmlYU2OgaF5ihYB1HJ40WbdL8mWtDC+5XmidVSiORgKlI6tr7
tko3iycDWpXyn+QuNeo/czNk53tz8KY7cIDyGYc+nI0ABJKKST8PkN892+Mdsh+tDTaGWSMjrKLt
G/apRG696vfU0xTc6hKZJpZMTTp9PGCORJW4zj4kmtyqrjkj1xbGqMxUKuq4HuFkrA005aP4d7gV
q1AwW7SMeAUBaH7wC0WMw2v1xDHgACks5KjXb3Jn1i2WYjm8WtAbP3uy55AYrrPgwzd+Ho9Ne9co
XOR8f+IT8Bxb0YtRKNtvrqxxjAlj081O7bYQqrPIgL9oz8mWKfj2TF0PKozA0xg4NSS3F3SAo/q/
Ox0CMwvoyohmXq0Tb0yY5K2RnJaQItumhhUdTHz5FyC1k9Baqi0+tcrXby+z9JyAKfbFDlffGzvv
OzeP7ts9Ki+wWrNR0r3ZaWnP7e2ZFq2Oy+bB0LMMimlF/F2XDYvDEybw+8cTpxwrRBtTVlemfIYq
QhvdPG5+eme+wf1PHb/C+U+0sV7goWUgV5kkrNx8OqENrTmey2qmcd5M/HsCosuzYyAAjhjHNla/
WVCqaPgOgJbwkrNlHZA6p3j9GZrUnnbhjXn6BSXQ3qQbwMivAr2tOOW392DgigRsaRwMAMrj0SnJ
mTmbuIH2sysnh+YICD9MmiTtPWg/7zCyBk37MzS8F/yn/VQphqq1c54ZZe4f/4bOPQg13DkXD0ao
f/TSsy1FJumeUoREoCJLx31+BYhZJj/dnTOBO1l0WjmcZ5fuKolRP96BUCXMQytRE4yNfEmAIV43
WHfeY9/Dgdei590pqwxWwhJOS7YagCFlvzAqKG/ZkvnCqrIe2ebbmki1Iua6fAk/69lBwppPwKpy
xxcvtrBvp3rU26V+mb5HBt+klmiR44+Ey9RBl7dx3sFVOfn23RFgBmU1G/Z3qhjHFsF0+hAru3wJ
VCFdOz0TxshmjLe7iDMfgRz0S7aNFl5X+3KnuPk/G6pv6bXt7y1Qj/9Aqqzfh+DMiAcrzbpsHh/l
Y93vDCoKiXNRKOOeVlWkzSpW8bJlPTXh4R+jbjH+IAn9HkKHz5FKi3RusUcZXI0Wk+WwrrkzcUPj
+11QviLyKDIkspCytmlcJmG7nm+Uu8306dJZ8DZHIgUCqVYgr0V+LcuY/jq7frwBJihoSA6sVA2r
VYxicPe11f5i+/v+1dk2x8uWaKWzJ6nXT48xI9q0iKg5wDVexW+evt9ZRUR1A9LzkCYfNdUjKMv3
+LCBusWyrlKWIJ30bhp/w7A3N93DFDAmwfcVru/ppTB5QEL4oiN+ajLxOn0uUG5hYB7SEYYendQu
BmbVodPPpJ1rYoS2qjz8jD3V8ouaROxCPkuO0AZSiqePquY2y5B8pEmm+be8DCUXNwzgq+ZiC3Uc
gsFqudElBNHD6dq2CTcG6IsP7IjZSz/GYvXzn1eGOHmmxouaDea0mfuBJSb3gAMu7aHyJ1r7+FCE
nKYCUBIqcoNA8f5eXOEKHyExgSoTfAF3K1we5pSsZ/MNrK74YVy1GauGn1PnbFu8+6Px3fi99Vyz
KLVydlLfqHSshpeSAgOCclm/cUtcacFE8qV0SmCnLB7GRo8+otvXsKy1ce7AdlZtnu+qQNmTY/UV
Biu3/fXBPIn2a7kKVkiqiC2ZAPJy08M9PZvr/8kA0iEXpW9A8uFI4A66p+DTuT+iRIxYVEM1En97
j0ySKyiMB6CdTja4k3ejyI0bBO1fUpOWlxoEwTeDn0dkD1lhhvkYNbS/+BkjpEFno80TAVWOECfJ
VU5TuBxicmYE1oAl+XXvFocLUahXyZmtom5L52skI2OG30a/9CN1CmBhIy4sOEIGMdWmZbnb+ZuA
w+r0SkrVSn6/w+4+sbjVgwr2indTRUHDoqfNa/sQLon+cFFQ2O7UbpQov/gwDoyIG5FMjblazu63
p7S9WXoJ7TDuen2r5j6AkCdyj3jCScAEM7jjIfXxZz6AGkG6D9W9IhULHNCMII3B4Y3Yk5j+vWMw
iB/gLsnpdPisvAt0YLyqwOwmlsXcAhgru/7eAN1C90Y/qY6SX20QJ3rKW0DfoyHe//RSA4d2Az1L
Ao0dqB3nOGf3weyz95kcRNTjT/pivpBqXWtpFX9tGy9A3QzLHgO9gc+FaamFu8R1I6oYCVyck0JD
Mzz85q9QXt9+l2sRYHrZ1fvRdo/SV+onQ6S9m8MXQFMTa4adU4Q+esA66shedyjRWMq80vSgzc80
3vXMQO4jr0kJDn0OfEu/sxECk8HkmikPs9NdtenR4GVlZckaUkgdi4BOuGzPifklwAL+ewXTM6iV
chHOoCC61GSGze1i27dA+2ZFmR+loutPJqMsP4/TpoFTZhpdeB1H1yfGDPuLwlDsbT2uue/jkr0Z
IOqzFY+a9IUxUbavPZDHJLjnCO6VEtbA7yLKgy8PDf/QbOXgjJuXmEGTxHq054rl7oqe223+AFWi
pC6DLTPmDy6D0YdDtpSUsDw2GPraH8GLC4vikbs8JclK2P1zBiSkD6U/Dx4A6Rm9eq5CRSxUa/YT
zMIMolSXdn2l/cHmjrwJ1qTHuZUf2hIBRZzrGvpM6lM4s9mQmaoHJtPRqh2w6tfifwvmOVHEHdsW
GI6P4xVheIVlCy6/JHv9lUO8S6Ti5TyNuyTODSj0lZaZ1zNQ/Mwszzd/CJrf82plkYUx6TAf9ht/
0edPNhwGvo8OtempsEqTdCSJ91kfvJP4KcEPvJ8GijXmn+lwxarvTYWn+zkizYGuwVq3qrCFsYsJ
xFHrENQrXnd4vLsJzrnhP+xMjr5bT7weWkWusm+IyxN+UtuHSohcy++Sb80ZNTX5SCsEOtGkFfcp
jhR5chAhC6sD5PfS/HXSxkYsCMqeVepialNO3KvIxyUcPuTxkfYGLqeFLsQz6BTMynzEQIpxARVR
JgmoDHmF9f6/U6aeoJlhuUWIrQpTJY/JeRSV/FXuKafwvgZoheTDwrAxvJSyq/gLGnOByb3C8V1b
Uhlw2SxWIjHpRiTbeJQ/BTbOji5Zs1+YFTpVqNRQkO7+m9mg86NKaOmgoDplcxFo0yIRrmjFfyK7
u7p9eba1RplLPRKHCHtZj7QE4Agk9uUaBEzoRAox3KAKIVpSlwgm8lNuO2zqqQHr1v7E3TR9UNoG
mjVFDq/DaNVTVBx+X0LAK/9u/3nuj9/P+IjO0b9s6FtUs+PTMahyeQmkxunwCMqn+DMNvn88IQzW
pnURyB2DLxK3JPQwaw43s1qBOXg4q1G3Jbk/fUhiT0UvoTReSdLr8g0U6zN3a8r/H8qtPt7CGMTb
cicJhR3Y++DqZkvS9tNVprENVoxmazqhK23o+I9zy2PBrER8wqzSoI7HgEtWoc5s1n/mWU6V66M1
ytBkAqxj6C7n+QveU9059SEAtV8jVNbToA/bWwfrTJJ7BFRKfytlnsg6JAbCeMs6hawnJ34/2/I4
YqWeXGAw2OGupsUde1OApm48DUs2TfmHYuCmvseNkv4uX4jSXQJU72z/itPVlsVLxkIqXjTR1fDq
9EJlNMbteQCn6CX4XzWGzQsqXNIWSt5RjhFlqRqpSZ8XfNppPEU/KcY5WHcyBfxVGACjNTcZ6cP2
y5zOktvl0vjZdcQZlOaIyI8qmCxcdNNIxsu/oJGG5a9w6MDhhfoWkrMZcu0jtlckpNBD3/wIC1bE
TeSRHpJ4ertC03WfD0YKfs/FjhjGgTTksrgrncb3IqmeYL5e6BdUEuNUq8kDvGYSsHDO0GXAVCQQ
LXSaUKIvXWlDMIxYCYhOYTjgZLS0HIuCo8RRY/QWrjrqPJln1o9yv52vsz/BlGs3Lj7h+j+EThTW
p0cZfZWQ+6XvB6gpABFIJKvAYx/ETEe45B0ZZZMOE43eb01KWic6Ykg/iGaXLnrkRuLDvr4DPab0
iBEGEfP9iOoLPEoW9bvZaakL1Zwzcx+/XWCQBoYdyPUyXi15WwMKpM3WIyRh3OufPexM7UNLzwSX
i/k8mdtlGtfB3V1DBDdszo7C31CZSuzr/MDaBtZF00U9fQxvjwkTdaaSnuBah/r0VUuCDGUcNdj6
uHRRCjeeNO7UuifEvlugbLl5aDSJR962+oM23p0UBm7wFbT/OlSfZcyjm5nKGsMO+XLlHj5gYLa0
GLsfbZAdyGKgw+OESOiNmuzqraao4buK1rc/NzW6lA9JVv0wq7qaWFEmyiwFTNqHpjFS9woyVpXT
6mwwS09g1g2kbM6Ta2lDsH0m2kUxZv5/cIhCv8TyaeaM5nt7ZhcGpalBq4/+eGZ3ggoxtLSBUax9
+q7DaQkrVyLwhIfHzcVz7EGgKVXo8z89OiSR0/OgKrIl3uz5rEL73TayNANF0piOppjysBHviX+5
+OomybQUCKA4fX6P4FAos9DNcSBveVLHciTJmXu1lRyvzTjMjSJdAZvPxWw0MzLbnfeDEjcNcc5+
yunRbi+j12Wpmpp5EEBsgwqsUlxFc0S3oWYicgnppNB4JxjYIg2LwZHqRge7uq11vfr+/YmCqoZ4
6J87siGVimcFaghm4AmtiVAs4vhlwA4KrqYPVq+h/Gu4L3O1UdjHrkW+dBi7hRt8vmev+ghf0Kx/
emaZXOJpSIBJK0YIgXN2a5J12f1t5r7cEjjIzI944pFAn0jy2Sa2kQAp2VUz2yu+4Rd3M3kjb/U1
Iv8rXWQ/oVEbFOOEkNrdwkgLRe6MPAq0RRBMyTIWdFFADSi9kQq859DjpEguBgUK2GcSNLd8/NfS
uSC4TA1ZbLf8mIeFxhhw9JTDp3XZ2AynehepXLI7FR1QDLb3uR+xDpJaBh+f0yWa1z4mZLawVRq0
Uzh4u/qQTjswYUlwbL8vZpUegNf2IFOCT69HNJR23iHQWsmFj+EGAf+ts+oW8ZBD/TMoPLxcto7o
pyWAL6qjUPdWs38ZDxo1vkBFCjBerMWNwjDtcmT7+mfNDRNSrdyekcSkeo721ad7Y+nQ8fzy9iHA
kDDtNv1usXlDg9tqqccmOXbHIw+B6ifMh+P2zA+87S2dvDapJ1VvXb4OCq8Ho+ID6MCgf/vCNzvj
FkP75zF/CLv5UIi5E98JOWro7e0+YHeFuOWtCy6QmkfTPbexBoG0O+80i0rGenG7DzN5s5cvZPrZ
Vsooo0YgXMut7uC7x0w7WuFCJSxiZdTKp0WV9hauq6wYgRzpFLtuW4weNMpjsyihVeo0xGNfYlLg
Y069cY3aH1fXQZE3DKbZ0nsYD4VAhio2Cnk2bjE1Hip6oIMmH0FH6mV3kZ2MkF3IUZZWl6I3aQUe
V+P4dVe9R2hr/4pBNFILIOOalVblhkotRZbyDD/C9hHtXKR8HS63O2JlITy9ga/SXYc1oHn1mhs3
Y56bMurw12EuwXaQg3zl0vkLFCw3j3iWQpnqksO2KKHZuTrzEiA42i/KFGqqF9uXlbkw0ik6YJRq
vUOGtY8/DyPO3KL2O+gI6cYH4DerFhA8NzcUtRk5V3aTAAhY2pFTPZvysETRJYTqJlwfe+VYoVgG
aV3SpIxrzr9MfTZZxDntcIF34rl93x7wrJj9Cag7t0AGqPj1QKWXQb6wluUKdxymKt9Ih2BdP4rO
6MV/Fcz1PrTZky3YXos/EGFlP5adJbmNSJ9ekVLc0099EHA1Bn+kpHNJtUlQMjnbEFNFDiD3Z58P
2+xNpWdd6grT69UuagFeqQDehTRnfXOzXXneOfmyeX+KjaJsQEZrnMjqEbPbeCb3C3iyAZeR2S1v
bLey1gYB9lUWTsWgyPsckuT+mJxI+9k4W+WjvWl8nDeF3U4/RaBbib2hNYc7JZJQbq216WYhdyl9
o/gUp61NYhy6LS0UiKwdu7Izf4v11WumXvo8hdZfSyWc4LT/wic6CZq2MhR7NCcDs2mI0T7vazum
x6ncKzt7SG394bO3ZylVH8Q/9Ful31UNIjOfuCfdsF+I4fIZKIEyY8egdl3Wz4qEG/lVd33Qdo9s
Q5cmsqKHNEZyWrejT1KB80CzULest6WlBj/O0RZKiBEBkuVRXqyUyXpadYfw6PIagLos4/57OGaO
Tc1ilGp/TSesifJKhxskJ7vZt91qr9RKKb7Kc0l82jd1M5Bgv2PsJ1+60qn07/0Q5YiOnA+34gwg
9TU0zi6TPtas1Usf02ix4xrYJqw2lNXXXVAP4uJPKbYB1UmNEy7lB6nBbKgcFC33On3cVcCsrS1O
XibNd0c+CqxeptWSnd+zFmvi0FLLYndDB2QbzB2FCr6e2E+IrGcIopOmeFcBYdH641qjqNjld3uZ
zI89jEfU6pRthQjLeGZmPAHuKynm3lYPoeGrCAHhPrG3zz0c1XwIOe1fcLSJQqNGkKqwvuC0BpRP
EUraYlGXcv31PhkS2OmTIQJ0o0nb5QZoQQXPYlAJn77rdNcHdI+9C+HRWRp2wKBmsMGD9RrDZP0W
vPkXqO2NXY5cV/8xIXXVyQfgdU8LS5gPujea8KRd/v29VoXep6qkApOTLWhLuK+daL9WCznoLH4H
EYSKykvZLPCPAb4B2D2N1XB7V6qCTsJU4MTuu3hZDn0TA+hlXw9NY49C2KU8B4gZ9Kc4Z8l2HQis
SI+NU1bqFfQXgndk0c2YIUJkanN9u8qrRxeSYEcw3jY3YV57b9gmUAFv4yxJM+aZBgw+Fn+wQ9Ik
r81G1edQ7ShXWquB6umCZ1BbF92jfj6p25yNSr40b5unnuLMIqG0QN/YaD2KxmJIl3O3NWa6Zhf/
MsiI+oQIFfNmUSbfQUoR0/flHrtplwhkgs1+wQxM7iLQGDj2Q4/mFy+3Fknk/p3yDLHzIKDbuNGW
gyMqKo6sR+QfCk3woAMnxpY0x3gkDnBJGsSK9rHdHv6hXpPrB1G0jLoleiqpXLyt394uHcGYwGXI
1eO5ww+C35MCjKSxrkoC0CW7YIXw2sNAMbDaOB0ZUcKw2SoLTSrRbbYM8kqal5bAaXIu4uDAM7b8
RA0o0lXQVzzan/3Ho3NqlmFJSYl7y0aepPoBvcXHY/uueuVfdNdWeVW4Yh42cW9FklApVlTMD9ip
t0/lmVx4rmlwgL1d89HUEM0NKNyT/wPmcBlXjRmWcADkduHEjB11kfW2voEVz28lLrQAuwNl5VL7
eKFgVwkOwFXK5Y1C5EriUyU8vqLobPT9rWEDKD2wM0L6w/QLGN1g7Q67ylvEtLjRLx8zOYtmbPyU
dAImZS9z9add/GAjLixSTfosSKzJRaV3FKOJWl9+5pONg+xPS637v2bZofv+fN/XyVp3iW2OoEMq
bHqhDZCGkHP4e7cNlnNXfDUlFh5DgsMQuaI+w+/rnwsU5WLjZZv+zqFVNt+nPaYdQIQlZQVBKo83
iZUTAYFLh7TGBV8P77EtZavccWPLPKIRfiSmEFEQCz5o4DJFbL8hVQNiXSgsEasXo7wHYZ61wpeS
MKbFTHU6PUKwVsRq6GTDsuEGqSpY341qyVj8HUU9UKmSVDzKRhWyL5juRZvJNwD2HMgJI3GPzsiE
x1pjns0iFnB2qlKpdVi6X68/v2PT0Ys/W7SF60U/WfxskoNk6eM4WUtG1zvo/SB4fisXAuYRtRwE
NtEnpdowJpLC0HtT13YAcJzCPdD/1vqrW8tpQjjVTl85w49Ba8dTEOIiNzlvu5Ol4D5VxmyMN84y
NVlzPMQkGA0XcbarhiYhZYVal5kLvpqXlid1fzpkZAps4RahgDEJR09kbFhyF39JNeBZtaLuu+L3
p+CGy6vo0K8RTc6gxlMnJJtvxr/nBbmgYF0EMsLgJTYmz8UH23GIvvHOJWEsZrbRbxCP+Ue1NLz5
MA72vXqI7A1AthttVJ32l1YScuFOnp7INOSVqfpUBVDKLgy3ApxeBWf4tuXEv2n9nIqD8LFaS8Fl
4g+SJvnXZT3IAzUY3k2BEcq2l3R3CUEHcJqycp05I1uj8VVZoDYUypO/RJQVHmNb9ql3P7C8ztiH
gNp9M4VTRG9Ndw1sd010F1Wfw9kt56Uiz/8hps+vaj+yNExXjbRClU0u63KrHy4WDwUFVgP9ffSk
TTkZloFczEeAz3XkIZWYwc23jbGxl6SysDmHMsSzE/sjsecG1QszQMGZouLrpAJW4UwspF/WdkuM
1woaWQXxV69HJQhT7Cfq3Hz54UqsQ+AiUG1VE0ZwwDDhKYXP3Vq16TxgIQZkUa0p8gwdhI58FNnt
NlfbyxekmJdZKauctH1P7SFuBkqpLUHeTs9F7U7mY0MxCQypLGJVj9xdHxRUQ0ppoOXyFwHYrpv6
g5q7BZZRkRM/GhRN60BXnyOUNOfEK5KGxKAAHP+6/OIcnhYOB4pHITmNAnJjIj0vIUQguV9MYM/P
pJNjQESfNU8IG91I+MrcNVQRz3qsNpQuNHnZ6JevthEQl12XMDAQFeDN+OTrminBiWgkPceoHTx7
Vk+YjjJrWWJ3PsSvTCDr2CUeigRCn+1xSfxGo2Jk5I8LFQGFJEPzpLlCOEhCbtSvLfqlCioKjqGe
EGd0r8aNjs0KQyzuRkTxbAB7MGfloBgGOqPXQ5+Dpmds0FHvkY/b4fmZBeKDa162O743X4MYsbQE
8cO3r1l7gNPl7M0tpDpZCkkDPdIRAC3kOXsfYid2WVitFcFjiH7ZSXgStKOoavOXefC9JnvfoW2I
fwj2/1aeAqEXHSL2S+26xT9vkuWnxrEajKm1WUGfZhVMJ7+HJgcje69Il7zw5i8Y2VdNYGDyQlIc
caN65kyEmJ3+zBmauBbJgubZXXzjbIAfi31KaVQuakrHBtPAM+PR0XmS+5UW3N8rRl7vKO4FDS1R
AiBlull6c0MvPlsVcTwePyybVgfMMm/S+8IJfRr3FeeVo6Pl5xmFVSIwaCFYZTkzGV1XFYA2+S7W
3QZFmpEq+EdBqMyZoFVsh2N1GiHmO7KPK57NzmaC0RFFOGJmw3P9m149YDj0ORqFvK8Mx17lgwyZ
WR9gsJ/fbzJ9cs1CrTySr/fTuLMM7aRaEFBkq/vbzi56i96Fj8c6XtWoQxsQvjposo6d0yONJHmQ
1FwfBl83w435S5gJKVXZnCR8PFUQ1R0MXzGt0GkKEYI4QD/QsvKb6G6o+/Yc/s8LoZyTcxQvRWno
47Sntv7GuSmVrVq5IvGBX2YTVd/sfW4PihXjGYpsiNEidLAe+RU6rEt3h1D1/KZaE14gLcPoIOyn
wlcBmSrJ0QprujAi+tBfqlW4cCMeDtrjMWVqoiM94vSTtIQ/w8RKM5lWfzU3EgqzDfuR/QAReNix
I+gKpLLHq03+8q3e3LqVsxOcC3wcAfk7GjTP4hIO18BeeDuOCM3e5/R17qmlxdynLpBp8akMmu3h
Wf6efh9/zmAc3g+ugqu2A8FXqSpBU9+PwuOdzlVBzZx2iFnwf/xVykxmKtysS4syE2JPhL2HgBHA
Y+31qfus5mYRDEdKB+BsqwsjgysLVJd7xNz2/4w52/79cjhd4zfdBmDdSx13Aj+gDgRTfBGZy42F
O1iaYz/5e1IxpRsJTia7WXO4qkyQzYRTmoxcP+nX288YKN7KtQEEvU3Ktg0MZdUn/1VflP4eHk25
4khLFrLC019ZzkoI85/GlkB+ZqiU2svog1bxM1o8kYuVrnWTeyPwKAgLSnie7cW89BGCnPwZksMW
z8USE7FAN3tDX5TsCmvRKu67q5yxMaG56+2R+zFlAsQj1wEDxM7UptT52YLRrmUMmqlcmNfEjIC/
GNtoi7W6USryw1VPYB+/vHSuQEdBzRhuc+vZztw/j6kdBFOViEvZg3v16bfO6MfxMhQ2Q/H3oGaE
dB3gKNTb1Onx4wDnFLUnWDMNR0iq/0LprIrL68TZhWoG6zOqElQrHiBweFTDk2fNqLm5NOgMYS8G
DUvsx2nJyL+ZXvaXgHTHPjPsB2s+6tKsA7V/X4jfg64wGLKXrdL2caVyqvqWtsZKuhGbH+oTyYLL
Qy2zLFVsB6vKXbGns2JmGJZjhDbt1j1qYicGO4wKBe0N64p8TVjGJcBRqWogY4ZztPetVvOLlW2V
aLBs8spyCdoSRa3plDss85z7rkJBueOtwmLQuDWyais1WKH4mn8lI/wPptullv9wqiH+W0iPwXDP
8513nGGIjVGTdBO09vwoKLvb9hAJse5N3Y/lYPeEsoKDKrenwRemyNHxIzIOM5sK4ztGXNEQp8s5
nWtn1ZE/x6djVT5JuVpUf/c0TbOORZca+Lu+UBZf/LhPqTasCkvPLCdqLj2mKmq0mQ06ca6sodIb
NgHmUMFgd4iNxlMi5xwm1swZBfZxsk7jSYTqJW3DTCPQ3mAfcbO9HxMsEbjqEDAMBmy4YkWT20bI
LhfxVhk/HBGwxTx8PrTTpSnP8eHfXk66vufJwwx+jNdxt7RQ9epLVr2kjQAL3Sq68EpsTWSI4svK
SRpX9aZbOiLa07dNWp29VwUsPmLJFBhsOLezHN+eczYfk63q8UkA+C4NjRBxLC7hs5Sd5VyrnpBR
ZVJNTP0hy7PzGlz26K0oOjpuoIeDyfQHCvzxmhCoDey5Ob6PHGwP+qA4Gss9MCTR0PeTnMF7LuPR
KRSQkO2NxQdMtuyicl2DZFFbJfCtVqUb5KatPiZkg3OTr4vT71hK3qXl1bVOi3jq30vaUt9/x3AJ
cYo3g73uUDF2J5vF8fkxI1EE8hIFiQBnsbZBY1RcrHEne/Ojfq8D9LO8fIss4pe0ZGeqmG4I3xej
aNbdOdvJEeoFn4L7QGVhEuKzGn05eDRDkoMU2Rb923vrIUaCho5hQS1A8m1DQg2eXenU4RThAT4C
TbIGz2SE1oDfh4fOcxIMMB2J+Nzt83rW9Q6pxtJjSzySH0WmFu3whqwHOWa+7QSFjyvTlx4311FJ
2IjEQvFLWsvj03l4Bo4YZrzoZHNw3mV60wlrC5K96HvsUvoxKOz8D2JkCq95LEDhmMs+N/0WruaL
ACwBZ8XGhMderMtoTQfqeqg6W996yalVUHZi9vWl+4bQ01zklk/rAgCON6G5A1iJ9Kpy/Hw1sVmH
syUSA+4QAR0tLBz0n5u1QTLWEb6lvTwfEEQqC0sfSE8Xs1c+QrV2q3ReabkeDRiQ/4yYwrcqHiOk
Q4GkxhXyA4jubFLXjDHf29zh7dS6P5OnkHeVODOuHFZw+muffftaRgcXKvl832iO3KD5+HLuQKSv
08ti6man0sJktTRpOlMquOe3WyxQvv3EaHFjOMPJV9T3EGGl6H4mpq0aNQRr3TuSJDn8qi5khfww
p4rgowx1EsMOWsVycPdmTwl8B4RIJSIfsWspTD6oP1kr6hC10hgXr81jlMQulEiyuhOacyhU/Hql
izr/kUFiOH/7epGg0zZmcdIOJ0q1uA0X0uudgPrnh4Vd70WHYG6yKotNlZunon3ashwCevTh7y6n
xaV7fEUjiKZUHzhqZSjfoYvmRlE0swYbpq2yMT7Mm17duG1FsG/bpjAR9j3zs4ffIlpNnkDVug0i
u5+7F6Db6YB32JkBL1h62q6SJ/icOfcjeG1t+SIhWJApRjOrBqQSMNzsAk7B6EuDNqWiJA5kjBdO
/jS0+Y98A8orCSCbMqZRm2XlKkNnpBJgBHwJmjzat3EnPxvzjjMxz04QsV4FQZlkfMaxa4V/Ubq2
D04CQYFZSxyiOrSd2hl4F7ZfgFdhBKID0sMsJosmiV8/Tx0nKel9n7/6gNez44wINyz+ReSN+Xdx
R4vylY/rnzubB3mnLLLt7uD8jUGneBYJ4y5BoGEiGCzx5ZlJVDiDwNsBOYJa77ZQKPOAQa8Y/9Bt
sFzx4uxzRTfbkIVVbFbW2xAur6AldG2WJh1xJT/BOIYfUvLBT69r4D9aAHGjIQWO7m2s+d6QaokJ
fCVTpaL737zbSTyZosQZiMzzs5wRowbHI0rXmrtgdgafuarCa0toMrqqkNX3rJV0UaCMS9Kho3n+
McCB2nkNp/7vkWwFk4m0LVqijiH4LIL88CvvSdcgOJiPgUcwnQFf6UFkps92gWCjVngMmHZvAq+X
9um/kYKQSQ0ZvrWOEFGIsAS9gNxZLFsVkpW56nSpUcZBfdZiB6XU//IM9yhobSOeRxiHmdSCcK9m
k1+gsm3pcZT3liPSaVSn0pQIKEJIwxG8XB2U0mpq/HMwimdfqWl6zUgecnNrtqZwlWGd0npbNu+z
D9kTBJ2rp6lnv2GKyZ5khLt+FDH+FlPNkYttmccdOp582whR5k/XCazOrJCv0fgOrZd8e6eXMWNA
vDApPTnyGiOvgzBVdmcBuiobmAHTML1vcoMTNahgkinrgpsV3vUXbVzLrsgRYRmVp4AZa/nk8fwQ
RK26yhVCV0fFWrNcqt2qyNSpEQVatX+81GByS65iBHX6nN6W+0/avUWYi7glZ9jb+mYizRqh0no8
8lwb4ZZc0pkQnE3BqJXJBE4ypWKgpzCCs9y+DtE+JqnF6ja/691BadophQws6TnlAC67TRE8JKvZ
FNvD/arY6l+pPF77ZrmhX5PD0W+aDsFXCZwnDiQwQje0B8UeMTIp4yqbxFgh+dG0Jv6GylDfX7t/
Kfa3G2V6HY81XPA/RzsVldY8OCs5/SgO2UJaNwxwq20WjhFXtKtFR7Z3ZWe3+PEaDQ/GRdztHXmY
+7kVYVuQ4JrV0jvYEEs+f485M+7x9yzjRx15FJhpYzDmYzbzOGNViJOTy9JNvCIJoV49Dkmfhoz2
g/J21JQrPE37h41d53aMmwxDfK+Fp+elekzFT4CAXHIddJRYlBUM+uHQsgnNQj5d124y36b5802f
wYJgD5JRteZEOkxSylLrBL+CBWgUmpMKr5LHyIrs2MrrtyWuieZjtMUwAI0m7stCFIFxTCxFb/eY
6BEPSGx6JHUXC/cfMJnSo7ywV9zRhAG88EsZ/+ZiAWGhNOP3ajm/xuAebBOd/VCYJbArgbiKakS1
1jLOxm157mhBw+WnRSXei6IjEJ9nfxmRzSuDrPIVAYrDK3GpVydqHrFDL8anWVpP51gIc9Fkyjcn
hIc7tikqMxDttNnWGqaJWZnEpe7bew+Syw8c5AXxfGrKESN8Ng1roTEkCP2mLEKZPPub4rWXCZd8
TrafzaVk/TKLd1vQvfGCCYPZ4deWGPv6p06XHPBMmQE4WMlZNAcunk5hk+Wjps6OpJNeAMfbTXio
MYuU95Bpgei/4vlV9Nca4sofQ/DggA878zKfD71LSMQSNSPzX8CP5HAT/CZi1VgjXT74/JYMEpvS
us89OLuuZlS3D6VYk6EOXCfyWnNcgNJUNsnh0AWz1dmNQ2P4HZGEHiTsvGqf3P+7j6DWvY0jVXti
QNYhqCu+JaAnFIlYmjZ+ZN2TaKrUpPInV7Z0sNfsfCLlg6xS5BxnthvxkEDGJhl368NreLVj0FZH
gJbSD6Nfw6hVqEW5Ug+gB/Nvps/R+4HsFF4nfc/YzSntY+IT9CJXdOUn818QlCp2rYsj13AWLqUn
F4OKVL4IeusHeOa/wwR+/DSVURfZWvGp3H4fqIzRHmqZ2rNU60Jcbtd5cdWuv4zlnqrA1bNRO2cP
U8KnnrQvarXJVH2WmEi6KLdLzJ1lyL+jgKPBjWoghJoJmBahGNu1jyJHSu+EmyiSD5ZiH4CieO+m
V8Yhg5nI8qUq3YsK+oui+T4FS3rw/yexz4YOar6X6Qcy3oEzjNn9WB8lAYjdBQ+1E8P/We3ZLc2R
F9lmDKxUEoZNpfKltCnSwTNDdx29gupf/Irt+LLBUmL8T1DJcQflyDj8acNf68URrzD7MVuYb1/M
a2jisUrke7qzsPOTxFbHb+5rVN5aFtEhMictmCB0yIHsmwF/IpIisrqO7V0OhKdcWeQVV3sEW7US
NIi7biMZfrEv+exlCL69jk49T0nQaCOaYxFH5qDw6rkJxo9IIhNr3U+JL97E/YEBp5R4sTTgj0xR
/Znv8RFqx5Q8hyQaE3oIyQ4V4tCCdtamfCcpIQIw/RwbmBdB6RuBoc+jkpNbHE8fbDcQGgYq7gt3
+9uAuLcSZWW+yqhWphu9sF0Cw/obageNsT8N3jojdztVYpQw6C/AZJkqY1KMNa3TbD3j4M+uaYFp
yZvvSJR4hik+Q/tNl2TxowaG52sRJ4eF0bwgjnM74b/q6SiDt4CigniR2nfXmVG+snOqJ9DDyILr
bJLJkHb8A8MhUF7u0SUnRAuyG8w6YchEP2uXsDj1chho34K9OwPshOCG1wUC1873M7XUVgQE0IHP
jXS46F1mFOMD0e2DJGfW8upajBgVUdipF3o3XRHWvSNKEKe8Zbx4DulGnSttd3puxOLiBZ1CmBut
HVY+qizRrzOHWVi/GbV9kncJit1jlR+coqvDfrz5MgGOal7rnLX0PL/Xl9c89Q+KgFl7qBR+Cf6a
6ayGcjuZ9YvFDde1fCb3tWjAgq082Udzl+Ju9m9vfsmLcDPdbwcpq4txozqW8hdHO8k/napRbfD4
RjFnHYt2ZG2x3gX6f82UbaIxOJ1tFzXKsANh165K7GuYHZ3NvpuzNg6O5Vu0A5NZo5/DVY6kf3v6
mAdWVWnYjNCWIQZbgD1xvzwRPYQsCC3cffUWoKM/xGhpiorn2GZmpwV7gqvbldmb9cTtp66wbBr3
xCJJ3Y3nfzdJHrE99hPPuoKYv7Dutt60J1HKf36m582KLNH3eyZH8IHhE4FLc3vi2UfED8t1EeVf
LT4Ku5hsoTMoj+iSjEX5Gz2BmR9uVITGfrqiFgbXk98j1jDkPo2rOIWF9Wp3u2bR9TZF9bE9FMQf
WdbP7dfLeFJzdBdXRA9/MRNT/eiUtNOp2rPBplqFq6kvRz7GyArISCi07kxkm0nvZAPPIA86rbkC
m67fCu5DkXGvN36baY/6dqHeIz2QfEkQSUuBT75z2+Y2RZBINS1dW2n585AiR9oP7xhnZ1yZTdEU
6EajeSdOl4sNuGAb3nY4anubUOpFWi4eC+6ArCrqb+n9f8ltycpRFep9rckRLmuQyjpr3XLmVHky
DA8z4ATO4ray5zCAI1ujqPwR4EyQmeM/jrntOZserzYcIbj/aJ+QMu28e+Z+3efFeaLjDK/Acpcx
mRXf/4qrkM5l5/+qBwGS9LGkLjde4uY3Js7cBOTJ2tpyo1oi919iTPPNmAGiOggKHKHVn9+OXz1c
+QzatahvMUq07E5cIo4Q3HIVPlUYGB2ww/h1lkgFLVRQ9mC485Gq/kEXhsAgoqdV6VyoT3vXqA5W
LOjox6TfMElLjt5hRvZuz61rcOes+eG2Y2f/7NlTOqQIHgLxrnB3vFGzisyW05zhUzP7G1w8hclO
7X5HM2kxs1Ut1CX1U0lSBpAI7+Lw0G1n1G1MqrTCmLK9hcDrE6l+g6TOllIheMorakiJOVcVKGiS
PYeYo513i0kMdQYBPqRXllRrZUBnqn3zGtOFjB7Plbg8w1y38z6RIRRWqpVVfVNVU3hOMF9FEPd1
bttFuJ0tKj/PCHYPE0/sfOKmaS6wbWckuooAmE5gRC0zTIYOJEwh55ow1rIowMMDp194lKB0ANlL
2Dcb5P/gzYnWtrA7qBnsuydNFgjz1fJQiEbD9vePX0wWtzruloiLYyZXzbEGwCtZsiitvcfm1jte
iBOKlZ6WCD1sfIHkp2y1pYzMIRu8yRFlSRMSluTcJBEYa7+/+wqTzB19/iLqvxEv3BimFfikcLE8
QpfH2X+omcVBaFyJyPm17eDQI13zVXsPQiY9QGIs9tmoFNVAKufJGmqYPaEeQeWZZ1OgeCmLsS8H
9BUxCRNsMTYDqUOH4ZCOh7mzUuC0ZXlMGoUO2/6YYvQMKLa+5d4pcghsAMK7HSE45DXzub2lHQAz
BxrWOvUjHYnnIqRbGdrY/w3/+fPvy0I7HMzZ9TpU97KzvIZeHH7SRsUhB2s9JzShHwRB+UQTsIG5
5RKNqILNGOOHunXnguAKO5q317a8BfBuJnJvMe/QK3gHiARFf7rbcOXg1hLXL/SdInfkm2Pido/f
SU5DFrQW+0AoClWEhm5EgPryOCUKEVRwenAkOnJfxdDc5jkMkt26EciuCs/HlLD3O+jR4TbxosKc
uINgGFqOjwa8Q9/Q05+JvQxRxPZMLSO7/MW4T/hweo/uhuAaTt9sY+oni3/R9s7d0pLzhu2JsQbz
0aWBL6MSLgnfQ6imqil6OfMWUpejDoKPy7di0r4+Jl1ATbp11Yxu+mXzSstfhnwW/vmYq/t6/Iqf
QqxHFzfKl8CM1mQYZytE9E0qzgboYrl8p63MgwWHKrAltX1HM13FUoJ9rlTem58yMiebzNvprFmg
qxKUTHnJ/RzcPP6YUNzYw3XsDdZTvZP6u0yX7HMN03gOENZM5r20dTFlqNXftfq+JM0hNrOu75Aw
6ETkDNygPQRrMnekU1Ruj7Sv2L6occrYtQLSBlqqJsS8bPNGUxrH5LwPNL9DCA1638oGCdgyrIxM
XCa7HeCVRRMWbWo1nGhNssygDncJT/cUboNwQbqkwqNII6/foLCwYK0Y6ahOc6xdv8sc7M5YrjI/
0ivaTtsscF/IpIvhxCbi7ZrsXcZmZX9YdDXFXJDJ3+xbI4KRr3GuCnYf3QeC0DuIO22GCpHxwGzz
ojQf5pRO7GMAI8wtnTD5MtTabH0xJPxZIo63vyKEO1h4NCrJebGBxMh6DHXiez54dCTxEaShOe3V
Y/0dX3PheHHlUujPTAO+je3QcLhMgxkADhpC4jqR/zG+DpQWXVd/ELFU9wtO8ilyL68O1WuIcfmq
r9nX7uzekCuOWac9xzK/41GQkEXacYVuupuzdllioR6gAG/dkZj27EBlfYistj3ogjx8iSiXz8Xh
dsw7E3TX6lBqrRHKqkvTI4zPTEKbM6kwhfqFaU1hpElyfnBzhe+oJAt7sqP97cmyyAc6xFUIb8q4
07OIW1EMGbH/OOLnzxcuFnUjQ/+5e243zXtOyErE8EwV4vs2cYj4OBQX/n6pjln70UDttZQkJpOi
6CL+kCfebB86aOGwZZm1ec4FyeLnHSdy6QtbmYnL4FE2HJslz00sfTjyQPg86SPt2L9J/MZmb/vz
2qjcqOZBykZoEtcGOl2LhqD9zWNax+clHH7iNehsZWs/T5CvKdb35EqcqMUM5PI9Ef3noADvixlR
0EoAAwejSyiRZT7yxIUoNl1VEIasOQGsDbWd8KyvtTutwT6AWHQsSFYQDfBdXsHBNGbykz3xXbX4
83lrn08gmwNO5JnynRJTiq6CpU6RubycG5oPxCjKVaEXjfFCBqPx0CeAhqA8qKQKn+ene15R20FO
KjL7Aqlk9jfeN3CRHR94ibvKLdZShp1zrM7V78kVpqWWxg2vrLwsyZTIeEzgZpexp+7Mdu/7G4cj
1fP2knEf2lXNpFQ/Nl1BuT/VHqGtCxpGlxN2m+8MzDumMhpCwA5C534nNfy+SXB3crenQxzL6KZq
QPI0aB3gn7N1kdnFSFdwGz8fDzKiGCmS97/412YDLUF6CeqOBqTiU57OFSzgkb95ohHi8Po/wObw
cHMqobEK0pbSwfkF1MElXi+CuIGUC82BaargyXrwo82nTN+Ntxz3UYWqDpwwD5WLnvghLOC/cQiG
cN3i7311GJgwoX5a1Eoc7s8tvGVXIrBmg1xP6M5NPlIG2rBvN3S+dsYfuzB8lruOP2KFXucrgy6e
c3PtLJk6vahN69bxKTCczqH9oqww+YvwNItPzvEat16tt0Nw0DZK+CTN2txwiUcSZ2JKVQHbaUIY
s5arAElcS15vZajrilCQANFwUoQ13act+XUkBFy3B8b8JcPNBiz1dSuWddWNpE1IssoUEha3ZtuH
s8lhtdg6jhwdRzhxhxqQPlPFa9GF96b7Ha0fFgoRCaLC33lG1MoWVN/ECwGKVm3HgAOhESxgoe0p
MJcmdTWmYmEm2ut41WbMGtZ58o1IbkK9kuao1UIX8euRF3AW67CZiIJyAyluS1CV8eXyFSxNStzg
B/sbrgw0Hr1r4/kFFDVdZGQGs91J8Hokjo8rXsVMDuERewGSHZ9Lf6aj1HWdRhra1Erygv738w5X
6aeMV0OtSXIPMd7TKDIz5MLjycMMSM2rkvJ4WoZ9MSs7ymCzMDXq+kk7Fnq/RErlWK8q3azXEXg3
311vNF9TZNRZoqVP4v5QNS//V/bgybAVmqHsCWVQpXMTSjggQ50rJf/rME2ugj7xHrMLXX+lCCsX
Qzsw27wR1rhqYjMzv+jtBAyp6xCD8NrRLJSw//d+sLZaJAotQBubCyanFi4u5m7O+mMgcPwJJKRh
rf7JH5ZxLL2xeq27XEo1pp53OhjZNNJC5dxO+Ar463XKbsiwBixAgLler7cD7RpkWTHDYpRgacVj
z2HyvMrzkWkrnMtZYW8MRw3hfbKvAfLEvtATr57ibxvjXdzf4qcLiZtpolU0JorJpTG0huV6qAPQ
R1GkaTVBNSF21IOj2jD0gIrwWpw2XOjnuCXhnAfJ7bOwLDcIh6cgdjR+mnZm4/xXBXr84ndiN+Nb
FZm0puaiqGsPQWixLfAd1IEYUxMxmOrSww9KSy3waBCgbPcHevEEStaNxbQyKI8XKygX7SkPQa4z
z9SiQleFOOIZsOmnWHldA2A8d58LDjXQAW6MLy9BMQu7TnfvE+5oAKE7QD0S9MmRF6Dwx+zgbIuZ
nKzTvc9pFHohLgN99pAjO3pvuDFRu38vIxSdAaHjXLHCNYtAsThrb9CqgwNo65NYfEn2iQQx91AZ
OJ28kExRkIQVlEQJ9ugwzXNKbvBG517i9O8xUj6wF9LaX13Q0muzBauRNjmNNoplbmDvuY88RVb/
cTArSWW8dj1nFK8N/Umgdki2FJnWvIwHH5Ud/TEXa+lYssuJLbACKFPrG2YGKFVYY4bXTzH7ZOxv
FJjgXYvFk0X2ek8IQ3A/3U5qDm3kIPZ/6rYcQGCEHULVn3m56BoJqXBgqKm4tvueU4bvyR04FQ3p
5qkAbZP0z1bNnUwM+4MtBScqub4RJeiSQqMi6sXg9Fxss54NBEh7KWV4zO9rnxb+q8AN1QkczqfD
ilNwEPSC70NxKxv4rZ/7r0AmmhDFdVLbqs2ixFR2QdK3msvpLpRTRp3900Au+qw+3QGuZ500nH9B
cp6buuSFSBB1WYvIlYGH0tX8CZ7l0obeXVdrpdAgHC2qhV+9y8zca+1gh9A+wlWd7CzbDgtP/ubL
UhPyYFr8f404VWj/3kY/aggLOFHuKU0Q6NNMk0aoA83Oltb5KS12m/qQgC5yO8q8zq5zD8tCfVHr
KKd9wI0w50/v76x8C3QVswFe8fMoJYY7luDPXCIOoOROwSrnX+uBIFqDvPi7ywMl+WlTsANiuXBh
pCM4qUWGhrmGsY7xoni8VSvUQ4dTQaQ8kxlSwU3dSYIXeCcZ1IVLsfWqKicixmuhhPVfBy0fs5fX
sH/2+I9Lnf2sFYOcn/rKggsN6RrshR0g807iRxo80l+Nn4GF46OOjAhfS9vSW0I9VX8T5zYbd1Iu
rEa1UFbt39wBQogL69YkL+RiPi9WfdaaZehRq6rld8PlnwhIY1/YQ5KIH9u6PjFkbwfh8L+xPS7d
MRVcrtYs3MNV3FDKFJ+iSab/YMLN7SznkqHfLFt/DTy5IeGwrs8PMcod5lDUqKFaYzuQw4L9qIzu
uaiOc+A/VKv0CL54xqdyyltqBiJMpoy7hE+H61yiwxgm3SEOqajaoMMMltyiQZnl9rENRY67QnHb
dB54nHWrF563xYEDDPdG+jct9mcOMEOtdIZ1YVSAkZ/Xbsby7vRIflGYeQGbw9aV8+MiXqJHQFx5
D6V/pxdfkaGR9PqaXh2y9iSfQVY3DF9GD4FjzNFKzVki3WCvSCo2pA+6f7dlkQdFjlNTn3W7yAgA
omndB36YGq7hoEuJoYpRRdXREjGMHbrix7j805/b6PFcXjNRoOAWyuTfxU6UdrvEfVAlthzGjVum
BwxaUFZMJqNy2ffP0WK/DitNSP+7/BTSOum8OcxWu9NPJV6fNOMdyZyQVF4M9u0pwyzZiARfUJ57
IdsgEzndDwL1eug+5v2E7nN0ex0UQi4c9ulXyZkH3kTdaFlDKKgH1rgRai94ARW/XHKWHOYdLVlG
mVyZW0h80xbFYVA08AJ7P4g2J5FRXG6EZJE+OXAGY1I39qhLNlztPY9RzGKYjQt5wRUDH2raiE47
XzTM3Ci01H7GXf0tAbZ4HtqLKoWp3lVxJWw4i4rQnw+4EDBV5TkJYptwm5CTtdXNuylXUBKOSEoh
zMYGmBZ2Wh02R7oeVxUXQUYxo/ArSjvuOge6ttww5DCpg2oxvmJ36jZTqY2JBA4yCI3LtxdxtNED
ChLOXu6oOk0gGIUDuUsrpsKUr1+U4vM4x0tYbSuX2MBUVz5A9Xrs3XT15V5KAj1eEgvPUs/X6WU3
GaCljkryVfPW0xhwbd5QIa5xU96Z+wgD8BoYzA4aomllXxQLssGSMy9vRaTeERZgRZjK7P/q1N7S
xlbgvM8plTSgRNtHhy67pqoOT4o6xQRRh6xslxmoGDeaYRaTSstmRvCAwS1A37qgXmhff+viql0f
jjBWDPuAT8SHdMSZD09Mu9jdg6MzGihXnk6iTd12IOHrqnPQMVx5jooL4vaMGKq3oTVqhOlHQVlj
jh+tTTGRcJSD976LlsBg9Xdc9b6JNgqb/CHiKYM5aK1R73cQBJpIGcc6sTeVjjQPqCZd69EcOrO7
wswgSlA+qyxalkn9jkuge/Oc7RGPAjEUHNfrl27YXCAzTlovbkHT313x5ERE6nCGMiJpPZti2EK7
F9dChYrSbV8Wn5ELu78AySC1CWff8oZhQYWPYGs26xiVv023AmPFWjSav75dWFs4/wAStBW0LaCM
o3XV46q5l1g0DWDVASjXG+KIfjqMV/qag+DG4xKyFjx29W518cqk6QiERtKdncVpvscUdq2igDWw
50An5KlsJx51+SOr/14jAx05MFyxS1SmcgtPOTLttUnJizOpmmYIebdgnEYf7/XM4mZdLRKG5Ky1
RY41H/xqfbrcYuVcG0vRhJJtBxIhlScbJjKjNrdcQpmQJjYWkPccaD/wsWHH+X6K5b4HS4SUFG2Y
Q3prvnUEk+cvOHNhIVsZwMdxGa5Dg/ZYlXJjoKQbhvW2DO6hVCaJDbxYU+MeKEwbDn3/xMMqP8yU
zgz9YGxPclUT+w3tlvZb5TapYRJu7LpYFp8yf4g8Ztt6d2lLywMMZ0K/Ydv29Bpx5qVqFPL5m4Ji
1re8cabuSHCJPODaD3Y5yy4Vyi3MdeVyD3ZhL0e6NoOHWSuThsG/WrJs+YlZMEQol3uhfD6e5FoH
xFryvvnoHey5i6n3UN92Dr4b3SDaAU/y0PkA7UXPu0TdP+Wg92iwPXM03IoyuC4UiOV5D/jyoTXk
Swn57bUlPBeCtl7sLLhYAn9Wy4ss4bIaVFpY7o67Q17Z6CkID7znIM0r0HnjuA4NulQ218x1HG59
RoHJ3h+OrJuhKZUUcmggLCVUdgeEuKguGiDddZWToSQYKBDBWDdPFI446hF98ZPl4QgaJOTzFtDS
Zr1rHi6eHoke5DoS/MYXKvKMqbt6lokxBrtGXD1OQF6D678XhAfVLTnTT/8ejXpb+PKY3WLfDXZ/
NrInw85STG6ucJxkRUbOd3LYjdZ90jUmgOr/daECtXVVHevCvyxII4h8j3pLSQ0dF29UD5L2Q7Y5
CpSgkEoIBUJV/+3dwrhyZvjr+n/f2m5ApUA5TW5dvEwRQGwtJpTwDtgCY8LNyxLItSevprU9YuGk
nbllDR7gGkV4kwPfBhBDeq3NW0SakPYjpZfaTi8eCYBj30sXPdda+LMNZC10v+jD9medZoQxJBhx
BqnEFyKp60en85PAS8SSl5NzNtvBlEjdS9Gr9hqbbjC617vOFHTy5GfZufRK1barhWDFc6Bq0jnf
7JA2+aCKA0pHEFyqCHP7UfZl62p2gw1rIH4M8MnQyT3CSADCmcF3ynBPYpx5rrfv6a8yK4w5mA+W
QonIX6LjK5N05KyRWxxAqUA7UuRdIjTBV360WUCHVo83X1UN9jkxYyC/2IsJFb17pWwwbUSKQa7P
AMguzTTFJkoQi3h3Xk4QQANzdpSPZ/HNp227ErdeOVy5FYb734989E0StyEOMNKtEuSlP0zyvwNl
v/D3KHROW7KOpd5YvWU4Km4o8ZpvZqOD2uoqIYOxrMTKNojc2mLgdmsTABI7EKykIOuZMPl1CkUn
m2J5pmy7YCRI0OZjIL8dLDfq5Ory1lT4mnaRPesu4beO7/rWUytwsx+u1EBuxq+E3lufBsUyClIE
1SJBf3fXYq8oKjK1QGf6hFyvkrJduTsRwpyCjV3zqcgtvaUjrWNx/+x90Ny5igugMYqCP6QAxvfB
eY/hgZLwGQdlk0t7VulBKRhGAebdEeImKN3jMg++cG8XvBXENHJkaTZ3Ban0Xs79cppsZtxHJxn7
f9B8qpaX+3G7V5Pc2Tl1iaDa0vYmPZTfVvaGtG6a2wSLJMNa4IohNv0eK1vVj8CRYvfadyYlJr7H
cCBOvDc9USv61l058VQZCmlibNFebepk4394+XqMTXwKk4mrNILtgeZIvh4ak3HnmWJIvS3QjWhh
76ilbJJzGt+8zWNkTytWMel1VJK6ptAsetyo+PXF8bEVYKjQsTD7t06DuRNd/6nPqezRYfzuboQu
02TazUkn6kPs14wE5T9rpAZC3Rzbtj6XdHUhMRSw9ZW9t50sX9mlXpxoUCbDzQbk3/hqEPcxcoGV
wBmhiEsdQwgpxHwtuQDiS9dEqbSXSnOXFyLBInaqSNqSEtCi2gn2KAQ5IZGDkGB8IE7yJFzqOjY2
fYfb1tbYa167J1CXB4Q7LjkfyVXoG5HIeLTjyPE1D3nJpJjwtUsE1VuoYa2Bzo9v3YHrAHvPPTJN
exvW5RgwnomL0tpCINbKmAylrASipysY8MRRhQjNOKh9SMOYge/II62GoRffxl2FVIX3WtaUqFhz
23a3OqdGha8F00Q/eHRThzaqN0GpNGqfmMJD7slMUCQRHainCa/dwHoEJ+zQ8UndPBUTa4LAufoq
hanRBX3DMaoB7xBjRsfN5mCUEllOzP1hgQgF9BWWeK7aUfzpLK1CJD9MvLg7FIF8qpPFtmd0AXXZ
RTwFPE5YCB9Fo2O9OPFhb9VvmMhfQ3wxplrNdD4jlOWLKVAl3Rcv5u01Ujw8LMyJMMsnjtetHGRX
PFeygSkW7NlKKUvR0UvOPQZocRKBy0gHedQHa7dVKyW/9/e3NnQZppzYsW7oVRBoZxl71o4h2xEi
9wqLsoMKQsZqbmf+H7yUw3qwmAZ07HoTUPR2bS4V8c0NoU+nGq3FXRr7g9qHexuRgJ2M/azSTuqe
CqDu8i0JNphYibQbEgcUu0lug70qlcA7qjsyzZzivfNOJ4viRW0JNaIhcCiBCFngm+i54iL3zMQ6
FNkC1WJ4C2gYOqIHCJfJVh4l15+Z1UxsbzZ+3jAZheampU80yiukDJU2d+3TWGeL0sby3tO12tvO
/W8lzC9OUAW2ufXlQbOGGE5RuuG6JJxZsTsdjAvMdhOImDH/cHjv3pbKtA90FuL6AuAyXRk/dLv2
ztVtrpgIv+nc97gYiLu5k4TbsVbEd0s+x7PjzCZavnRIUViEgSuPZMst5/B44PoHUumVGrofAv0S
yNvG4IJARVREk0lp1JWLFHS0NtWDtBjFK/LFvH0gN8t773SCJ5NjbbsejDfH0nDBD/1AdWcale66
uMYZ1rzsABt0eTtRyAnkWlAC2HuHVr1PD2w5c2y14mwTPgX1Yq3Qn78ggB2fvwiJXEb/AgeO2lYD
5zkYzQTQz7OQmimQVto7J5RHjpERM+4tTElD/ZVT5zbc8jPEI7jvwmJKes9JHz2k0oAsabfZ3Doj
0bUMUxYPbgp7u+EI/3qu2rz7YiFfhdwYB/kONn7eWRQtGRRlgWjxJi4qSAfjMjxoF0BsaOCLKGtT
Qx5NS8qSCHBMnvSckUpI57Z+EORKvSBNc7yjea9NsMPMr9zR9cgM2FYVfR+4YKoDh2l8K8eOLBUQ
SmZTZCXMQXnBGw55vb+1XoQxscb9PxSstyyblKHrTVNVCfW6Z4khIBM/XEjgA7OjSSPcXwKR0mQ8
AJpgb6bI+nD76ge6BiiKN2A2gY3W15RWjw32oLFKgQZBkXHAcSHKFkKrJ4us71xJV8ARnxHAZ+Kl
nyWO7mmXhh0qE85efAieDNd8n80kFqSKipjLsDwcO47tiYQAgrI5hBfNrcHwFHLYVf2w6jvbDN0Y
8x59e3PQE6dbW8HXaAxck73wqRYOlUKP34mw+N56kBMfYauiFBbdIH1DL1n8VnKXvrq9SGRMVjwb
Y+NmjbkLBp74r6sErIXbif483mfvuMIXPT1cbH/h9czkSXgnmyDtF4AleS3XYIesdJVzKsRF5Zwk
ahnJS+N9DZeEYXiI8I0CdtmSsMuDFdC3/4lGCO6Y0msH2JtF/LMW8YH9gO/aImhT8ISI9s8MLVXQ
50QgHeC+WyurkJC1EeW2iRguproHJ+pwSz52q/waEzNlBOhtP9SM8jAyhhhwh8hdv/GKfmIp3bO+
QyMNOBl6dtBUsVpcG8LGgNbcsi9zm4wjkaXxjq8N2sfVKdzKI+kSFpzSDxKpnZqOir406cJT0wdv
ZfsFIgt/1M6jNAH3yCEUfe722iACwZ9hE9dtbC9VNkwWprakit6EwpGL0dK+Ut5io6qzm8b2hmGp
npGZKlwx5GExRTWp8sUPUrBpSNnyNa3+Mi73JATxxE5OGWDxtifiBSqrJkAkWk74t5CoxoYPfW7y
IM8kduS7OzSbNoE9LZoPFASN7jQPMxHq7lS7pb7h4iSDR1cqNiXExTyBoWiXfDWS2JqHsRO6pvJn
BlOno4sRLHaxUgP/ADO7lUX4he4UWKyFhLh92ws7mUNhLPFZFVSypXa7rMtxFM9sF2M3qV967koF
g/9vWd5m5XovbH5EpkfTIkruMuWZB1uRi3X4bsOPljEf2qcl7S2nRcIVuqygDgY9g+PvRILS1Fa2
ckI3w+zZH1TKjPJ2i9ThDr7jTURD/yW7k7A08jcrfyH4dUwIyD5+kWt2+a9B18wwcbESkq/Gqx4d
GjLdxXbdfwMp4JCxZvz0GESb30vF+Zye8nH6RWdYm+jfptBMEKqs3SXgFqxX3ri9LpwUGAUP4DxX
zKDaiabcKuE9wO1b/Ph0mTmhCYrC2iX1LKoHk9BEYjHtZGbb8aMYzeLkaihh56jn3FNupiwX8/d9
1wbEXdbtwiQ3ajMm9gvmcCkT/WMnwuJodS6RBfLBGCKQ9JKaw0NcaNv619pCWvekBv92A14yDCgq
86C+8fvAv0fy2dfXAfRhyrGZJarznxkkVZz4rpMtMkh3tUb+zqZUBm9SvA9IyApkaU8lUubn6zWH
hvbpUzYERh1h9gKS7LvDQb5uqWAazq7r6AGuGZSqdFlQpbGcp5MJLEyCPqt9twABSfMyv4TcoOgC
+PeOpRbf8HnL1lu7YXhn5p2YId3939zGx7Gy6e5ATydguVl8ALTBQqUJYYLTyM8vbY2US4hU15Q8
UzHTaOubENTn+FFZiNCw9hEz/sHwwCv99OfvXpvLKEbpDkzO0J4XTAxedhGV77uEOSKXEh5pZcjZ
pvWxSNFKfWEvECwONomzyaJNTT4rdATnUBBPZWEncFf/N4OPrtzgB8Y2pDF6jjgD2KRofXJ/2DUx
r87jhCJOrl7plYgyIAVGCFzWlQ7kbfwQCxIVocEZ025Ew6qxsMOQorvlF7A2enKKoBxIRYVR5mg4
Y7ZDUdysJFbmIglgV5p9rdj1IwR5H/U3NzLnHhpFc44yRhgbbZV5gbuRvKWfQOq4yEVrzOMlWcww
dBM16sJsAsfVe6V2YXHDCrb9FlTLKPU23l83v4KYHZnPUM4ljsHQRtHoXelJIV7QKLjCvxM97lJS
3Ry/QseNbfFeBH6vOZQdzvPEL4A66XLnfgph5vSDxIDHGHBKdyWk0QA75n7D/re2bmg1Ftz5zud3
AgQ6NrJkMOQggyJsck8sgjDN0Fu29FmtuNmX+fcmmIH2rwBIc9mpjO+MN+y17W36hrp4rE+1yMFR
c5VQoXeoRg9R51lKM5/+FAzWlozJb9nqOei5JPJMDleEVla6Q9Org99wltT5u3jqMczKr1yx/JSF
K9lMy29XLIyJF98Ls0R1xKtn02euglzgHBwNphkuW8fCoAZ4yLRCYUKKogLpgAvWCvQ4uBNsk2JF
w8J/dWl3aHbDB57L7WV9O2XRX90MgoD1tYKa5rNROeU0DwYJbMS70uRNJQqZu8HL0TSap/cud2p1
HzMkGzwr2rYvi463ZniAsGqIXX9jiOriaaSo2B4rzFVmLm5PjYD9BRW8XcsrKG0KxknPXO2PkdHW
Gvb+B/q3SfJODjODuijESbhpeqfDce1Z/Xb/Nb4cHU9Tjbv3wdjUS2ifxJ6UzT1lyg+GBztNYFX2
nd+jsH4lu2dDChJDqHA+iqZCc7Ow6HevMQZ2QUMbjqUWiVbiirZ4IGH2y6epaFSywFvIGJ9SIyov
CSDdB9NxHolW9TlVZzRZuKmPq8suBdVMHUA1uyMaNex7cTlTZTOERmjUYY/vHQT1gytxnyKUuKl/
kZ94AqiCQzKtBRcd1edjZ9afpGS3sQ4FsEpIlpODFxIrGJ6nl3yJosRVwDZxNuHGP85RxM/8zquc
dFdWPDAhIxxETPAmdkpXCrX2zszSw96fmR/M0/g16DtFePXzmWIChkWq0hMUv7Wv+PP69kEzd4lR
hQFK5LIn3X5LtneFP01GNFaj8GV3SLtdsqHv8V3AfYmRjDiHzVyafeGtZ7wE7gvd/aW+3qWe1GLk
nKCO2/0GvJoJQWDe2qe83F2AfHLhyQ3nSe7h+5d9Ue3itxo3CxxWqd3W8XaRn16Q4BNGdtlf3BxO
wtfSyuewT/AEghr9Dlq/+bdb57zSM41rnYAkUciRDvZm7nh0O0vHc74vkcmInpWtTe+ZC+VGk7aD
inISGVeai5u8ecH+UXta1Mm8+ibnGWVwAPN3jIN8qjdk6uZuO1EITDBTSJoPxsikMOmC6Zpm4CjE
9PKwu5dGEXmKX95abIQt2tsjqxYklyeTcA0kFFnaM8WcmCqfSGbPZNfeddBs4FlLtPrhz6kj0gTO
pUJjvOtg6DoeTyTjcu67prj35mEcDvVjk4JAMmb6bgyczcQIbbh+ZcJqqL1sLfyuOaX2nsh9Uhwe
E0CoRpH1fCC7i4weHghzdDjwLnQt6pKrOenu5a7SLVctP6R9cnMWlCDFkIjN1Coj3oE/eGFYGS5H
cTV8tMY9IKLK0C6f0Q0OpgkwCX4rYy7KVIGCfV+fj5TxQt0EVtcIXUcNrMtU30Xd0t+cmI2y5Ix6
EzJ6K1P3/eJwqFu78EKtBRdHjxPH+f9XLSkuJSdXDW4OEjcRivODQ3DgzjjyVFFB46UnmVdP3bgQ
oh7LieR6+pTxWpyWCY1M+xeJgnWJi2V7Jq/ivCbH6FzD+FrJjR7+RWhxC+NG188RW/l/nC4xIBHo
EB4a43vUcyQARaPTjNphR+jZpVDj5W7SA+xOfcs4022zL9gA1JjZkRlmvEknjh4JB+oheQPCU2HD
nolg3Pv/C0K0nTv+IrJ6NTv9TUSuqUYnmxqWbXDZPqv8mMbBoNsgqVtM5PCstiFeiMzx3R5DY7yN
4NmcEQb5TLmiIxNdPqgCKMQQ0EBM4lzW/WmSV5hy0jG5qab3wV5vYA6CrgtVE7mWc+qSzWtkRiYy
Zwz0ZB5DXeZkBCTL2xY41umWe4x7g2L2TeFfsKl4gYuOY+o/uLDWjg5f4DfHR9jMd481q8iLqaXC
IK9CRViZj+QJXgP3ERmpcEzJ93ufZjoV7MwdnT7YjoQYWJtMH8q8sxvm6CARQn33H6wXpEt/+R2p
oM1s1ykOPC9yG61ZZXTG/FiEL0Pef6Dl0/38SNIU61iwhhjDMwNUvxN6lTqGC4/3DTvE4GUjcQmB
i6W9jPPfeSLVSQRbWJH7OfuCIYKBI7f532PxM09MnPp9ovjO2/FNiPdc5FEZseuVGxSCCWtmz84l
Xb4ZtfPLqyEM5p29LZ6G1HDpEb0KiXmr7bxEuNG4lazPSuLT6a7zduNbGrzoiw20gjvuBMz0Gdkj
k/25hkJ+2lVPJ4MQ9v8QX6N06RZ3CFkiRAIcDOeAQ6am7lIoeX5lIB14+vf6URZQDOT/CLh681fh
8u0z/QHSXsGsAvnZc7JxBjkVypgR0/KqnA83eotI+/zKYCrTfe06FG81YDeltkuvlBN820UxtCWr
7N/wUJGXVsD+iaWv5cr05HYx/6nLiUgImZfd+llihXyjpBP6/FjtJBsK/YIjaoxG89jY0HAlSCgA
VUgI4i/1hYhL/eOfPhfGc/10b3KeG4ms23c2/yyIPH0a5SOBjLMMV+BWgBcIUoOPCajyHwPPm7BW
Qzt6Bpq1vCyQY/2x7EObxVfiWindnRcw2HWZT2vNwDN63FZmtRS/zhWIfrKhi+UltTmJeYzKfjQF
c37expd2yRnxETddW9Up9OrvPE4OdrZnAeP1JoIadrhJay71xPiBQ2SUI8c2GBQFrEIfjYDi6tMU
KOUmCVnBWeP8oqvmFWnA+KtjoQSBpL2aN1eEPBTOcgWlih0W3MRm3pLV3VHmp4PD10deANAyu1pu
MGNDP1lBeBNT+0pT5RkqIz5GpEyQSrJ51f7HFk0bUh3pGH5f0PljMrYMm8byVjEoPnw66gKvPRr7
VHHFnwaVy1bmrYqlZf5vbM0TZvdbtvi/OL74Z+Z/lGfS8ihaWvpDggBExVDTBoC1RFjzGMH4jJl2
osRNlQr9pkK+itb7eTEsdaKpfTA137pW2+xcUimgxb/hJNuMluB6GtDuGlyGD0Q+5gEvIq29J2Wq
vZlWT94nEZ6bjf3HKTg58/DB0melLc8fFlVWKkXS9GLBchaiAi87F9OJhPajRbq9h4O9DRq88Mgx
6d3sjNMjSOaSE7ZSgfSoWnKVIPlKxgE6XE3rLEi7uaKxHTjXQjyLUS/aWIE/jol6gwhN6GKceaRz
9g/S9jwqG7fzHdUjR+D94SL7+LJBok73tPJoUCM60XCDZ0tLdOxE3IgaURSNf3Z8h58Yi3rQP3sH
WVmZX/aHqPJewC1gbD5khuH9DfOr7+FDirRVas3C5oTa21ThLZJ1zZ0SHqD8Cmnn1KXuQDl+I4vB
4uzTOB0MSAt+wZucXsZZWTzGFC35boPBsV21FMq+to4RB4+0w/5yRAPvEpCj+/2wkkLQ3/hldmPd
xmQwg1CXGlfGnOd7GI93MwA0EshXRDBx5oWprK5KWmqGjeQm87qvuWkw6p7kOwI9gJ5eWUU55tPX
izqQ7WYy9IZ8ObJ0ZlHlbp0ZAlUwKd8/aB4CnCSXyVCpmRM2gVCy+9UB9oc8BELtNEEaHZ/SCr6d
bRdb2V+qlbk12NNhy0YbF9FtPZ9EHtamYj1r+hl/n5dku4RlqyRAZCD61pJxPYhzvkfnLaiXh+rW
K63XFwRlpj/SkM+jhLPQquEmOAZ50cjQhYZC8XdbNoTlQ7lcdLed9DljPfUGcaX5sb9239sp0tvv
bQlIqxDagB8xUoDHch8TTU6cthjEu6tSI5Ne7W/9DsAyOeMFnQum4EB0xSxzMIrJ0m+qqRdc8huG
F3RLo7ciVxpd0Zpz8464bJ5bFAUHDaBwwhbxAH+IwGIGs62CKctLq+p5BHrpvmdHbqe6JVYRA9/n
RaFapVZ3Zm/Rbazv1DlPnRyNZZIut63yJUZtGjL9MeuOB+181FIzY9u+hWDCLCKuD1CRo9wUirn4
lu4N7w+omfEsPUyLsWkROWPiYc9iAOXF70O6x4j7E12CYkt/OXzgYM3DFqaEs08OH03+FFu8qAd/
VRH9i85PaUMI2bnEHSARbW2Q1yzKzEqLeyVcSLqIXeoFSbYM4DTp2h2Njg3dgg502tcAKBQdRZuH
4BPF5ttfZlsCJm4mYRVu67xyhkSfvujXlsLiLPiDBQ/fHMcCbIGOS6ry0kk4jRK8+TNxZ3uVg+i4
2mIT02GE/HgDWLjVYr49oTVwypfyQaRXYjbRn9Q4VTew7cN031/ZxaQi08POIw9RtqrPYVi4P8qi
5LpWymrIn7qHkYv0K6+XkVM2PS2dkmtAvVnJwkt1Gnqb9UFjpHKzDWUVZLjx02LP+nCu3Oedac/9
hcGlNqasehkThBvCt6AQEvLfa/YwKRPxMKgLiWzprOA+HnAWoFPlfC79/Ku/dKtwPYaKWgyg4Fk/
RBOlugZh7F+GY7CKfHmOuuk9wOE8N0Qi/MFMTjxqYBrdEc9+avbjzgftc8dJFjpoRGozzOrQCkrO
tP1o2NErbxk3xlrZvXqQDMs8uXSOdtbjkkdmRCLW4JdqQeLP+smB4y9NYU/okrm8mBGUu8nF1b/G
l1PHz+7mKI3L9q195FwKdFLgrdEUhkBvKgUKE1LICsefkseUqWsLxWX54eXGtrZzqW7YhD5jJaO/
E2ixuy/xxLFIV4zsIhUdm13ITqkxSTFelA9depuaZtDO/qKybH9bToWePwcvt95YSr2bOtLEYgEx
dnOrBav922YcoWUgppeba5uoeXmwr2Y6+ExjG0wUZgmudEsS7QTFcIXw6w+rrZ4NJJMwjgFoo375
F3yA5VRYjpEg+bi2RgJaHLAghK7J4CNtU3tati/wYCMKGZKR0QRLuEXHE4haUF+r9pLA1xD8MEgI
OZODxpF8oIYaMWiiSE9RZcDtwNj0/2kXZ5uPVDa9N1cD4Xm5sAb4kBHS4MauLpiQm37tFAI9Yprd
tPxeKKMqbbdUmaYKH2brRnFPGSDmfvO3M0ZLaNjInXvyZvkk7HSuytGcklEunJgGydPXzw38E209
azjXigE9rR0pgqVU84nxCv1OOJav3No5hUFWm95zluX6QVkPVrBxeGt6yINCT43FC1cuDahvBIrz
JIs1xPuwaWX7P1oI3ebAebqpqGXtYZ1fGMQbzj+eM83Lm+C8gzy3zOtT0rbLpwM9DCGv5UZJ2/d7
OxZYNY38qg7/IMtj0LM0fjw3mGl4dS8olo/BJuDJ+soRkDeS8FKp+PMC3/HZR9CiX2jbinrxytt5
64cUuh4nPaZIRDNw46kjD9aYTBXauVq3qzDHRxER7Uee5p/XdEr2ngWyV/H0Coy4451Z0urXy5if
Q8MzXpZ7OfLFmEzZ6BnQOTUspL0LAAVT6rYDvg/OG2L4lAUQBe04sC3Z9RmMOJEyGWHvCdpTYvkh
j4zD+ndKaRBHS9PQCup+vNZUUqXokD4oZQNOLKaSgxyv+z+QviU0X90/tr1Go5Ti+BlNWyYvjoat
Dk2l52qF/XOyJszKEM0ilifluOBcXCY0yYpYOurdZYkQBrAgj6XQxaH9sKZLkXIpqjsgz1bEpyRv
H5GmVqAGZgraoqUELLQ2lqt1Zi8oKjmQHzioc3P8ygUnG22h/I2eXLeMjBrmi74dr5QClEUoFadW
CbphQt9glDVtQb1XW/a1qddF8jCiztmssl1YjUPmEbCo4zfRoertyoFIgrCRDussskTRKS1SWI6q
h8xtXf1bVrW49cE4cljedCEOPocxqKCb7U6+wfvNR5Nu0NzOSIdpyS359pC9p7SENkg6noW1IFeH
L9z5YJvRB2YkZkcZySY3EMq1pRIBIpjkz7SWBfMoh2EnrmwhjT59TtGiOFMQNlaXSr7AutHalxsT
DIRoAqNRPBYUgNawrU3x+0N7N/0EnCqjhtOeewGI1Q8eKzBfq+OcY7rfgfFYb68NN4Lf19tUMO0F
/AQ0Z5l3l7ufQukN7C+5J41mTrbaSa5qX/nwyDspNMpy1dZEDPNd1tdkIoTMch1075Eprrqw6/QY
nMxU06DckSEUVVAx4CUR1awICIeNJt+ff0Mjdjdzu3Fl/I4dCvLPysuRUXUM0X1/RIgo9fhpdzrJ
vTJHiO3gDPRuRwwD6KWMIkUW6eW72CiYTy+CAm4EXsG+OmYQiaI4VDVItg+d/qJE5D0Tpks5oh/9
7HM3Na+7mK6XYq4JJj1NKd12JLm2WTqjJQ++YuRcE7uC3fbcsaQFeHhkqD9gToDwm4we9bzpnVrb
8ya5X8tC9oDct5VyDIlBEM2qIe/FZ72dyEmkU3hHug7S0ZyTWgK0V522R/rtfYAhpuS2zX4QocF8
b7p8nFtcNIaxGPediiXmGgIprUIyb4TBt3R7oosCakeunPmTWJWig5iAW+C3gwaQZP1u+gZTtC33
MAHTGXSpsN8G/Q6wCpFWuhdrQGdLZHib113qARBuMFvzoI+KuQvQHUUn26R1fQZDaV42JoE87Fko
faoY7Py2c/QPQqIO1TFaTQw9Ak5vKUhxyr3oGpzjHThUUJtO5Ygvn/Ugb2UhiC01NiFut4FGrvIf
LcuDICc2QJtA/yciOlkC89O9hcgWerwKquRt6k8FrObuc0gjcfERCZhP5GUXHuj+00No2BIsUUce
JDGZbD8PPMXnmVbumnG87fqUisSYItccGqiQ2upPcy8AiT9FvC/jluYD6EynnhZYwal+xpD0up4u
JZwwviu+dbfKnZvshQaHKcTYox2KG/06U641zM7V1B8aEuh7pMUXlNpXyU1Wf6PvNh9YtT4oFmOw
mwKP01IDO9n6hqp171MwMVtH7mE7cTujLwLR5vMyIQ9hs0+K6IfSHcmFOZVnHO1qM76vsLH0JiUj
lfVEIUbCPJad9R5SwaHud4hACd8BB0tqVu0ajZKND0i4W+8cue8LebZpAs2lRllqPUHeOm7V3hSH
2HgFF9VQE2FKrR0vDKnwwzzKddHwSIg9l4uUTxXfj2jQVmyxi6A6TWhSNoE+hXstg/75G5lvpZNW
6wvSQQ4NLpTmWXP9bTET1+QB7yX202+RQdeNCZGZQsqvEcFhEby8s2xhT28ps9MfsIMtL2TlXc9L
GfrS5oF2dPpxQLzE6zNJwQlW4RlfIvodahpfmtMgsIvG8hsV5g9W8+1FS+FLdpAiFcAI7uznGW2y
nRp9N/8DSV07KXe40pI+A6yaS4trTsZENZmppmp7kDNB+44mSiRCf2mTVL8i7S47uFbJfNO7Tb0H
v6f8ch9TmjBzCzgFIvMd1lcZaq59/taiv2Ky8NPQ9XlHA0WUec4t3OkVL/meuURNXzxxOW9AV8Lp
yUV/IRKQw5jxptg19eXDRLuzpfj7hKtrlTKHGNKJRPZrYyeouH8ndQmNOH5l9LeyJohWq7XrGw8h
mKroN6x1Z/J9wNrFikQVLfJ7LrfHk6KkXE+4S5wpTMR9ZxsPzBLaNJWiQX+/7Ic02/FcoZJg3dDC
OhzbEO1AJgcDmOatE8spxrDrqlEedD4JS38PmYcyN4JBAtmOcqqCm0tVYYN+eUauHpzuBeXqXqUV
6tLPlGbzPI9M44XiiF2NAMchPTUNvdtU0xaOAk276LRgiuACnkFkyfXbbEU14zmdEPu47y6mdk5J
rnz9PlWSnH+IqtEfvVoX+RI4YWGAxNrOz6xR2rx/qiVZHK5PMAOB68wZxmWjBFqvox2LArC6Jeog
Qt/iYOZK4Qn5OxakntvsSxmFwsazrWlVqofU2JayX4sfD4p2ebyQqicmI8wPrm8goNOFJOjCep9S
YKRy4hW4+PyilXfW/yAdK2X3c3JOxrzVtzO1830kqySCOgvfdRnnLAufI3/+nl+d6nYFqicMWRWZ
hro+W/DZwMzc1xBvnFZPoxqSkJMjn7bpxs0bLB4axmBkOev2vRE34qn5uIRsxHcfJdTGqOG9UzE+
hNYuTHgKcEUiYOad9zB2d/uJUyA+S+TfjnQ0mlwBFrlvvp4ftCICLnl5rdzAn/3I/LZ/Uf9r17rR
/xCPB3udSYDD1+jVKJBbwye/G/g7sb6ocziZKftqme+A0brE9pkyINcLmYQmzvu9PhaV9tC7ZRG+
bLNwHWMQU4gP69ngjitN3sy4mAMh32xbXpn57jbBsyz8WzVpzFPq9SsIp9cpGV4dyL2TmTfZhqPz
1yhpPo4i6U8iFFFG3zue5rJvoZBhglyIP/jlovVFZb0yv0ZOgbaOoC+0pH1ixpTDqEU27Lw+2Ga6
4CP/RHVdhLptJ4m1V23eDJ6dT2JsCge3q0aX3bI5f+Kofh9b75cJccj7ub+Bsq0aPOY1MhDb4E7N
5PvvPNe+kfijcPkjwOQJGcJ8bJrP4eoDSOxSY3+Gi0YjaguT/yEtt2felyFQrTRGAMKZTdJx1124
z4hovUAzkOCTxsGjZ3pm7U/v1bWSKTyPPdlSQj759YBTp/K2SuPU4PrePh8fogpQGKCcv64TZ0Mv
4EFlUdliHBUvgMOkNMfZNtzlHKghpQhiOKcsdq3qftPngZyLA5yG0m8xWaUSZuZU55Sbmhw8S847
BGl41z7kTbMxLnIAaPJ91B/ImlHdT+eQcdHPeUlBxjTxjZqfcsdf/7+UVnA72aVnFi+8tYQmgTRN
fkgUNt4VgMXAyBcRYGU6p4pUy3pUE30fxZ6kmycTDF5i6KxH0SWl+iFbQQ5KiE7r/UrDWbDDs0AA
wzpYmzKbGR+a3zGqvNhdahsMgAPN++VBluydBwG9O8me6Sde4vX+PdA2e7wpEvwjSHiqGwA+jno3
o8yze5/0uOQpZh2eD5Z4Arjx5BACgM5u5TNsk2jzIdBH8MHoE+DxagUyhanvV4nkBP/5uBzDruhU
artOT2xbHhJphz1iDqumM4PJXELxZ8SUulRvlRqRIzLHaXncUgkkVcsqr5KzgzLdEWoiBZosIgvE
lxCZNcDodcn/T/dIRvwC6EaTpQv4J3lm2ESBnl2qROOwVrvT1ikfLSVcq7SnHrp4i4n9BkMok8MN
9kGLv2BbGwbtyNB/TnOrUCszna2s77omdZzeKVnTDmSD+RGDNmpQS117VnVB4cv5VgFHZk0963mf
3QLA0QxbkPRDaQLA6okOdbfwwZEi0Em8l2pe2Px5Q5aTOTtJT2qTnvIJdM6GYf9L3dYTfrK8pr6F
SguyPvcsRy/QYlNiBZRZBVfNK/90AVIdCb16zq3JavSM3Dc+tX2HOK2nnhy8guJX4EVUVww5lQqB
+yMowU07G2Fdej/66uzRLXi6LZy5+ffTlRIq62Yc5KlTuXE3qhVlE4juT68X/+u08QF8gcebdWyA
b1ydeaX9kYzHf5WL2iSdbO07UsjpGRp8Q1YduoHOUfqaFLKuemwJrINplr1yQlDAhsAgstDvGfqR
Qyeq6qsXv3kMPBoCub825CyqKgVT6ZfNcmgOwYez+BJTDI5fI1gQ7BpYKO3To36YHnv0Qto0NcUI
NeAprKC3CW5fRokPHDqU+mqGa8jXsYey8QZgJ6rLCDE8GB0cOhl0YaqvI0HZP8pOQ3b1N9xCmrUD
u6MuILnEGCO/O7Mxg3AJfX7LNPbrE+OlDREYLYuuoyHAsmSNW4JAh5k59R1UvW2xWXvyH46Zuw7w
GJWDu6mF7ZH1jarOVkQm2rmhiE0lr/toTv0uQIKEvv2OGYsX+5aYmsPAiIddTR9lTWb6oPUNsU8l
N9AOei2bsRJk1QpT1rK9vRMtEAKAmSkF9/KZ8KTppvakNbIpk04o91YANdecLgjW+FpzdCHLQrNI
IlZIs9DOtj7wfgvO6rlJS0XCzImKxZ/5XNX8kF1L0vglc/owP9RlK+3E7N1YtMHGHzYnvQ2hOw9p
kKucd/8H5z0MuSgH4/LGrMTtrwD3S04rZEVcoYP1zSn8dThi1zbxU+OswPtgT2lKDhkbAK4SDmf5
ucE4u/YkKPeIHcH9jma2FbTW4HrFv41eye/dSMNK7+uw709kBIsz1/7lWYrBqfmkspFDKXO9NVSR
2DxZD0ymr46ooZonimIkQsimcrMR9Nq7aSegJiT9f5Dvt+g29dG+SzYdJ4G28IZn5X8HLsoXYi+t
TjMwKEUUd5A2qaaWyRV6nif31P/+uW7nRhctKwGHtXUjPRHY35ghaFEQhRXiux60ZV5pAvwvIsUx
W0GEgO/W1RaEOVT6+FALC+GAsznpuYtSzrzQBkNs9ebR9lcJaat+LbzscYQlPdGa1haTiT8mLGDm
6EzfMgVHjJ0CXZ8nAeWuNhy5fgnwLOnzD4uU2rCvBkBkcXgyLWR9o/bIsJrqkE+DKvXVk1iaXyIr
vRA3nqEmg9fSi8sEwAiZswrWNKi+oSlSLdAn2E1aO4Ws37x7z3GB2vTzRx0mJ7NZV3MWJQLe5tIX
+pvyMX83HXQCJa4cjkZwnH6uLheePqCCH8vE/iWwCNY4lJabTRjWpBiKETEHnk5GY1eIMXmNliKB
oe0cBsaXt3H//X1uKens/vpmI8Es6rbar2kcqeW8zGd7MmfsdpLCPniDmM4M3L1nBPqRHeDD8XNq
WprgTOP62eLjFhv1B2bNRdJrXXcfge32OHkNZ+mZIFqP9b78RPRzGVmOgT8zQo6LtlCeCdGW3wvz
dHpHPtlZmURvltmJJ0w8n6as3KasF5IzY4UCu/qbIk5e023brXWsQTZChIjecxkdIhhlo40s4n3O
ofyunJ636T8SDTfW1Ix4r1jh6r/OAg216vlPlWMg4cqeUrwcdPLnbrBcH1BF06kgHUczJibHya3J
Pxn055x+pByFexB31ddfJtg0OtUvWenNaKt55x3Zx4e77tvr7T5HoG2UY8+Tp6uKIrAf9men5Itm
+10DB/cOzcvkx3q3b15TtnnKMN5C3OTDqRZeJnfkCTKGY3ITuQbfsrWc01DdGTtrxOOp4MMqGrLU
+WDc0drnMzxCKvQlm+oiv97QPt5pdEqdeD2UkojTBZ9vhZyXV53vHqtQzXVYU24qXZwH17ZzQ4Jl
Qg3BeBzujmMOWtYR0W+XiyxXdNtZGVkifVRVP6dCTyGzba2Jl/Ic5iC8fTfNq/eHr4wj8o7q5M3h
R9Pkw7mZxS6c+PBoFEV0HyaHp90RjFHfVpddn8FuD01r47cI/CdDFkV/CPk5c7ojeBwaIj9N0Tx6
xRRpIlwnoKFhfNNBH91dOUMVyXW0ZeByV+xgj8vL6ne2z47FnNnw804xCR1IG9dXrOOmH/xYr/pT
lopHMv2Wrm1vf4NutQcRWmQaTlPCfXs41/fQQUnPhj2HCm7QZQWx2QVVm7kQ9jqLN9pP9mcUIqqq
Ba3YBrHCioPTs6mIWzdU4NiZJoqOQzzZFjgzDEZPs/7IwhXld+RFhIPg03ZNVP5APblZX5tda2O1
5AsdcDJ6+A2NXPNOKn0d90I2c2sIETTA1lczFOsp9EA5akpAegSHsFP/0VWtUvmDFnRjHvkrh3cd
NHM84bmtGxmXLBpmcTtkor+BViOusNlQMTFg7IVaR/IXdd8Gu1h/nV+N5pSoM3BVGXomZ9HE9Adp
W1Mm+AvsL2j02wpN8Q2KckEGXIq8y3CxLbjWl6RExqIeOihS9+x3sV5G4jivAGgHW9Mc3GG7WTAx
qnl//Rk7vcmm1aQk/bEgrw4L6pbpauu7QinO4ybC1BXF3RHchQClZHEHPNehT6N+lG/iBPRG7URX
Qzdg3hplTS0C01JZBj6ZMnIa54rVflaA2mIwWzcqdX0CfKD5Kj+BoDlJvcYlJcM9x/i9IViir+8S
iGV7J9HVHpIDlJ2IbLzERzIx0lw6BPUBggXVUqXa/LZckUQU6y6T62n10JvW4MvRYWuRMXYvhnwr
hHx6nKZjkZ792eMxCXpfy3XzzeN21hsga1RdOStOtQK6ZA1Z5cDEqPNQCQrblajZXzJF9ETK1oTF
CA/Rrxv6RvbXxyYpsqUrf6knFAVjbvxEpokjRSV9cvmvRFs4f/CGM5+iCqOOBnluGOEDHHAJ7u5g
6ghn2oqc5whohcLQC90UTMU3PNkC8cgqx5jhPqgapcJ6UDHUpZ+xaJf3yIVRnyPTj7hajn2dxJng
sIVO1L29Lq+38z+oGxo0o/ZF9k/Y38nFHbb4Wy/njeDa8LkRm9GIjukBgLwXyVG9meBdlzUPn3IL
hpkapmelay6prb2eC3ms578frIOuYzfBUlHF7lye73l3C3C6Z27S3YqIgy8mlddQkDCt1Bv23h8u
Jap1F/JxbFymNaxcbYM8tsTMs3qr9grUJrCySy75V/pyGPXym+iux7WH1faHkyC9K450axL3H1y2
gFcegXFf3smCacIl7/78D+WRafw8ExTkSuP1mnzPrmVGcq/vbrUjINWCMlGPE5F6WYv4cW73vgcE
bqSAtFAH5VSpFM03Anlk8ZB3OA8atXYrdUlPnLyThuGihwjM7HiY1C/koJj8SxrWauOGosukAdpU
TR5CN0qfHj2rq3dzNFq3NWh5aOSCRjHnEAXoJBLqqqbX99U2XhdofU2eLlmRqmNEnN/zDlFJ1rKk
7EC7TvWOyrASpiUMMUMBaoph0i+JCIZbNkIHbeLwGHIkIXH83fmhrnj9+B60ZB+kugq4AEM1irHw
zZAHv46/ByPbgb90wwSB1yFQupM4b93uDWuwVucYcKaxArsdckncvX2h+Pg+Q0Z7wXroXnN7ui3Y
/My68clgw17ChnlelKxCgXJBsqE5qKcj/wvvtaiabgh8MVpa3WROLNJD9DVhMj9wAP35vpq5J1HF
OxI3BaO/qDlwppIC4JO/12ISM1fwQLBByuDEMdirXTPNslslPVVyzBmDbWbfp31w6ZzftGgANjsK
5/xDax9oxiBn4pcircMW0o8LtpA31r8GL5jBDrKxq62iRlrydhZ0DjGEIoSWTpGTt9itQawgOdX4
23w8zy374Avfhg+Ztff+Dy9INoRRgEgx8gGpir9bAC+lFl1aS19yYxrywiMzf/NZBkYcbrLYf3VJ
ccHS4YwFNZC5dU6P5V5FURMK+5NL+LPSzASo/tx8JlOj29BPZ99sX/dAcFeTijHiTEhR0nyKymhJ
g68duo0hpEMN40B4cS8++DNZquH1rfJOBTBfaPkZz/ta+IiCjtluhNlSOGqoXrfVoB7+1h59mUcm
FG8TGkH508Goybzy/t1MWl3hgU3rw015xQFe8HlTw6xcVTVFfj0XRqdARLejJSeWkLBRkDw+X75o
QXSDdkBo/pSpIr5DYWaZHCMPMpIXWtsrI6Sof6myw8AMIcmm3S78S+t/JWlLG/6RVHpT6qOR0+Gh
qgSDnZ4+4CREgvZimHVqjgboHSpxsbBrXHjqO+ptziS4mxEL1GPBF6yMbNpHbd+wnYmRdqXuXVrt
1mSVbbf9qH49bDP9qt5mG6rMGNNjmutJ4IFeH94BYolUmBx3nGNfmJAcjz9fgrk0+9dQUpf7iGqS
LURR+XAh6GIOIxHn7IqD2Jk1t8R9lsFhKIlf2kiDKny47ThXStihvIgfuIzRErpHtYdcoVFrnuTJ
t07hQa/sJ5tcv2yzp5Q63Aj/Q7dAmZA8+uodsZ0I6/FQAVE5nUhYFDH1dAwVE8NM+4SajVERggHM
25B7a66STSwkSUHgRlkV9O4rCtZdD0g7lvB+wUxhxVEVcUYZeIePGdWtWvm+H8xnhU+aT7s+CPlb
skoIGkOqe8BEw+g0KiIRSEX0sTUYtc5JIb+49vYRh+LYlnsMCglXMmLx81MhQPDyCO54kTO/w6+O
VoGCgn2SNoiiq/YDcAsHjbzasiVoB2eNxc8MHvfep8mmstcKMh2ZpretJZaJaYKIAc8+1WVF/LsT
58MwAwJT9WvqnJszM8GEi8m4My5+RsIg8Ytj2DO9H33blMx2zsIVRvNvCSZ23u5RmupuBUKuGpmE
cSirn0jlTsGqDyroQjWag/tHayCoymjeGFBBvDdDvTpRJxyTaE2fl2Umu/GSqKGqmJKsWQfn6wOQ
HQ8tTCAKCudYbsi4ASSrAtaMOIkGON+yk4UAFs6oyg6XMFvN9VmCs0bgVLu9TED/m5zwGpsDOxPl
ylOYhKLkFRm8lYg9yCeBWoBya/ilcX8xowwQ7zehcmja15wyN6dvZmjMX5+HCwD7jlXJynOmKAFR
2EvA70+4BrNsyvs885uYkdV5snivtxe+cemw9GyqIoLCQXtraJesrjT1rCc3V+PSL1W38lBMXsDs
OtpLlTEFPg5CRQ4acpDjUdMzh09r2b840gOiLvjJMszU9piMF8idzfiqeKDF832epGyrfsK1oFzO
QpUVFFWfks88vvqo3lRVN+eI6ZR8crJkVBPuHpd88iYHS3cYKpQFfNGMQx8gJwgQ7FoIDEyOBHhT
exw2RXGVKzxQNnsIASNib2oh5A6rsycYHUVF2/52zBQpAL8ZrSqLPQP8VgWmbiEiKXp6m3DkY5Yr
Bg77z80oNGnhLx0LppLOkHtTJG7zVY2Iid1MX8QtObXJ57e39tVzOKXsmCV3BI2WldNy6w0+VCn7
ChRF0Mb9B4xqDOyeKCyTVEZOo+EOY5Kzn5WfUuvMOgPo/qbF9wjLk9uLg+htJdWGdPu/wQifEurH
MWl651PGFL9NtJ1yPU3fo1XhallsWLNUgLjJZ2VPWZ9GdWxDLqNGht+lnuiuX3I4uxD5WACMVmE4
vxKXq5l4pQwDUvhKYSnF5MzsUtWjn9r528LojoHr6dZe4LfcDfzby9GPyPanhNuyNUKoVc89P0Sb
Z6WguXXYGpeMKihjPlzzrvmdgi6TtwHIyaMF1VLE657YUHvHP8KXbLL+XF+PlXMV22CHoFmyxECl
473/ue3eHEOOl39EDWRzuD6soXHjYCpTpvOQFSInZTSp12Mu34QiQsnGOn3clMbbHbJSGxTuHo5+
pEoxJ20UKk5kRR+OC9xnI6Hywwyly03zwAKqusJnfXVxYtzl3SOt2Rh6Wu8tFh9eUf/f2ekDOtHg
EgjaTkVFtAut+upYq3ZHfxNHdnqZa+N+YIoG1VhXHijIPHPsdPfd962txF2qks038PZ309+q+wvA
CYKwf8kmCWFa3OqBgRsFjLO32HSnVcxtc1Xrr0FX1UsPdMYWXuWRgwd+WeCL8EfZxdzXUxyJ2zqY
1xAsFq8HEopDSUPUr/jVX5cN5EaZO8WWRhF3nkuqHV8b3F0CarRoLdNm7lfTCbzW0MKsxh4zQpDj
VpRwmU8ZNnsfXnfqvIDdZlARdh4v+cOTzw9hJK/V3cEdTczOgGJbv15EbEzJCkT++vVJH8GyeHSh
dr56wGrK6OWaOm/jY9BKNBn1PN7w2QPEjEdL6+seQxzz7NEGR3NQomQ4qLnE2qCDw2hCAAOUbflF
8iIOXp/h0dNb6w7iYWRV5zl2BtG95tRgixyb3vqpI5AdIAUztC0OiHejN2nHGfpMwsKL3he/sBpX
mOfHRNMBsnXufB+qEBCDh+UgqtZOYmC8Vi6T3UjWnpz3o3UI11kIjXRFWcyIduk/em16ewnrY6TX
T87et3FgRv0Yh3B3x9QRS77N5XtcC+jrl+gXCExb9CkbDJbobIGqFCNwkEsCIBt6RDCDs5dX9wiR
9fUD3oj6qGvkMm8swmJDpfcxZpNkR0edrFqlVUdmx08VC6rxlgEJUB3HYs69zUACzlfFA9riZc8n
zWBNtFg0XOyJem1SPz0WBsuCmvdkTt+KbEEHb7iP4Jls5wWuaRY7XZL50pJf6bW9nuTAxujToirw
GmxcZ6P0GkVMZtByUz9AoK8XL6F4ZdlYCbamudZnpoiL4ABrEGRA4qoB9HTTtia/+JocQW61Vdpd
GjYWsm7r6QYKZpH6YYPjQreqRF9c4oLtuzmdh/dSHfu8FXZM+9Lub/ccgZkE6hYeDx9yl02djzzD
oWYNVu/hGKIP1FpXK6azZeQq96wZGjnvzGa7DQoUTZHQYNzwcHU/Uf4v+fnE9QhLwuuC0Pm8bqnA
SGF/UudqSlx/LEhDINi5A4pyKyjst9lxxyRmXf+Dj5MZJggcNmorOFEXcziAySw4+CiLmOopflwj
LwPtaY/tDG7/WOXtwj7Ljn/DaakkNeZtABbU8j1qLqjcfrTXtQhS1Ojzqgx0KAUa32faCcnTTY8U
0IK0c4GelSHKNyOmoTvyQEiSLYnwwSe3M1sqNVIqO5R0vHXfyV1D+OJGA63oAtT3s9zKmfDg04wG
2bhKvFERQWe+yuIb8nIhW5WiUQ0KNysfmWLAu8a3i6o8VMK6mN/a4s688pZpc53xe5XKHHnc4asf
Lc/PxUExs9Uj62E3x3Sd8W9cArl/tkU4bFOhfi+v9eHkE9WmglvmO7r+lTlvd5KazxFZQcDVqJ6W
azBNINYncuGt5zBGxSaAPdAxizyyIfpOTWSr6/qmLeTvQrYVlMpL2ahgliSwtJOB73ch4a6jDnA1
XP8kCrge0BUkxbdPZLnaCYIlU/38Xn/VBkBVIFUskq4IxR0v6lCcazviv5nmSaZp+z3910RPqx4f
37SuQyScSOnLwN8nAa+tp4nTQn1n8pNxVeWeYy99tuHy9UgIJaZKdUdcTM7qtf1HIdIOhsDqwgiz
dDrAn7pQ8ydLLe4SSmuFbRPPT/2Zo/b1clnRv90zxxO+NDT3G1WKmM3kp2fBMH41QXyfRTgX4Yu5
+N+BYcQ9ZxDoDiUNiQ5FLxWY7+ieOvIb01u5ta+qAXTH55KhnDdqIVBGJzCVjZ1t+gLBZZvD40J9
mrj3jX2lYvZkNtMKK+jbAC63yqFz8zJ5kDBBTOpnEA9ftaWeyFFd2leP+K/HetKkS63izf11k0CQ
A+kFuKb+5lhg7byFLCK/Vj/8UfuGGll3/ANpYFOzuNNfimzmBVc+UkE85qjuH13Iz0HHcoYG/Bed
J9IzGsiga2t6aeaF7p0re8uxCH8Y5u8YFXUWLqUCZ+jywHG+m5rLmPsJANk6gOFluyP3+wBzYAPo
QnxmYzBrYC9zNnIVdQfeace7V6RcWos3j+cpnNtIR/zW54tEX44XgGK0OJfVL8u2KSU6UptikxHC
Udz9GRfMJGM39rD7c6XsWXfiuCwNRMKWtF22wr+oqMS9GBkkRwE8NaynCrE1OrxsFDNokYVYeLj+
I1EdKa8TMcDGMBzXM+mIdr1YIgzTzXY3wTx38wzPw0l6hzSvkK2gSALAIbZ5gA/JhS2vnFcWc4Kg
/mbKqSOMk6Vm+s/b/2WQyBosWxA6gsZztrYuBQbzNGouIJvnl0HpNDUqiLyvXGQJTJPYyuoQofPl
0gQ2Q5rnwg6fL2oyR4XOYm36qwzMXATKmH8/LXzBWPjYcMZLB5a45agmxz7jZ8yp4+lys7cf/0Fx
vMSEUDIICfQ8nijDv7WbrBbIi8JeKU2Vy5J+EtO/Mp8Qv59BZXk75Ggda/Wc8Dpo99uJ3ds7BND6
e6UsVhum29zzAU0wMw0eTUH/EYc0Wmo9S8XWw9w4XlchYpU4db6JMKfXaOK2a5lStDpZarIsYmPT
q7kJeFRpkCsxZUagd0ZkvO6nfeYaf3IUKZL8UuqIgx2IyLzPLVcVwPaE8Y1Q5vO7rcvdEbYFTpfF
QojK4XUWA/29F970t+68WwYPPsWERIGNsjdporQmteZ5ygGhHLukFHsWLjPJcHEvMarZC8Z4Jy7V
a+X5hLsTJdd89ydbPcudaCt1rkVwDfsSTDd8jFs3159uOU+lnUrtOs6ZSZDNREU05Xg9z0LW+ix6
btFc0nHM+ALwL/xp37R/bJbLI5fOdyNZiZi8CVQC++8VLFQQHN4WBtdJZHkjBkbsts7Oaagqj82x
GNgvEJtd1vgx+nufcbneN2rGJtolXSImP+dlJLqurlWcct2asN2KUEzMr+gPugQQmva+yYqK1IQY
c48VFSDMapIvZ5L/6DbHMsFfJ6D2X0yf9ztJKergQbilegqoImDIF/nN7O7E+z2sMvvOum6yVj0B
VPRch+dQRBZP3aXo1Qa4HcBCfjg+T/zKxF5ZbMm8W0pLqmo/jSTcO1Qn+fpgYlgEB9n1RLSaHxM5
eRTIpREFTC3Fthg6aHY0SYang0Mp8ytoEnLAvlckar65MKyL30+gPdqsqlo9rynucprUzf8W/DCv
0mbQJrXqm3OfdoATVtbfcol6+fqamWf7EONoLSa6ID9kj8snQnY0j62iXhUD9B87dDxuba722J1q
G4UzUeo9wjT+svMJAzxzf9BzEPAJ0AlR+j69pAilCUKnxYyVaFqaHZrZGCjLw2Jdu4BQRHUw+Fg/
t8jhXMCfOXBKe8j2Nu1yBEmmpXztsURVVU5cx/hZ/lnvnF3oq2e4P1jzUCpUZphTJERpBItIaW9t
Ziznr+c9FTwNXUkMaQ4ZdZW9cR4n6buAQKP5/Zs6RAW9I9z7F5Y07QXo2sRb0CEfTo1g2dJXWoU1
JnvMeo8tTMZAhz/rpHMidD4aEbMuFULgxVKl5arouxqAmo2P8bkq6SQ8ud8jjzSlYeixiKo9Kn6b
AkcriE42k6FNpho0FYmI5u6JOVSwfD9soVikaB1MOEU87NYgkXgwQV+evOw6SMGm7j5knGjRSjgI
tatokx+kybj9na+p+An4VsLAC/T5LJdsEUy7UQG3fppW04CRE8O6Eh6jKTpCYopkQwuYpRndkWpv
H7OwUSz6MnaGem0xacVFJiyvq63z/+D/GbsvQr0wGuEzufDhJ9UGRtz06lYEpqUTD0lfJNGAWDa6
6iGA/DZ1Cn6Aj1k9+UAMKns00Hujv+IZpNrYpnkY6rfD+uLjMfVK1pQY1scP9pC2zXlmUB9/XHzA
nfeDl7rSxsDNxNeHxe/k+gZWqI9rs0MGxwdjAvHkF7UUgKdvt3gm3zdCkPOxKc+MYCwlTuJuZ163
NlYKFPaPXrAXZwjIY0CbwDf3u1rchk/IW/j+HYjPPpR+tbl7JWAK/iLeojNs/RdhYe3ZrmLDL8S9
HzED77IHFrONdfTq86K/q/qKZH56CtXKlvL3FNntWpYlXqJtvYfCS9Qhfo5w367zjeKJyVubJuLj
G9LkZOWmCziZ5O0FIkYmdBj3V8AI25txbz2af7K5IDd5L7DhO0I9CCMqA6sG3Gkz6XhYGvqHGWLT
vXs2FpvoEJX/ul7jRikV1tDYRs1pE9jDvRcl9zUKIi9ZGJNTTkRMzt6wPihBk/O2KuVH78EhiV08
MyHQSjnMo+iWh5FTLzGwiMkBwacRZ+9SnQOmsareikGSNA1DOSbO0fZUcF1hzgHdDlIhORHKQjAq
W8GgfDcyupF9ShB0FSt0WVKtKuXjd6Jxc9oBeQ6o39OkIsQnuEtJXE8F/UerjSvZ7SM3+6kEY7r4
tbrR36WyTvCz1cyWQQvF1ovyOLrrsMjwkXm0ZSg0zxbmxh+FXAX8hvTQ14XHi90TshGTNr19NVrq
UukktDW3vzWPygDBP0WWlJtblVCZ/9OAECHNYmkoUkSKc+XaUoiiiU5HW1TYQUsphc6XY/a5ugA0
r42ScSFhkzF6AGo9YmTpufEA1FpwyKaunu2XyGDLgfQS2bnuwjAulwN1vwFR12clCQb9aibh1Ukn
FLoeGMK77VPqjTuqHf5ca4gPFlCsJNmPJKAoCRqbpci/TP3tnqtk5RT7KDCEPf8mQ4Vr8vvyCHbf
Z7ayLD+cfY4Mu32GvQ12l6euAOKLjG4fOM7PmpKZEHyOtkP90EhI406LJuWLzxtc9jk1LM37oV0Y
2cMzmVr4cJyEQ5CSotNZmA2B3ZudBhTAGMyguU+pV4DbDMxtnBaj7slW6z7dWLeodAXWs0+CVJaF
lNmVcRuxTv7oM+L7eNsn/lWObqNwUj5GZla49/+rXaV5EnVw66wHmMx49QG+ITFmKZzdFI3m+fby
TdoigU1GT4laOehZ1lxtnb4ODbzIl19t13i4GE+8r+OgI5bMFKXbv2Urs5bdZ8O3uUQnAp51caf8
zusGnu5peZ5tKuKS3KylZfLvFMZFkuIOYzCTbClqyaEXy9AzVOrCuNy6/bLT6kCrE26dvzlzefKN
EDAqv0d9fzlrTXuJyXnC1JHWTX5bpNLjRhU3AETALyP9J3ToaKAO4NYmfCL6tPuAYUX4d1EkT2Xw
3P9xTGKT4sEiarxt3swkG05J3tmmRyUn0dJ8JYDzKFg67E9fSOUMb2poTuNpUAjvM+sf3VvjJv0j
WLoYvE55CQ3LJqK1CDIktQ7IsHw2v0hAx94pOEHKttiOm6F34BmFMjkLPVsc8E7p82tGdPNMRMl4
e8ZIjfUufZpEsNdrsAAx5vF/DEDRaEmGr9t1dkgZVbIHe457G3yKBR0ZpLFXcou2WwnQW4BHTAXU
Mlb57bGfRkZIlccqmaZ93Be8mP77Ym3hL/OGnY/kqRO7kLXwKuU7k1eeArZ88CkNsWxiQvUwfTD0
e7Rw6EdJxk1KZ5jdPXrhO5P4PAtFkHtaP2wzQcslZdedA+2oq39G31lqrTVZv6rXVSA+6JWu4P4J
P+PrPfr2srtUzyVIIgk33J+x9QThsecSxveHMwdr9RDbLXlxxm+TdOAqY+nM8QcTFGp83cSAhkfI
V9JTKEAk28S4Tv+376p3jpJ9FI7mVBP8Xgn7d/1+atR9i5to+DRdOBYOOnoo3cFWZqmGRSRLB6M/
ZjhAST2ESlpJKb9aC40puJtLnECZpbSgAv3RT1jyfwIanjYos1r9edBkOUhKeo57jRqeSHbPOZNb
P3FcGaD67fYLmv2ij/4NJUv3BN3GywPP2vJI1y5r+C3GBXpxtuirF4R5W+xIzT+eO0Io5tUCbyfH
FtzpZwoihGyfD3pLTnJhzs5o1IqpzYWXVZNIFk5mDb2ynpxZK9vWA9A0gVK3MNSiInFCLdcaZxP0
093JcIENo64EtBFbf2UzHIrng9ne0QnELyLIkoQsbqxq2PNOagVN2u6zYw0FlFoXwuj0VpbopUVn
tC0BrWJyh+Cic/sqHfuTBN51fNJf7gBuI9TxT7BwqWXzs6Z2dxuvFduatnmx7NRdNYr28UJmjZVU
fXwgZ0qcs+vyMf74D4PCwbpc6/lNqUJpo/uAHRJ0AdpPXK6d3FN3JZ+22NaWBUQckcaq3yzCanR4
gSx7s7sHGkMj6zbF32DjYCRYw5bBI2j+fZ1fXizMO555bpxyKdjh8aNIqsVNn12m9syykYId2jfZ
/KUFu7/1WrvJNucjsjAa8pzasM+Uonab/6C/jRyf4dhAt19H3PpHwiBOC7/9VsXig5COxwicDgfI
ETZAc1qXxDDMausEXwcMgGwWd3Xmm9uoMNQemb6g6bEifoZEh8TqYWeNPfPOzUYYUevuZJuEQtzn
oK911udMFWYtOaCiI2mrzMujDDWYZt4xSc+kDCw9XumUvLrJvYi+PfMi4UuGaCwMdfXiHU3GiLkq
m4LCl2YKPHcCFpmoPi2hpXq0ungc7z6n9MWKl44KxRbMroiPtuJ3bedLx26tCl38/QWXOwDvof2L
vl+9wFf1i2+XVyg7hXB/vn/h5dsJWaDipFhnwz0WxdHDrC7rpMbOKyl+HUNkhdbbINErLwB6/w6m
W6OHVptDd1FjB5SzkkLliAN9j7hn2yT1pmajw+HvxndQs4bfYj3JKLNYGDWHfuXMOmPX6H+rCp/H
VT4CTaeMLfZaDuLoI1/ZUl+AYmCiCvD5R9j+KZR3txvFRbfYCm/MGWR2vFUk7WGXMTgx4GRAthee
yqs4loPVkqWd6S0jSuUI1aBHtFQmewrVSLdM38ei6+agkaLy2KAPueJqTIKpOLn27OFa4TyyPsSn
Gzgy1Y+b/4tUbc/Xn0JlqqIAzJAxmgAuFfFYSfaT3SDi7BLhm+E8OQf4uQPj8uh7+B2pLsYPhdfD
jsX1zP2X2keasA21yXAUkEiJqJ53avipN0fB6dSchdJvMEx+gpxsYkusz25rGZA9lTmU4gn0qogV
Dyy+zfG8ZsOwNvwGeYaEml5GSN8AsHV6cg13ntp4iSod3qrjRkGMOmRj029IjLyJ3M077f5PFjHB
YCD/2St3WdVllHlQ1wLaJ3UifmKmkpPsstkEadV7yj1UsIlW+jk9sOlU+0Kcc+eP5x8EAxjIM+wr
AUOT+I3cbAo64Rb4GPtX1rdsithCq/wf0EkVREaeZAQzMH5hFSBN4vLv9FvF2QYhZN1Sr1n8eSUi
6b8kQ25+m6LW6Zt9Z5VVVw0iDcunsZ57V934Vn2j6VL5IqsU65h9DfI/fNCpwU0Z7RrxugmYN6Xd
przXWW+53M8bnivDML0I80IqiKVuLIL+yGwsKCeGxuoL2GWaxjCCSeIPpokAPkrwMTU0GuUJoLqw
qtVhHE0xqgWkRurw/yltEvgjlardAKhAPe1bSMiMByh4NsN9UUiYu4snbmzgkgMIMNQ1/uyEUjR0
mgey1pm3FyjC5AnOyfPTosAj2U7Rdjefwc39KcvoG/helA1Letr9cBl8hZSpRD3WjT2YA03/uxc+
MvtnksUvfoqn668cxBmUGY/WTZFK59c3255l5gVj5U7jEqEDiuKWq/j6+vsEgRyYv/9rJHHrhpap
0MlOwiP3hInB0ymPMWlNVdUVEE1LYbqKGt/ZApVxWcY23jlZakVNDJBbrHY124EEIXInWVrpzxyQ
VQ9lCMTtzYO6Zklvcwo9FEDmQ00JROZ+Dg31WdKWN7iWNa3OJuadfVM0gTxJHVUuFYMoXCnwESgk
hsMrYG9lwkJ2l4AbPavOXEO4WBt1YDkLZCIJa0sCVD1XEg4u/hrMa/9d0omr2//HlQqiTd4nSFbN
E0FcmLwUxlyG5h9ktdBoFT1nwiYOx4GC6Gb8d+fTljScHEXKwvkANXC8DaaOT7NXrIHVfPN8jgJQ
5G6fffI9RIonOyXOga5s0/gyBTx/cAxhsE9NfdPIsuipqTyDnM+pJXmzoDYuAXqJk7Z/ibOy8KUo
9NfOyyLSuqu54WJSQanyPxX/80qEbMSG3i6cfW+WcaiabkmP8FhFkOM9WsMj1ug0gS0LSsa6DyhN
bbeXsuu5F0jK+sTgsZHYEpiU/xPRHTNa2ZojQGEjSR+aLwfMY1qJ8cgqBR1yFbKxln2wAM602Iui
Zx0NoQPSVzoOW8r4yx0/Y0vHehrjy7edI299FwqsrPehrGfL33wBTGJcy7U3iIP07MXXBmhpEMLY
Op7osXoTOzPwpi9XwJtq0RxYnp1FqczLJWHy1w1lx4eCjsU4c1c/v6NucOZaED2Ckb+hO//ZDzAH
wUevjRtUOOJsqSMnKU9f/DzKyuMDrL0SjednBiPyp9z2Lbe7GJSNfpXkzUL5lr5BDxcpF5FTypAf
w7UDuIAzr4QgY89Eydzg84Yrjn2p4QxZU+wcbnUC7m4+msxazmTUDgSSYq8635Ef8lAL0QXwr2vR
HhDRlc0+4qRli12mnQTDElTlt3ZLwqfgMA71r/HDBB4DhYs5gPSQu/AHnR/9erc7Dd49tZ+NzJf3
nrR6bi18+MqzjeGbP1JHAQZUFNR+9MaiqcZvV+XGuPQxmsKT8ZicQp7RaYfQq+dqmfl0Rx8kD6sx
nW+vPqMdQ23dZm6pe1wQ9YdS7s//sKriCveis4DBbE2EGzfb9QogJ91KsBhXicR8ZOAEVT3XlQLv
xCg39McFgCs1iFRbZcB7WNG/RGAEsnaq6OPu3pPO4/Bb7dcQfHbPnkZBRhtN5syEei9xdLR9YBZp
bDBJZr5TLpEV3jdO1osKn/7qU0J2Fgv5nKdOWf/wquWC6qp5rMrZT3QtPmmt2F8VMVe389hg5tMi
U/SETVgBzGs9AmQqKIdE1+wH520kQgpmW69HtnEN0WTI4rggirWsOaXa23SkUR+M+rRxXutdUBPP
oMKkkzdCKjF4GRkaKBf51aANaoNRP6v1zypzn2AJkoUBEIE6XKhaUYTkgYRMu7eUZ/UGZ9lMOU91
j+YwXcIlg1vmxR5e3tsHTH9LOS4Gd70Zmfj/yyjerslVAKmqBHXaz5vGqatf4H2tiiD8dvqjH+Vw
ARt0Zl6q23fyCUCHnZ4modnLkMtuwuctpEsdH5hm8OFy2VDhibpQn15lSc92LsrncLf0TUFDBiPJ
mcrriQ94t0+Wnw/zjoPJ+KWRYuSPc0bPcWWNXhx8Il28dBdLdRDQh4mPygXtn8uYNFACC3pSsqI4
5p53yeYCzayD54J8SdtxK1AQk6p3CyVgLG+Jdl+aXMsReNc5wYR98TGzk9NaEC0nYpEXxzk6rx8d
hAYEqU1Vf+Wwld8wJreq1P4lCuCb1obg2wiMwiggXt7OWPvSjS5w8eOHlyoNEQx5iF1GTjLuiMwW
rdQ1PNuO7rE5wIafGHleIe6PdfR7c1/OookVunfcVzLCNYuHTKxxZVFBfGKoc1FLlza2kltfDeWc
6OrF/cjGRgt9+hBgnrw8Q5GKVgDUXmk/86BlOAipNwTlWixwbkmd8a9c4RBsaWubS2zWYRs8lDrG
7wCYmV9CkhL2gIB3FFU4qH3Kcqy7g5jtQFmRSCqkPf2LDQTY36x9ah0YeOJcJ+kGC+EBDEpXx04O
1Qb9CKssWAGFqt03ChBfFp5QxueysHKqLqNyQeJLKQBYtEjsw5XAd067TJ7o2NDJDhuQEODoQrjc
DU/7aeEvZLRakQwzmdrXa/qJBFOaHQR16sd4umtbnECLYVx/PRaBB4/+cJDUzj/ZX6C9EX4wY6aH
PYEJ2zYwMdefhzeia16c+adaD0JWUgPpKzBiuIBtpPYL28wGqQ5ldtTzTaTfD6EuAWZh0QGdfyfa
8SUQJ5lrnvf8bSyhgpZy2IpBrV7DOofA4/5w565a/hd5v/Ci/6G0CCcS6ouEn3MU6rJQOV5H5oza
3OVzalFLCScVckiYddeRFY74VLgv+ABK5fEec5KylEeYR0LJOGBpHDMH9s6j0viV3h3wiBvgg94+
MmhdB1CU2CCY8nOqD08piNoHyS0/u88IBheNyGearnG6a9dhL7WESFtHcjmM/JKPEVWK5vtEJsHi
+176FGy9B16aNF8maWXmCohLHyjKckNtdSr2QmX8OMCF9kEXR+AQyaP/oTdPmWlZj2kRhbjScsl+
RPSgfqHO3UxY38tEVruj03IKyN/ghfR34oErZz38/oTsBw1KckCTngQ531SxtVWguquiF66lTsA4
ZDOS2/glO1yucErqT25o5B2kqmeT0DsJTzZgpZljIdFBxIfTXcp5ppRgQeUBuBoC3kLRvmhOurJl
i3lI17hh9u0B6Pc6mKi27Kdr+ktZQAIyDxSHE98GlQ2zm28FZZC+gJojh4V05QWGBqdy87Mg9g8x
2AACejP+Tkbx7fV8p1G1aol8QSXHZWrduH2m4913Ug9s02YhXjRWWGZqZYLvMBU1vxD71VKJ4KWv
A4BbluAgWbYRLWlzYkKd7pd9ceSmxjZ36bwNKl8JQfGnLqPMCDm5sgDNu0XIQ5ZeCd2zV1enGluk
yhyUaDCsm60/DG2jbS5L6djMqHmKL0fPzk4sBRhU05MevsjswiXhoN4mUGgZxyEvuOLIdrGAYlcx
VwlAuscDxqcv+saBbSKyaVKkDhWcfvfU6YoLJnJXgTyMS51kacVnb20fZ4UZYeiaYJuOO3jvov/2
4d3ZJZHfJjUr7Nr3Ya3myS1q2k3E4e7l3aAOYev3ZCT0xgEtjOky8tJV7Zxd4bq/6JiCFC2QgmZe
WFvDLEpA9vjjo9jpilZIbe2c/QGpXwFZAXOZbMqUX5UoC7+rtOhFUuj/tPN9WcRjTnJDCcCxMGUj
zghTsvwqWhROVUVxH30Xw3RTHKuGaxnYgwXy0zZqYlvCGnoP+axhRM9xQUwM0GnoVcwxBnWDuxyE
6FWNgtvo6jmqJakgsBSgk7OP81Yu0PlaGGO1vJxp1VsJ/Fakd7VrTarKPvZyZwDmAsVjAhBUwU2r
7Cyn13a0T3FaOj8PdaxvnNd0GC/h9EO7YPoqjtxOYLhInWj7p4UQXecCMELbvbTRGIMTyRkfldcN
GOjs9OTGh6ffY9oRBN/HLbrlCTj9DtN7njgKkh8o47WLcGWxUwIKZ4sL+6Npq5rfp0dZUpFuiJMY
+BF3tmeQiw4kvV5dNN2qF6rD32HKtcL+z4oYfc+c6j0Dl2nZaYRuRx56+JnKLQ27fqaeVo94AcBK
0Wp36TCV6u9KQrno8vcVXpGAM8YpApfT4mrGDzIbC4B3riXdInd9pucSrGfjTX/bKKz/AQbL315D
EQlALbQbHsSurFny4ij6OICKDopbrsnX5eO1Hk/r1/UDnQf4hhhmKN2mX7mfNhMpm0jWTB9GUC59
QaQf4XKfmswtel7fjEkHGJWSgBP37vZEMJsHk1hxRzoFaS0CMF5rMrHaaD/kh8yXuWh3z5aIzvbT
YupuEEwc/jYc6c1l/v37LvZUiFq5CJxFKOunHnmBI/mU82GezuuUG6XflGfIkZkU1wflhptd0rNi
mS7hQDyXLMr7b7XdSjNDh7mldulBLj+ruAMrx+rgmnzpCcIlG3sNpACfM0Wsb+xaniPri/zjISJV
saIPKxnaYmLGsRuLgsOrZc8mhkyKhW6FEEoqmvwo8wpHNj0zv4UzG+nv2PjaFixIlWzFOcOVjKwx
x1GrpE3YJuG+H0nrJAA0PqQyBVy3ttL4zxPIolRk//V4HUXo+O/hDMC4VMbf51Fn1O8otPiS3H5u
au3r1rq6cv6YOHYEbBbBlUIy+oqygN1KSeoCRkvmTvRE3HxrLfnTCrSAbQGRq5fvxatpFp58cvKi
eYVgEGEqSxmQhqPOqcD10c3UyL74cmU570HbcCw3UrKlBSeTf6QEwPcXQQMMXPURBvXZIDP2rd4s
6xtZbvrvXeN7mXH4AIgADCy6CIk48xkuan+JIIxmRDNVzBPTpKcIjZuu9ToDO6SB2/f3ooc/jUbW
HX+xpXv0byWI9w3Jv+lsYA177sEzym/L3OFBy+Ox1YdlVA8sW2mNYXVt0ahBqKnjiaTck5DBmtMy
eLtlX7gVIpBAaiutmSE58IsWRV3lxrk2MAdh4G/RudPAO5QrEbRIBptcfbNWVfqRUfFP1krUukgp
Li4ftFtm39VjasZM+xOSZySzDkHY9nWMp0yEaqCrzgqlDahoTAVfCuVexxB4IbmP4hXmob4RMHkP
MVIzc3Ld7MHGQ5xInP9fYoPYjRR1UZCq6jAa9ce4jrcg9Z3D0aCKXSMmyY92wtjSWwt0N8r1v0V1
tf4UWDEu6Ofo282CIRXAyMYwOulEob71MHYesUhL2M2N5RVG3/xyY/0kg2CVN3RKGBtGhQrMilO3
I5G//B6z8F/KoOlYnAW8i4lhbCVSUnGuhNyt4UBODGVmzfB360dIQ7xQeicz6wz7LfQVUaJTNAOL
J7CQPRt6zOoG8P5hrSipTjEh31XqmJxGQHA2os7OBrppLbuSsW+jdMfDmv1/g+HF/LNmFxEbHxwV
IxBK3hsMt/PxyXq4Kfmm4Uv69Gw3W3G5qpTMPjpUH0BifynDLThvsxznAFtjZ7utAfe4swH2T82M
C12XEX2HPGs+1BuZerlKuOEK+sCSh66AqCBpLpgZLrdF5jSCB2l044tH8L6tzkwnoILyp/7kTbxp
Net7C+KSeuRED6y8jkmaryblEcregc6uZcKs9FdEYnvN/cdZb9Mce7elD8aF/9kGosk9o2Qz10zA
sfB/iMPO0U3Y4Z6T8gg1Wa72SFNlwS6Kju7FiJV48FtzlrOhqtGiA3KPY7+y4mujuaWAycoRswxX
vwOkRtf5wYt6AwMKlbz443q5w6OH1XFvt+xR6jL+FXXz3a59sCkv3R4k2CSvpv1lXW7HyEwh5QDo
p5QlPXn4SiRceTdDql5ZGGkxoXG2JfQy4Uam+tsytWMhVfhsY1cxF+LL6BAVxI2QtGTurMcuZte4
cUO3za1H716AH4IQIXGYeFReMj64b6ewnCKcUWQgQS2pBI9tfyZ6yewjXK5csD+LP9ieqZdFPno6
n+10XaPxJ5Twr864XBUedsn0e1I2fLmwjnkpO+3TiF0lVxEhB2LV57lAQdarLYOGskjv1b6pNHmC
oa7rJmzFeUkzyhlZaQtFrh9YH/IvIeDRb4xZvxES6r6YoxF7JPy5GOXg8PI0mDM3hLAsa8jzvfPC
GoR1dEzSc22psDhYO/baIeW1F5m2873NqmrvX40weUV8bHMdbuDk97VEn0Yvvrpm6yImRIK3iN9G
WXgInHudiEORzwAWgHhdjMDKhvgt343sN5o+lf9Q+oKq0MQVFqA+efcN58XIUnRqhJ79VJ/5YZ+Y
J55txy3dIJ8mmCXZCSybiW3EukNfXbRP5S5QAi0+JuhJeu/qYvUe84ZePNMPbuFdSSmGhgbcEerg
SAFHIhmmXE0b9VdY5XbKka4lROMrWOfO8e5AMKXEjmppxO8CisfQdxsIL/GlxeDmZPzXN9kZ7PkQ
qJTSB6GhzD73At6KFLKStpVflNiXYjSvSWIiBdZvBRqYVQ+QUpLA1iQbjR2BIGZJ8/ljc/bPs5dd
M9mtFKc+7yvyQKeGaqWmocedublx4cXXHpx80Zf2Aw3Degy22S9kT5nYxoWfIV3geFuJAn5EEfFW
HsS6LbZLF/MmI51NvxUqjKz7Ckv2b5lrcNGOhBpyMiNQ6rKD7PL9Cy5wlaWIi6SdDsyvYb1qlztS
vxfFC4BLsvPBAmhGefTf1hjjaA6VINfCVCvSx9FO298a71h0nrmHiQPbZ2A/7e7iyz9E/7KfN3N8
MEkTqfvXCxZ+HO6drurJ6FCNwmg/3owh1gIguY7A+MyH8yDFTJA9dl3CD18S10H0ekKjPKZYgEXL
RaCgUy1PKu2yko+Dbr0l3XSW00tPK58qCWWNcacdZOdwkljmEGtAUPS7f5tGaaI7blzsrBZAx5BJ
RPEKS8UZyqSrSpoxc5GPk9EzlNDN2zNKl/PYfNpOKKG1rIMSzJ5lQZwOXyJ3gl6VMxduLYpqn8eG
Fe5PsDcCRz27pZGGyS3srrI7IL9N9a9kkJtymkre0y6WVJYqrJjfG9M27piu38UcG3ySJ/81N4AK
F/pxXHPGOH2+yFP/yF3RDTL8zU2OtSfePO7CU7sWIi05LNnfQYsbgA7Tj5N0XZGLEc5WrQq+zNBM
MlgMymmTs56Ng8F8ovN/lTGM/If20fCepCRRoTWzrcI4vigSNbFEPhLYmorNZ/tNpJJMfcxmwckI
hYU6oGM4pxSzmHWca2Kw+CcCuCzSSoHxq87/OzK5UU4ry6CFcs2TS+afyMVHw3Km1hHKT8X02i/e
EfB+IECkYrJZgaR+fBMK58djPJ7LAwGFt/GgC1jYl6KpXPmMPHF+h8jOaisKVd64RLM6XNCkZBXD
g9PkF3klu7HrGrJfyjbc54gmOk+UypfisdDRhlvHikaR5TR2joWGZ+9ggVbqsLbvIMjysja2sYfb
7cHZAAECDZhnA0iEDQ1hQ+ePxl+Je8mIUSt33I7P9gIrC6gh84TKBdZ7S9ZNZxB2RbfTmUbZTIri
9Ao63BT3dXIC0d7VXtc4ndyvbOP4OU8J8ADG3o+0t+D+FNDTg5omxhplSHW71yo6UJDSylJtL8H0
3LVfB962XeHU2+iRTETaU4dny4n5Hqq+HTtc/3L+pQnSHROWC+7ZZSvx9yRIPzZ/aQJmNhEwmXqC
6SMvN7fpNZSA4HH12iIS4/IUD1fFH4aB3CrUdOe5dIxp7P+xnSvwsalwhjFVKuMfan25/OnH+FGG
kZyHtD7ZauStlWRmPwqiEiTQB4k9i3HfGeRpWJwUd96RF02d55O5OlqzMed8u+fw1/5939RquzQ/
GzSfNpQOoHymM1aY3GN9gDcP7oeoMeSFo0gQ/APYH7Z8ZTmTTgtEYbzowMLzCx66CtweJmfbc4+f
9p1bdIIfIKFsNQCSVQqcmHWy+hrDt/DdTm+jxF+XCck8XVnC4KGowXkC5i7dF1xQn6+Fa6rbMA73
tHa+cBkJrvhGBoVCs1YRU52OMqkFsg1JN4j2OFSgr6+L5zrFldMtUaR9ckD7bAN3FiaNoow/Gpgd
deUFDhON+AXf6yCnn7tnNQejlw0FNhjO1Wa60iydGI95VmFpGyaCd3si/EgJBioqHm5wZpnoYVOh
LFqThZoRiCrBwqSbKnmC7QxqMhaAo++bl/Zo3+1RXGthK7lEFpxfOFARdQf/YEYv6hVeVfZZkhI5
iLguLJV8RY/m4ShKoQh/HfHnPNuw2UXgnuv+Ie1gPbcXoZyW3v3o9YBi2VgcQHlerW2bGehS+JS1
Gtf5cOWhmyb0+fqF/4oW7Q1hwmlpKbTdI3YSfVb5isRGQEnspdJ6iVWVqlC7aBCsqEvujFbMdFac
Y8GL32SVtw79bnQyu099TJI6GMHuGD/auFq4gBbY2b5ZemQFtxrWsni1zPjTla2xg/UdmS+UtpE9
2IC3um0WwJsF9vOpwD9bGAbNrntnVxZnyKWELF+dI1b5EjucpVUX/NJRPAQP0sz5EYOU4hUjwHBs
BvQo3gnud6LKbi0B3Ews31X/Ox8eVDF5GNrS3a7O3NNUUTTTc8Dk+kzwQx4YYjXFPgqPER791y8B
/Ad3qASYWsrCQlquz1NUkDWb3ZfjYAjOHhdvXD7LBsn2ZICsUJDnxhIk+40dYzQ9e2MtN5jSL0gJ
jD8FadmvX9nAF2v1LKUrMdnfQ4Iirsr2ZNptb7VAnY9dzJa1bug7pRwkmrWnjsZ9S0dp6sE2I0HJ
88hCuxR5/sLsrI9XJP5Ew3Utbunz/LU3UUmgb6/hYR4Yr3bsuGjnG6M0ZgM2aiRxLNvC82aAflpU
y2QkuT5z7VwFChuxKJ7GmyNPQIwI3AaCqxEsTyYHE0aua4CUXKWsa2DkcU1o3dEo35yRecBGNxZv
8xQyjFky+cda0mA/amNbwYmad37wf/7JRrpApDT6IRMb1UwnypA3gqS940bq8dQl9SPiioK2LAAY
5Zhzu7OwO7aAsfnBqqZByb5g3w+sY7rPaAUOZGzZbK4L+AaODdOQklXYdEd1x+ax6twpiuNwXJ0X
PgSEVf+MparnDiRpUBtwWI4Ngyvx2xNYWoljeoZJzILho3Ul2IOHSEi8ILWigXr6zZLa3vmuaJnc
487oh8ZWSovaDQMYI3IY/r1uD56cBdfQnEIFgey1O/wKnGO+ync+jv4cu3oUyosmPabprYiuBT4f
axfYGaWs5GkSFaXNHsK5jUwvGYWpdAjZzbOekzVGlfxvtINsbsWLyfAIVN1ow3yMLPsE/eq8Ot/u
hDULxX1+Ph6QlL7Fy4EthrQpjk03okqg1hEfzKEK4HqydFxbTQRgqTy7ePuwTQKyuwza2SuiB7B6
txa5sPqGdDUNygc+sy8S5ZICfMNzEB79ivPiXul225PRwbzZoRLJKROYpoNtUFqKuw+3jLzzSPKr
XGjzGhfU6FzugDWAg5X2+ZJ0Ni92F9TTBYjN8kqqOgdVld0OhaNDyiJIQSl63qkXYRDB+5gqGukd
EU/djoTYsjzhlWdtAqeC+b1XqXXVGsAhNd1NXvB5vfMQl6U37DZS2NP1SC2RDCbuESV2Mw/Q9Yxp
UxeBjolYEMj4JiKg5TVgnwb1ZtcG0joQCArDncpNLiYVPvg7XLVpG+7DfkxLXvhCeweopEkQYTXo
P90FzT80X4ebiDU0/eUMIERmvWqXx6hYxRQEaS6w1WqtMkBe6g/Cx0wEmWmiT57qXiDFlPzO5CG0
QcHKWnA+dY373L+346MG0osLO1sBd7Gk69+LBcCfHFTWjLSp2EWrFPUukcJDNaVuzqnllcWRa3cX
j2ywn8yR3M/DLxImNOobr7I2z+VV0U6TOOvNTlseYfNC+rJCubZ7xOowFZYjcjfWQICiAd7lLXEC
SzcJE6z1bG4qj/UFjt/XZa4WDZPVaYXKZkME2V6Y52iMGdlM1jNCxk8hTkdhS5ROVuPyxeAuu1Zg
DVq6IgSm8I7PuDfzz2Je2mfpj49Q7YoKZ8y50lrd+CqWZBVaPYYT/xrwZi1eJkM3BnPFhGt+/ED7
OwYpPaEnkQsyzeJPFBPgsOENHlgbOW9NVRQ7i50pYGSr1yIfzdaX/SOO7ngtlD/Vp7SG2wHp7fZl
IlJNiR6bsdtlk6hA94yFl+3KfBJV4adFylxHhJe6nhKYSReXUuVMTLvEcUqcNhUGoKI2fFSsyEZI
hVc/s/2wXZknCG4MDwTvq7YbzccyKkzLGm0RFMdWBj0pYk47A4IjOzX2f6Y3z4jY4iQgpiIlLngc
hotlKpAF5/Sg8wmaADFtkxeULSxmsHWagF9l2Es/5QamX7nTdxDiqEwGmT26hC19hiG0LJs8Vfhn
0RBChmYf0fdUL3UU5mbYB+YcAO9s7HQPTMr1INZph25Jvfj7PLEBhjpYuuIe01tp8nYdTNaLmRS5
+37iYUCtHBAu/DlHRELEDW+B1BUdkCElkUjxdtRrdfUTMpMn1/I8HhMoa16qOKWbiKRZSjZ1gugZ
I7t8XHBsQH9KppqDx5PGJQe9ue+Zfdaxb7/ArlrNaHmXccOdC4KV3ckzX5NjodHL8khYyZsGqEE3
iFez5rcbn7faw3lSS0fyFbmFJh6ijxOQD5yXLLp7akwT+O/qcOwsJ+90hLVmGk1nmianNtoWoTLm
LK1q9PKCMFL5M0v8pR8sL2531D9BL/BMu6O/7VSxHPIwJYiRw78w/lsdn0sLALvYpJ6r/+5vTozk
Dvk95CuTxYKIC/Na/2s7OjQVv7HENy2pcJmSAlsEYsBptF7U61ikbD01wE0vWhiEaTvYha/RqRf7
mTsI2L899kvMwtU7B9b9n6vUCxr+f7Dpl1NdBU6Nnt/jAvVCMxZF4/aZjpZ9bcZcs+VEEcnD4F4U
YBlimynrJMBR6NSdCwohmiZzZi8df1YYRpkjx3Of+bI7sYn0G5+mKV7Q2yScvHZ/M/ks81FugKcH
YVx90xvvrzYepqycvbnk8pt0FvCXWzfn9hXCgOG/TpOgj/53nGUzNsSCYNsiaPmF7oL3zZObbGtS
og2Ely+Vsa9jGQSPPOgJ4DXyEcHwjkoEZ0E8Y6yqPdv577k70gJVHPa8vYHbQqg8wDoyYDUiOhuI
rGA3UG8cwYm90M2FqorfWX1LzYZW0d/y1KnXyFnpjRDzQMNmqUTDX61PRT2QS9cJnQtk/tVquXI2
Ix28OyFAVRwgHTWbxplBk2lym0W3KDrv2CMweAaP89VsvBX/2n+mXu3KMfe77+UcgxMrZi0kCBv2
v1MEXtThRIKdynMAckKFdcm5aJ970jfgStzHQ84T/iypZnRspYl6SKXitS6rTy1iVHpDu8bc7Acy
gopekTm7Mx1C73udC5rZSaLwXOmz+JuHtvW+F2+V/zA4kYp6P2Tf7ch/pjXlKAr6V6KKnKqLUo5c
yZtoYJGt67B/FhHgk9ewZbye0b/fxA98o9JkjMGXnnKiSojMa9gBcjz1vUSp6MpQ0VeR1J0c9fUC
TqHk43lxrg4R8nz49pPBHiQpD4s5y/eKKqdMd3QmKfE0wvQ+aSIxf2ttB9KwtiLeI3BkbXLhqT3N
4Ym9qr6Vp4ej6oYqLgkq0LEL5vA6yu3Tcyj2qplg6QhK0Pha3tnTsBdnSJtY1J0vnV3Qf1B80LH8
+/JYXxMMarAr9qSmEGbDgwh+Ajs5xIlLCe1OAVhM/w8WWXPtwhEPOkDn4a+E6LCutoU+iJJLvNeY
lwg2NVPIqRE7luixR529tndztLgz7xrvuePfhThllmpDUIxwxk9DYQJBGJ8kIo3+c69CSM17EBt1
yBLAMVmEsvUdUC8NFfwkqozn15mj9toM5e4uPwUe3eJUzzE257IEsBzRJJgjW2/RE8Qvhr6Jiexd
zs6OjKhjSZlk5cw7V5X6zTWBgxqrUnC139KYbw99Bk31b2RjTIcEBLL0sVA2qWmCEBlj/PGVRiAO
9+cAIwwcMJ/U9a90zYm9mFTRXNfpn+cqXQgKAcCfoCfp19xixeljBi9fz9jYVcA2/RNBfGFV3R4h
o8UE78fs28O8gvSLiCWIwkukcb8RhqZ04soF91749UG6nLKs8RqZ5x1Pw5+QsQZYQP+Gxs9TQJsY
CBlVKGq/hZQ8Iq67rE+dcYF7rDnfK0e/x+jc50TCpFwuxKr9HhclluYhl8StIeQHO05VRMee1E5T
H7A7OZY9x2/hHscdMd5Zva/kBZ6SlEKbb4vuZSIO/nWUdN4XE37Dwyr93/wGD5N1aSxgqHpq6aE8
chj+ZWTtDwQQpJrcqoPcw5Lik7XspvrUS49hXF5fLWIFsQgxJS02hSUbqpSp4nZyyVdfOw3JJaE5
LoQTd/YP9XwfcE6j5R3dmRCatPfh2P8AfrinRO5F6TjnkKO9J6AtvL2yeR0fqihGAfd0Q0SMi6Vb
bN/m/KCjit6T0GLdYwJqbY9Q25qwu3cA3eDNpzR3NnaF0w3EYZ3QVL5zKbqbEBE0w17HXR6QDf8q
kfTNOEzULFxfLKVToCWu2voJOI/xI1SFoGHTKAOlgZnl4ZvvdHh80JnmQQPcZc65xBj6xa3iZjle
FfZT8DyXlAQCFTL3Pse9aBWN8R+ZG3x1wiSUhaecwmQA3hViTAtYIUXFDRdDh1ZCdhAB23crufuD
YPwrmRprGLLilYbfRjOAJ3cDv0n+3X6Q2a58dUkHJRStny/0ae3MWy2pNgKJ6XYyhd9SfFseUMmW
tvS7/j9gHcyDeWCmhBUztSxFmcszl72Zso/oEsZHxNeohHXpze22wb2gBUKWVyQNU5sxBnBcKGa2
0huS4a415C1baKMwTWWz+R4W4Nkj59wD3rf7xlxGTb1gUsfY/KSPJiKQSzBJr/mnF3CEhjrqSPTQ
O3xVn5lD3jjMorfg6w9rS9v8HDEVSIDKvWPB6VDcNIl5oyyFJ3aMqLgX9kmtFNx3UHrtMU1JurAz
AGsJXUqh5oL4XujFIE6Y2MwvP+ep/HTNl0cZRe8yBd/6hcG80jMYSsBW6EcshG7ppx0sDfUbbLui
/NG2ncZVLgRAxZz50RyoHVW9tEUA/NVPzbK2fHqZLbjhG0EgTlDvx92EkrOvM8V2aWS4lTZvmlQ7
Z9A2devsqpu6zylzzibKygIQKK7H/3Rt4TiX8VvWwiqotVAl4m4d886pjpyDlREZVUuTc1hRaTkV
dBCSAVuIeupfUhyZBz2UeOfRpzbfFGpftruJV5i7sDXBZtG3We3DxPzVc4zNK/K5culD/qdZYOXA
XOYeBFvwTXICDLUGslfP8EzcuRMrHYtpzqQQE71XEW0iBWP6T47obw91QaS+YosfRC9az60n4nt7
W/MG0tm3IgxirXlqi/Qzwu14/tF+uZBvySKAcoZKS3TzJ4jhNifwA7cUYZyYy81JpgAMXx85V9xM
i+41bVih41ssjMM4YvCaRMZaH9ulICt1oYjoIOPxYJb5WFKe7hmR1u/KWh2cEIuFsuuIisws6FTr
Df3Jildltd2jkVcxYkvoegFDGXq8egrr2sa8rg6cHzrllU4zJufcb55cdHkJKgNZlwDvYklpi/B4
KMo/0Xtx7AOroS0ZN2Mu5syavxhMSgNtqxcwavHH/Yd/LagIOrDLhvpR6e2pGhNY9tATkSbh09Z5
203Pd1JRdY4kWEKG+a/AHHDJ42SxEh0VjpvC5vp8YU129S/4nY1HBzwxXAWKgxuqUnvmjnTxb/cV
AT6AePZu8ExoFpZT9Rx/rk0zRjbqUhG2aK5GvzgiyOduJ5YiD+Js6C0XF9vIB9oOu6yTV5t65nIQ
LlRCSumjYWvSQAlrq7Z5e/K6TsCqfz5WYxFAJ90/Zg4lphpMzol5QuOh5R8C/1u9RNpnHk6Z/ex3
ywSPxqpaqAafKcO8W6trFUYjUVR7qAjcQSzOLVpmhKbIlR1g99xW+lTNmQADkBU3e/FXXBeYtlyG
AZT7E1OmZlTP10AyNryjsbScqyaOkmSVi/B77+EYxb9v1Olt0/WWMuciQWXcYukOObcauUigI+Zh
4ejz3859hBY4AK+BxR5GOoHOb+mn8qhy2ff5iljIo5ONBUYkxbNudtEDVITyHY1UQ2qq240KX4rX
4nLOW2C+Iie7JPBoKknJGY6eeDLImP/3zDfC3yKTouzTd6cyqzjMxCclE5MthyCARWqJ+SB/N7pH
XT+11Ra9f1Wz0QX+LnPcifq8jZ9t34cBOj/hJxyzhSx/rsgAvcbSY4fETmu2Qgbc35U04UikJfr7
95NO04mJcYx4qyeZ8dIwUHmqQbQN3AQBFPAiWbgMf0zFxMR1Yc8vIuIJuj9X4ER1fiarnz6tQto3
DjYc+EFQe5HAdcRYncGTnvmNUtW63qG6JS+vzYNfaajN/ZU4KblWljNRPB8OUUhK4L8QXy09rtIL
LnXZxE45qWwV+8LzgMZr0+LVQZNj6QvbGHwWHoDndUclIssW71gIhT1unoakZ6IEWG1l0uNMfQQ4
ia7qpfeEgBjv41XdjM/mx6v21Bcp4JZ5xgQQD/oeUoy4QuqwO/aS5jgiiBee38AJpBaBIwu5dmIL
suKwKqdTDzPOvzx3rd7zTYBTk4Y9bMcPsGwi1unPpF3Wqt2Epkjdj0Jlg0clhpL1jVenrX2sc2iC
6F9ye2dLw16+Uct/19LsXV+LhpqMHCH6l2p6APfiE6uKnWpC88Psy6BMxit7RRfSDhlDVMpXH/Gu
Bxa/hKoEM6mrcI+p7JYrhaG4u+j0gggadQfYAj3+vIktyN5GBL65WNAhQofePRcAp87wESYM9qXN
3CCf+dVuLFu2XUJDZMFn5lXVinrMUH92Hwq0hdtL3kCS2EJ4I1R5dAS3YxCwQM8ZdmmLO1ZUOy6c
FCfHIi3SOtXZe83FUX8zOsTbjqz4ZNP/guZ0GfZQ9BQY0l5BcMJ6ofGPYdMbdZb+5RVDaWxzBX/3
GKzEvMgwUyLsHH0aNGo8fPMON/FD1QJXEPQBPTqF7T5KnBzZmhJzNyNX7kF1dSDzPGnZGdf9C9Pk
PnG+6VgOfQ8jW0Nu0CrENaJWOWSLFWOtMRVnz3/Z6d3uNHds2INKccup4uo+thav/1lfBms5V1Nt
xjFClPSagvPTfftUFnYY6mc8ap+BfD0vRaq/y/U1K5my0mXuNUUupdAKgohTM+L3WnqHUEj78TFa
C229TmgPuKKmfNLpHwaoLbf7qf6J3zBzXVYMtijaR01Dn3t6xbcoFlmj8ALADShBn3kOosDJiR89
JLFDQkeJvtx78qhsEsMSfJZ/jEjSKoDtBv5Kq500/QEF3YgHk+4LJfOOIhlsell+HOEopC/UX9cF
ed7BZn7S7CT3ncLgpq+8G7XVH2mhIxGxlSk1nOQFIoyo5oM9uWz5mrOFPiSyyIpj54pP1b+gXyO/
xGHedt46GAkW4QajMALk1pp1pXyFB3X5w6T0c9jL20IOzcLy3OmSLqXKQl5gNA28obfBCU+LRtio
+vIM0pb7+wLBH46fOkPraKICpKd51/36TB6DzLAZ5Lm7fzNiPh6OEjgA1tsiNfTeS07hkljfVtAo
bXH7lk98h9lD8Gh6GKjopO3IQ8l6JsL7xQZxD7Sl/dTC/QyMYUgzaIRZYlaWgbjt9dyRGDAmbjRG
M57hNg48lLALHGXtXKwP1N8G3qvRFH9x0WJsOypYpjFN6SpYWubGaizsrS4bmdAiFb629mQJ0gIC
rCYatP3GR8rgf0xZrbsQti0iVc7Ss0Ek8nD5oTfrlCEmSEsLmCAm6cTTRcNGyZHUMzabQny88JWE
SeepRqKDqXOe7jMyOWvjR1LhPRrRyAOqTXXOlNPspW4Glls/IX7zoFCeB4Tor2UqBJHc12xvdJJ4
1pRTIwV1ziBkRrD11r5L9FkI9+jInGL95ODV0R1gRoSNP9idSD/qsnTwhAIgQQLdaEF1u/dUO87k
mYeErf1vgwMTzhoC86ZdOaZUDNmyDOXuBlHns40oETNmdCsP1VB+xUON64AAzZRYuLj6w6Cm7G77
EOd9J2jOWOm62rpYPrPLyLhBqPhcpowToW+CYJbg4M/oicGy0OOAclyR/lOKoyHu5OQfLPxVzvUI
njiIsnrP13QUpaFjQJ27PohtSyEty4ZZ3NX/6rth832IADOf4iPjlCsp688uig90hVkKrPDw1PED
qiajtfjGBhfeslTsD4Nid+q0t25SEggilXOf+ONB6ZN1+2ekHJbiFdQdJT5D5P0Y6xl8mURkHOA5
F/O65FcdkSqqpEuFtEZR4pDntIDKPOvmPZDZe8KvK+I3z9CWvZHTWxXWZBUutK0KT/tDIZ7TXLOy
Y0OsjVQ2pO9jpLjlxlPrJnihEU1W+mwvwIP/+qdA26e4/0FClwQw6ioxH+1ePe/e0RpZNALXPvrG
2Kln6ul14I6JjVCOik4hiI1/tg/RDzugk9oEqnrQWEOnNCNfc7WROA2U/t27TyWvfTDn6tZWeDDQ
wCgh6dEa+abB9TbHnHSB4hrLaIvtl1TJVD+hLriMsEOJcfYXJ6qPsbWNsEKet23rTvi8QKkEG4Gh
l+J4cSRWgSgrrOVr6GUe1wKwjUaO6ErlFDyN+3wQSuyTwXXON6QyTAoBXTHkCMZvrOahFuc+zfr5
ty23zJPLa3mWavVOECReVc+AoNpTGXE+tfygNNqnaKzZCcRm97SiyXASK/s5pqCwacjq4+IKvVmH
hyk3YT0LoYYAPmGml1dGlsR9nWm9XAso2A1BD/+zkhx7qdrOlxM9ldAXJ/aZ42br9RkuyWGRBv7+
WH1QtJrvGXrTj9YQFCf9rW3+bdqGLmk/+QPn6Ua++Pe2YWOzXxUv+Emhibz+rF20aujBW2+kJZWy
7bd5XSZBiho55XNTssU3fkfVSPcFOeBho7Kki+xDLrtwJxKte3tKPpGThpOhWCDLznFUAXXRiaM4
wOpKEzLkB4eloq2LXBOdY6ojeE2/koU6RShdWWAuteHCDPlyb39OBpL5Mu2KfHzI24nc3BXLSI0B
Ng77mNqjySP0VOMjwuGrlCE7V6JCKk/JI2we5xQ+Fuu/5Ne6kltNJxx7lvmR2amfxcE49g58I6FB
KYar8cfFbzq9aC/LJUNNuIFm0gn+yyVk8AWnLhwYrNvIswe2EEI56ad0r12JhXQ7gk4cMbCcp8S+
wridSviOtAbKUYyMmQsSa3sS55SJl4QW/YMIRlAFGJ/OUGlZCqH4yP6gXRFBWX7r4YW4Ep3mkrwn
q/BRGFqCASEcH5RAtEjSFI4KVkG3gzUs5F2OsJ39CRa4371MWAi0xlFNa3tYLngn2vdQPEZi46uy
YJGKCCFWkSK15jfAHADVursrd3CG+KROHICmgR7N0X3xpygPhELX4Gijf8f9QeS9ws0PlwIc7mFo
J7s9aHBdc55KsP30jsnxQN8w2aTsdwUHByaO7/QOqwlSMvRr1HUyz88Q6saSuNpF90sPdJ5QGxei
IiJFUfOA4HkS0pEioEY64vbefSxkWYaEPO5ZBcHByspkCvgiHxBPkOMjXghiopQ0MRUHCTLlIGOu
tecYYiktSx45u8RfDqLiJ7LPO0w7Yr+jV0zwlQR12pRqrZrNX6/NNNTObq+dhqKOpVdU99ErZxkL
tQAei51SVKqiyyBdSVCZYURwSj2ikBVkwdzCDe1Xx6iaXuIdEVi60+f8X0yHkf+BNYOzQuci7APJ
6bhGxE3KPB3cnAUg5D+OY7rekJ5o1u3wX6DyUZX4JM0HPFYxb2wg9xZHFTglwqcqA74AdT1XxPsF
9m5P3WnwrU2e6mvJDDOLsiF4VrMqXxjvVVkZPLsM5qWrvAF/H/391rlJ3LxpDIHRjKY1sNgTvBsi
f+2GDzf5APTRzQ+E56MCV4oXPOxfYOczZYNrpVRxlCytVbGw8MylLWqlYosA2x9c8FCpNSQATXMZ
Cw7JkQO5iKxE8VeT0dfUel2VB+ahaiYORC7SsfArIixINKBUucP5uiCjkhZ4D8oSTlfMnQfaOTpr
1wuVRtEv06vZyK+eEE4BzdBc1jcLTpfr/WJDEtlL29sm8sGYzwdzNmN0HczettoP+8/8/yhvSWnf
cvhq4y7IL+lHPp6Nh3oVtMD9I10UvM5xwWtNsIUNkWfYBtLsi/aAJJ8/NuYYf/tO05RDQpUDrYKp
pDpjnHIqqVzMrIHMAjDDEtBP8K4xsuSwZCtYfNAsf7iPmd59MkMJczaYH6gYQEbNBfq6SXvijq+p
lR2k2j/UfIQZnPPaiprAJliU9h+sArff4QqhFEf+gYR9UBIQEvSq1Sv7K2gsm2igkmpDYvFtrAft
YPuisyv71sEAY+stqq1qpQ03hH2M3AF2fvxAzWAO3xcg9XFBZY2FmmvF5cWShRgqqd/3tPhCGCPy
YcVczasm5H/3I0kUTDVx80xc7mcNtJEdiWKZlHGDZwnr/FFn7dN5107UsWm+LGsQGMMzw+zWSLh7
6Y1+F7NGPfhWOpQYhz52TGAe8J8WJeEVeQ5sqNzR78bW7ydjwDNHjql8o7i6Y/ikb2fLMfEuUrT5
JnQC9ZpaPnTNiCqdE2LlDc7yZ0j1ZBkczJHYWX0C5CrtPk1EfASeLXvVrvWsPTBGkXzRe4Je3tqr
mX6xpDKC//9yImloo4fx7awVWncMCgZyYmG/+J3p3QlAdtz0mfCejjylZ+UIr9GXGk6AnolTxNZZ
2u09Pjj9YoLXLl0Y6JYV8kJeIvb22jd1NXJhlqjxAL4HCmopH3xLLsjXKF+ut29hzIBiBTIj7MeY
0yZZ7/N9ldsgqZnjqz76WEgr6rgNVXkkWZsLzZtHX6U4YOv3LAHyh31afexU8rnj/VPtCHNiCEb4
oLeRygpgPJiUmCOpw70192exbCYIh+x/8FPEbqVltuDVIABNbnpFZEaRD8khu7Y0Fp7ti6hsTYqx
nDEA4gjUQfux/DrUXv4YL0TdpD6XtBlCU1gJ5QNqQolcNzwO7a8Qz9ThGwXiVRucoU7m7PUdOwQF
qFND33VTjxI/NxGySmJ2Hg0P6LsLvel0p5aZSQaxp3fxe5uVM3TR903oFowK/Ny1A42Cp7A9HReY
OOLGCLNxm6XJad3xynIkoaCTd70dfkCehcFAXGKD3hduhIp3qPurEipXcoJIuZ6NEQstd7Ba3pwG
OV2ghFEgnz1Ym6pYlMoZyahNWrwFuVf5HSEY5vl21qooUii6S4ZvNa9Tcym1RpPxvbEvZnxsvx8n
rhb4dcJWFVFYTVEVAV+vvxelFAkqDr7Nf2cbq8+K+rYFrg6jw9ao6rmf9HxoK41KAfTM3m1ylDEu
9+y1liBXla5Y+BI8GllbzjqRQ0JxCQJdK+u3pkowtjswDu8uUGQBTEQ9OULyXZlrQnfUp6DwbEtt
9ZazJr0vWpB4CTqOvgLhr/GS/7fQsiYIDvZUCSxSq9n/SUBJJn1kxPgbc4JlHvFh2bqeyNKkOZQk
67JdoRN8+KN0hmvt2pVQhUzLVtSXEJ0L6b0c1a+2B4nR6eBStsKc8UfJJIV+laBz6bgQx8VgVfdW
3ufNqgYCs7pNfGkeTZd8mGMFtcrYQVH+P/vfh52toSGRI+0v7jkGo+/uthuFlB4+Btdl+mgN9Zex
H89PQ5HjFcM1fQyDk4Dswq5F9KGeU4FIipNFs1bYkAUSvusDVIv1vV6EP6u2hxN0zRKT7SPKTQl9
bm1cLSIqf9iTEpTWRkTX5PgvtNb24BZBTDvieHtlfk7vK0AFR8DPPL5ogXgPEyN6tnMNwWVbGW7n
tREytV9HHx6Ngmt3NHQex9Sn6EoaSRgC5aEf6TxXL6/D6eZ+98nYEXA9yyqCoVy2JkJ1jHdCdT3H
t9DpP9cdtaEIu8nk5dfh7+u9qFoPRpg51vmghIHQHUPOo68lbyKqfzxSiQ5owNHy+OWF+Jc5PQCH
RGk7NjSsxk9m9OgHnXCy8j+oaicblhnng6Hdi1sWbmNBhRP41XNclCj28ue0RkJSofKm/7RGR3HD
/JH7jx74x9RokbGRnVLAjPHPszSEuW+wQQ2E+cZQxWqSVkUR2tsfKVprKA+ErpDzW8vybAz8gxIC
bp48ynLrIZmYcWQlfs7ZrIpNLtPQQtSjgE92qZCDTFwYiYmI5tudnLnATlx8Zy8gWXEDlxKotjgO
7Yhzt8uO8kaksVX5iCyCfiFElu9E+C/h9GD7uNbPqqqO/RExjr+2W8jKpNSMdVDMoeLncPbR9fyN
IkX4pa7Di3VCANx6lyHmu0Rw8PZM22Zoc5CcyHiw3USH+GUIiwqdEx8e7bUMOkWAWya+B6PrE59+
KM2jdiCbM9mqBcz1KrYSdqZ1pIX9b4+LIjYAHLzIoDpv0SVQkMOvlzJR1oTcoS/awqFvAIXWm8P8
cDtM755biCD5AdvvuyJhaT4NI+uWeOThiykfDNV8UX0VcpKk+6XGhX7fnpimhE3MXIs4VBN+oGgs
i8BmXoZeN/cwkjhlAEzCBsZdzYEAjZN7VEslp30zapFKXGfpxXZZQph6peXBJaK6rMBECTtUvUVp
jzxkIFx62G9kGgbgxsahVJaYYwENmZyHDBNkwxyJes+Ha97IWgLSkRaydMaSKpO5gxEzvd9as+QV
OMA38kH9JnRiFFYomF0+eY5CNPyi9/hqjY0zLl6113zPKU0TJSVuRnn62SeGHcYupRgsdly2sdzJ
7rHQsiYI9Ltd8WpR2hxyChHYhaMspopR08A+Og7C88IzxDekX8bRdFNcLzoh4DO0HOGM5OhneUYI
gK+nv31QALPAKhTHQJiexmqhUy6JkZCxm5kL1gB2AwHQyYqY0hE/y98GNXGET1CF5mOnUTc6Ws8o
z6VFIaUc9PfCyx/u+qLpEv8grQCfjEFP8QUnsYDHytb8BYW8A2nYKSsEMdNa7E7Yw4HhWy7RaEhd
SHAkcZkDRlQDxfxWLlBhqwoZP7iBdtNO2pvyA9M316OHmRM8AQVfnBEL4/qfGBjz+A+d9EzrqthX
BnHvLHChWKG2oytwgdV3d8Vtblc3d0wzSqAvN4jOG2odB4Csrk3KkPfST1NpkGbvKtEWJ4Sq1fB6
8I5K1oagrdjr4/k9a6GKOVpKQ5o86+KVkJtJkoh09b3x68+wbBYko1GOPMiZNGxVHDgG2BpQN8Wc
oWrXXmW0K3ol8Tq3Skgi3cwJHBRr+juKGl3+jnrKOn9iACSCSB0izTtOEhOCRNFJ+qonULDDNipW
6kO2xidwHWI6uOYSS6SmbIiI/LH1Y+x010n2EXmIout2XQPk23FePspDhcNkn3j/67msJXXOXHyu
ZUU3/Gjume5UHru6VKNycNXmwZnKOqKLuvJBoZTiE03wPHdL0YZu1p9fpxwdjZV1JH/wO7oQVRuW
rv3KZ9L4nwZoF8BhtyA3HWNJCpm1IhBD7SZt302wBEacLC/sThhOBTAdayjrJr2p+WWMtFuGyNZJ
AnJwJZowtFZ5dSzgeMyvWDtlwwZsEWxHhEr/xIYIMBZfNRNTEWjtkNgWp7KewVMfMt79OvX3QKQs
9RmPMlkl7SvprmvgsY2uNacQ4J8b6m/2hZG4TbmQSbruLPsivgwILNGXpDq8nXO0TIsgYXjc6ql4
yjwgUV2g9QOZsaLounjI0BzD5Kqe+Eexda9k2CisyY2Dcn2WvyCIZpZzn8w0JyfZoS7bmPAKLf7o
JavVSuQuhfdglLCAO8c3tyUIdORxtbIJvM1vD4OgLUPL/BTKB/nqkARBViyZ0L3YqkDP6jsCotWn
llCLJA3aR6YS8c7gIfLPoyVs/7LNFvzFe8VvnSR/JGV7MpwsxwJiVqDjPnPLE5evUvRkiRpZBcaB
dyPwl2k9OQ9UPMpaySls/51e2xrJIo821dbwTBQeinH8QP6MMVfgyHOu7wlhBj8RtIA4EFBRad80
n3BTZV2vAxbhbetqx9hYXC0Bl+Udj6I0zNevJfhD+lWk4HW5kQJdM7um3JyW7RrUM7n3YSXdv8u8
N3bicLIDpdWGaa96hniAYS4yFD0KOFERg/ywG7bzf5ieJZ3ksSrAPvMtVdV/kbN1w9404X8a8gI/
e5Qn4ckLdqGRvwhye6iHiJjtmObNypilwryAMlRXTa5ZN/ne1g7am34GxQ9eSaMeB9QMSe9HnlOo
5PMXXlu+vrsjFBEJRxXTs+CBm0Kl4N//WyxaTc6EOKh8LH2erQnWVs3SYwaY2FsVDoYXDjL/JKkm
1unKDBpRvy3YbL9g0hdjWR4LsmPaif1aZuPMyGQw6XMaCPIBJeUroholS++eLH2dd3qlGzG9Y6M1
HIgLUVqYvV/XtKmTI2SEAnySH79r2F8gGl6K5c+kjsQF4vWizh617DSzJwX29yV89kAh8euxClph
vXaNPMsZkYbxu+A5A6nphGEOf4QyfQ4cMW+NLdH/DAtwJNxyALmHVGtpXD04IQWf5kgWbAWMc+gN
7AIgfErF2T0DrSo+5mJmzH2rgV+iW50XHCZjah1cg4e1nuGhtqo3O5Gn//ELHk309UaFTlIR2xPG
I6E5gufRz1q6wtYZzJAUJ01C1nej9fab9rQQdLog/mCY320GjKAesLUd4qgKyUptSVjpLLyO4Tns
JOPUI6RGGABxejl0Nttu21bFqXxAZnCOCKozyghzASaf+sDL9sSqwPFDUkys55nx4BnLR/ervhUI
kyeONaC7sZqHHrOVko5BqUozbjYAvodEhBNWVf6j3Xt3r1OMEhIyGOxLdQE4JrG2hXvx/r3yTnWX
oWZASTRGc9Kv9WCLvJS9RLvV5NVJ4Tr9OaCT0YmgLfoWI2CFlLbOi9qLVm+xQVN68rS5FdBGuPmq
HKLe61XYh+I/whF5aGcI7+tGsUuCLZ16CK64hhSqV3yBW1/GvqsFbttnMAffJlU1BhO01VGWDv+e
u5Ql9nc8Zn/02u6HeX9SrP7oLgpH65G8nD5+WlxeHaaCgsm5bkOVwTGhJJzRbgMAC04055GFTlrX
qwL8lnG67qSVl0bvhQ1SaUezHbszNR6b2GAKjxH5iyCcyyrXERnKCcHoYT3UQmsmAMFw+wTuoogB
chBIkW7khZSeIPwcGFgFtB0xteT1zud5I5m80uvLh2CWg4OGS8+yGyxxtBYSVgTP6n+CDQon2oVN
MSmkVCtrBf2snY47O+PHuMp0Av3gR2sQE+hX+VtSKKj/7ZYcDT/j5Wa27V27jVxgzjsXLdyBmJD3
yDGTYRrUr4CU1W/HfDtaWi+uqGuiAK7aO33IKMhsE3aYNCPhofEcctyQ/iV2uYYjtvDAXq5Vhql3
oUW8R3lupfint+Z/2CDpjsp/3SaNmIBgXFei/KvWXCpLl3ZJYtz9SDHRkpgid5j7QsOEJkudYAl/
/vy1SOmn6YmSdO4aW+UcBOe7gJixe6m8M/QXnky4H+/jOZhv4eFoOaNl3Ipf8fXWx8Fw0EPG1WaB
3UeGwvXrxmXQQRttm7LWLpj4CpTKyyHXFLDEtfTQkHha/vUO7L0NigTI7d+wMiPuUIYShLQO5I6l
J4LADy25zdQamFtzCnMqsYmIKZbMhbfbjS135L+XNLE6H3heK6QjGwV7Yj9J21T6cKE0T9wyDwc+
sID1RcB02ejea4gXhMb+J7WMN73XUkimEy+LhMJyLtYEg8MtzwCpti3veIoaJNEtm9SNV3ynyy+C
/QY4A4tADYjCMbevlMX6cirCYpR9U5o+x2PHzbDMqdbgmFfCrARU1FyYrl31bjZyk4+04sfoRMbo
JyI2UARNk3yFaX2LXVNCCVD6yGa+/afW4NBHRrO6lepKOWlQJv4GCQ+z5CN4LDC3pcx3NMZtcv4k
vmfnOFyhkRCGR+AZ4CkFKakZyM+sJXf4KusOCC87WOtMO/Z92MADapeyltheil1LAXPxX9Evy1Xc
sa6daeoO7sCASHBTsk7MRY//bQS/dW/sfEueyC1qf0uMixPfT4eOMVq42+PW8TG1loPGFOJinItK
595DdvyA/JooiyVe5nEiBMKgtMdFl9Za/G704LzFBpenS4UV5SuLktUylr0AieVATgL6+R3W8CWH
Kuc+dsjfAzZOg9q3yh0g1r+ZVyPmch4gwVb4A8X+Ll7n/52j4VOhgFJQwTYUUbqYqjJ/x0b6rfA9
UwhqHevmbiBRf6Bb/UnrGAMu70UIyfAdePuF0w1PwIRMN5UPSZUWNUFmnCafSdVuVW4cZ7Mwth10
s2P7TRmhD6JEFRjfIARuKByG4tQlfpaxHECvDV4mAxR63YDFM8PgqMzzUbXAtRUvCLzbla9mIKM5
M0WDeba/e1Va1Hon1sKPFXWyo7vpHWcPQYU0D+t1jmFQjcFHxM0JQ6TPvnezfmaSXefh7jzFQZSH
RXutDUJxdsPvJQFQ1YuvUUqRyvO1tZFwY88GRCc8jiuuCK6bzLlwTB3tdgmA1V/Ft/UReS+NylYH
iW6ZjS6OEd55F2roLmkaT3pEdxaKwTT+rIJRi/OhtZzna4E5y8e/z4tgYgzhNFIjnjHsAx9wWE/7
ud+u4wayHqRRzlN7kyw4ELSFXUkLWmWvOWvIrXdAwN0Qwxn8f3cX1WcxRM7s8zRXiEZ3JDry9mCz
5wd3mLExroF7URwHili4wCA4kWui0+MRE9qyzKSpGG97GxM3a+77AYTW3tRYshmpubVOgbJMCLdz
mcS0qc0AISsoixsNquEIiSQaY+ORhnU3Hq4vIKwJf0Cm4yRD5/zMkHayCGT9rDxSFpG1NaFrWyfb
FulZCn/Lh8uHPIWXr7zz9XGmuuKIAzlrJHA/49+xxdOfPOLVtsMCCt7jacceM9KhHx4sg/6y3Q8g
zovif3Elji9Qt64ZelKwznGBr9WlF8foYKrSJQ/z62UH+IryoNNvSBk4aAy3z1wAjyxPGGKXD2DJ
3RQzk/G25VxvJ0338vPMSK+0VnxNvHWSI1PKZAz0TTPlhxcUXWuiudwl0Iq2CuSj6AxjzeqxInrr
N4yQVi/aS5Irmk2zo6bck7oZFjtnKBc9wdthzk1Sh2Qrn4hykJFDcFthMj82xk47PwyiZge3t3Hi
Nih+2i5YVyXUQ8+2syFSOhflSMLyb7rq+b2mb4s48E4ZFIGLeVRE3i3gDmO7kKMb3G2ljxlX6lQc
+eOjX8XR7EhHPmOu2huVm0vmQx1JtV65pOxy5yHl58Mu9G8pPBQow5VPR6MI25Q0j+CD9w+0Rta4
T0p9GVeRwRgKLwsxmg0SGNwY0ro/OmUc2FcI6cPuE4X32zqvTIXxKZgMxdKniGsoZHXfvAbPLwAf
hn+mEw+uSa5q+J5KOv0cgQ5zGHFTUhGZJibKrfhcmUaGzvWltsWI4qsJw7zJt1BLmNbt1gp8d1np
We8X/3Wvtqoav8MMGHVoCk/+9fLSS823fnynsIrHLK5+t15ABJWmKX5ZJCWFEt/0IEAi+wIwGsIw
yP7TNqoE5QP6mLJwHJKad01lgMdLag5C8RZDIpQ6dWPz/E7VgXOcw7m7Yj7yGDrSsEW8fq8QriKQ
LYqHUT3KbL/Gtg2H8YtX8glW5VEL5xLGZCN0pyplWn+EWk0ny0TlH9Is/8mtaovu45hqZglpO50x
3IHmawawA5bvgagDuImiq+C39PmogIOCaIoaejm2qfAS98wbzF+6v7hpiNcDg/7ZZHgdLaxTlsnz
S+woV9trF+7we49RuUYimm2qqyvvlgdoHRrEMBMFzk1H9btaVjv/HoD+64hnv4OAARjhrURC7+Nj
20k8WiYjEsXZuoVsHoFihc/cLrEh/hqNCfG7AAgB9ARwphvSFEYej/2eVOpytY5uihfp+Mu5hxAz
YK1AB4Zc15YQMBIf89QukVEy2glN/Cz2Jh25HyUpmTLIcAHLJhMQAlIwGdUnfcmkL4WJdOlkIIXg
BkSKW/n32xfSkdg/hDlyzgebVrBKSAI5Z21kLxsJCQ++Vn322yL0gpWNOPP10OaFZhTAZawE8954
XVGT96fh4d+PaWEoGAo8dKrvfyXSrbwwbX39V4iKBp/G+4nuZjFlCZ+/PbTDC3NRi3z8lGrjdkFR
6T313flmCofUuL5GyN64t56WpguRsh7NbDicwmdJuYEUJVg6xpwuRFUgi6K0ZUM3Bsg+IZBWVCyx
/rxTixWG6zEiSQKj3Tnm9NgewU/KnWK3qj5R/i264MauIMy9IfCzTGRi+FrTEtrS3niwu0FRZb+3
+av8KwbtF0uYa+BDr658MQQu97SgwohlKagMtooR+cpnjQknhr9lB+ZCGD7qSYvM/rHAUzKSPadz
5sfgcV9UKl2v1zGbD3jPV3grUsdBwWOjVDflrfLtbdnldffrAvU/gBB89crO2TsrSCC9W3Q7HteT
Q3lz7c9XpJxu1tkrv7/tf1UE8PXR74HoU6PkV370ulu79LXBYZ3TUFIx72QZUoN8kHb8r/tJRzST
44qle70z9RwTdsVUHTF+55h1hpXte7VbWMK0bGLngPBqivaBYkd+B02BL27i/ndWKf1v73QtcbeV
3ebx8JT0LbCAvgiqXFN6yMjmeOHyCz3Kb+CI5oHdfpChNGnFwiFKrp2hIMvEIDyoCGJtrp/YaCTk
u2Ae0pKGTyCf53FnYwZ5BJnCTTTVD9env5odk/ilnXo+lHxwryg1gn1RtqSHrLOZqRSzkkMiOjKY
ZaNaKTV/4Qh/JDhDJK4SyK3RAThOlg5iXBE4C6+hCSh1bMa8CqTtfxEg7e+I97ij+3yIC59hdwku
eVVd4RTRQedraUHwEI4kqroma9gErckZzz+3ufSQlsPO7lh/g75CGKvxalLGeU6d+GU8d/Om7XRR
6pv82Wocf4Pr+7190XAgGQaM05l2gnu0wUjK2UFUsxMT3u/BaQdJyX48o8Lm5QBwh2B6/psCUn9x
+ilYA0qoc0PriqP2i3DfFI3rektrByQ68be2cHNa6c333Fr4v0LgIKXyq7LHmD0FAiv2QAoRLUxf
osBSin722RgI7b90s31egapo0j3LFaGi3M4p5y5ZfBEXAMlON9hXtl/8H9XhOxcvSeop7IrNZ9sc
Y0YBzVSOS9e7Tgqc7Q6nPiVoajmo6rqk/+hPC3sOID2cMbNJ/eXAF+hXK6zXar/31SbLBqR2zU6M
dzN/avZ3tBhVaiiNCjQl8pxrzC/IgGoAOq/92KkH2UCKBcohxOelygsyJfj6trAJ/gJeLZAWDGf8
phyd8rfI/SNsS+OdvRwdIkbGvvOrH3mR10HIhERwDG6of8k2uyNTiBOxZ7bc8hRN5b+R+TIUqrzk
y3vGGngex9J4gI04X+t6raMlORiO92cKHG3J5ZNWUdOMFLPOmsK2Cf3SXzTGzVy7YrvKuYli7bu6
lCLSBths35e84mlG/mmmS0VYFg71sK1pfAlwryrwKSbkYpVQTn7cwELAQMnPFoPGvHutw3ddjhJI
Fxz2lq4T6mWlj/Iv0+59qqh0Q26TaKg3BEdNoiZzZs4q++6BsDtrS/i0bfVc7ldIaoJ3qjNUFbVK
5PKkzRH2dzY75fI2A0fGSC1OKGWMmXzjW2jFiJovo7OCs3icBMb8rInHZVhDfXSZTj1XI/q3G+CP
W6FtlT9ksEHiUhXVBgXktBoB3T0QnBtbjulI1rEXENWbJ9fPKpalSCMq3A1zcx2NLjToh7ikoXc0
T5dze098gA9qke/Ecez6XppIA7Z3XmaIAReSe8eYJWdUQTtP6hrMVMtWfNDgk289CDUS1qk+f/SW
HDzVwDM/jKZnvIC2MK9InHzp3NVHRZ7eW0K5s9dxfzQ/j2IbQmygWY2czQ1UqKRm1F0RtPPCiIou
GO6CLJ8cao7rZw5TPOCHARIE3ADDWYA7WLDW46/z22nQJt5a0qJ5yICxRvJQGiOCeDsHVsFmrIA/
b0YMB5Z8YFxhwi3dqlrMvhwEgkHPxll/0XrcRvoFu47SCawaKo2Npi5gqNK2ghHLmMec08o5v8DW
NpmsUo88cu42GLNdYnlmWO1BS0cYOGdUVDKhQqaTuzTY9m9jXFBQZZCt6hKMkofT1jNImHsfdXYn
UVFygS82lnqyimGQvxlObXIzmEMahwR/O1NPHpCaZ8YZFxMGRIpD6G0q5wbtL9d8CruBEt3tg+Hv
VRqTll8PZs17RVE/VQCKLfURyby1DlXdOdcPshOHMMAK48SFcqtUuKeZqwHgXogho1F32Px++GmR
KhDEXbRpF2n0MBAfhisrfzt1+ZbKUjvHE5dEgwyHHKzGZAUSDQ6ZYID31D0IjqsGd7mCngKmfLXU
2GHx4HkNAT/OQpDoM7wz3zLO6D9+GbzR6I/Gi+m5HAjw+RhUsirz0VBbzkQxkJXyyIwKbE5y6fU6
/xWxzYPzP24MERYi4cuQTWCYkYRTtr6AZ3C1XVkSd2S3OHPHXpqDZA2h3jlDQgaNYTUIy+DV7xtn
z7SX0Ez5hllZGEc8KndQOlp2Dc8ZTFyqN0aucLQ31TvLrLyzEGn9N45RkFU80Vt3p/haoFF1LVK7
nxJj2fqd++DPWO7sKH99zYGcevr9PZDipCB8zaZ6e7uJfys0MKaR9jcvauhawgCYR/AojtN/lm3+
e9O4aJm+PTEz1i9q75ryFJg7QEjon1hvjIX8oaDlUZfq+PzFtV9SzYesQKdnGAqjSUTpQpwPCEeg
PtGj3aJUHArIvDbGENkaPrOXy0Av4v3Vyq2Y4Xd2vAR8LyUXaWNDqmUTNOMd6UdmMbp11wjRLsLp
qOxC5HtWCC7iqrS7azvPXZKb63Bye5jtz5Dc4Ze27eCv6ZzMy8MMqqcT70Xo2DRT2rjc+ZqgnECE
TIZM+8zOonk6LLUUdv9vJ5lMrkePPLlHLGQVKB5dgZPq/cdX0qK+PD1/G8kGma+aJaXvQ3RqdYBK
Z2TvUR2r4ANnuQnFbaQraL4s8mfmpg3wsSHS7aD/1QYg3nAZRGGgDEZDe2ZSS7WCHI/brDhFuoQ6
q1WouN6+SLaVRd0aejVz0f5W4pxffKRgxuDrZc5zSfFzTIfz+axJl5snGuGofECkos3LJQyVUEtN
OJ/LSjLVi5xT0ejT8RblKqYynHRiPmA6z2Zz0lU3Re5JNBX+HKMBtEIiESF99z4dwIhgI8GOEZBz
O5L6y6f2qHPa+RZyd3eJbaoSG8+9Quo6VM+ftMaiQgUsW7Zf1UMZB67Miic7NSOtBY5d6Q09r3E2
6Jl6gxFjO4xtd4kiLUK1Zcg7Vw5XnWuRRh8FbxfvTMz6hyafGaC4MZ3TVjZWa9S8YHCpPCkUNOjc
kYk7KhJ+HyuQbczAk8e1+cRLdmxjywTDCY9ypFLi91y4IRWxCg3a3vFTIc6JL6X/1ZZ33suOy2l6
tU8aFP6FIwm8Bw343Nq01b5tFF44+IKNI6TYCTE1MFEcJpkklgt7qeMI9HUpq7Q5PHiMRQJRvEoL
KeWhkc4ykZ5icZ+s9focSgxy/GgoZquTIAWKNiGUg5I0088PKAGkdZkMyAwUoF7cy0q60gCgcm0b
pGkvm8ASTtjLvplAbMqBYxE8zNXY5SZ/XyGqgGIFQed+aXlpMO7F+m4utF/0uid5F3sWGI8hIXkI
BsLvax/pqj3nuErJzx6ngFvEgw0XJmWEUJVNV/1LYK9SGPgwAHhefPR2UBMV/j1zScAmeyaSnLqI
bN72XSIpwNKak5lu7QKnNnfspITmhswYAErdL8UwbVFSfxInKELvv2GQMRI/MJYP7KMw26IYtEPz
10DPwOi1bffY+27hWc+NVGoULV6hdMvAWsnTKmUNFikROS288sZN27R5/ZG/bqe1HmJmRP1619nk
pYVwvaNtE0lZ9Bhowl+ic4pwek0vyGMVPW1jMbG0R774DTLTc4TvwvvJ4t/qbMMnwCTF1wXQs5/h
thDzwVxTCGuThcgMksGXQU3Y9W42BOC3x0V2fkwOcY9MoA3sUOEkM9BsL84R3e6f9bwtJuK0foMG
XMxTLn5THTSewa4cYV5wHXMGL/H8gq6S3a9lvNP5J6ZcgY8wuWv+hY0pAaMnkhLT1dVrALLQp6HN
NVN0L6GqCRdqRpBNj3DBFrBg+QM908hWUP1oXk/2f4CkqJLjCTAfNhSoYdFGseTCNl+TMoRkf4VV
bcnj57aJTwpLXY/T6iQms9mdQr39CWwy3kGwCSQ95Y240YdVbqUrndSHgdW04gZy1jyNp5dgSS6e
x6Rks5zPQ6apPDuIjVhRqDtJXbJ4w/T3LAO+rFjedbYtCJJnA1mvnjTNEgiK0ZnuzSnFjkcY2mIQ
NEiBQj01OuFnKiXKv+vHqLQrF4uOWd0/yFsZ1wPzdUqGJPaVrhAepp8WCCVyO2E9AjS7udaa84t5
U4bU0SnQn3LD1zckioLGM34i0LcVLu7NEz5J3KpsHkZmXnOhEpzPhVA501912t/0wEmqIA2t/vKH
fRRj7iW0/TmRDGD6zKqRuctnhP+88U2lzoVBNcHv3DzGKnp5zOHEKxDUBh9HFPR1aHGyUURC7U5A
i/R6WfXb85NUjNyKBDS15LKgaE58i+iePxztOAVlQK4SQypKHkUW7RCSo8vySdIyWz9NHypz7taa
leGqJ/m/2bv6y+n9m89mn/fwlAXB+LAr7+8NwjoK665lpIRSzIEesaUwFYcyxBwhSn0pwWH/wOBm
0AycMm/reJd69TdhPQmsAvKTDQoL2DP1hNiuCPwrU2qwVj+7erj6Lvuw/s+7hmTD6635srtkh0vr
den+Gz59eaHcZgNCwGZ6fX/hmOPdWZ8i/7scM5MdIgIMlyZ0t3sgiYuitWUpJJ84mdyld5+iNIC+
XB1Aptw+zJjyXodilIg/etsZjb5Xn1EsvqdQLr/zAi/aDzDW9GI24HBaWNx2YHgmgT+5wSrOVroX
QEy6FoA9jeyA3InuOW2oJV8gWfn+mBhBrHIA44N+hp0y0k+dHpp9rYQQgssixvnv4rjrO9rU0rJ+
K6DPPLnH4x48SNU3n899iR8Om4QJS1a2RDFsA060bpiATtjk4I0OAj0TnVGVvvZZJFKtsmv+BA6y
j6aNl4omyJKrWyFGq9Q8hqH0A+lobk9pBUz1Q9hPbOnch7RwCJEnijFuSoK7JYv3xB4dvIzqbNq/
2mS/D1AtszQhoKmgJ4+A55OAEmNvlboSFpTtrW/2m2vvvIHWp2egFfl7QFUjU0Xq1uezOH1loxxt
TiFGzyKmDPMi9BPJKi5OGpJrSvVAJx0/Gcax97jjGk50y6fkNylUOfNGWczG8JwDHSfuEH3KQizw
AnqjopvY0Wvj6KF4yPHIaMGR1VYYlbuBKqgcuX/Gt3CEHUqLoYU/m+JAq+r3ouZfkdLAc6ua7OD3
XCUcj6MlP583Uahbm1VfSNYu74H1dO9yKaIdw85mJAAchQJ2rEmUpKrt6bvDoI2oMiiI+wCe703A
G0okwgCSGmCedhUdrlhT/8sDoZy/8Z+PwnAyPAe2RoeKQcll6ckMHo82l/Kc/ReWS/ZehYal/Fbm
9H1ctXo95K1xObtgTj/G2O0klhTCuZm7ZdhTWlOsijTuqxE0eZB2rFO0aOHPKDmZgSziN2VdJL1d
VDlXCNQbE3E9gBA+ypPHPeARxaJw7SSyQIJOzFSQXIvDBS7UAyN5t25ZtRNEuC14q/s+f1a0B5uk
GGfNJIw2KnpuX9lU8MFmhFyViq9XRuAPRbFyX73unZmvchUptDG+sXUYTujXUwo2Z/EA0Yob8Xge
Yt/nvlbvMd8tmr1aunrO1ZrE6uqs2yMdAdbm413I1PEisSnS/CoYSD8F6MSccNBXISR/lFh8bPSg
/OSr6KkPvwpQSVGbchtmmiFZwdrTOOS8c92CTYbnn1/gD0ncmqODNTs4P83nL5i6va4AU8M/5sA5
Bn4z3l5He9U7+mYs5r4s3mpRTjxliCdq0Amg3y/tIpjA3mf24jZehHIcSImkXL7bMLTTJh1W24YD
mW+/TRNTw8Kack1JIfeMxy291K4FwCDUcNvV57qrtn+fNc7romQ1EBJLHhjZa5wJWV551V4xTdWt
lz/Ez2SqIInNCkxOE8bb6Efd1EQwMXg89ykBma4LbGCXEdu3SKZPRlefbYJP620PgtsL6edpJ5yq
Y950kE5UI94ry36mNlv6WOaGuR52iqrc65lq00MuT59KiyEieqtRpKXAAgYshHC233+7g67je755
TYI2mIYFq2BxCe/bLvoMNggKBZOD1AohW5SltwUAzC9kGgMBnFbzgn5iaO67j8TQHQ4B99ZnJjhK
xQe18tQVADswO66Qy5B4SrGa/RL7llZV0AT+CIdThE6Kw8EcxqqmI1MoA6t6aVHTLvhjMoINmEKw
w947HAb2rl/IG0qytHlSOdbXa08EnSk5dIe2qrK7tftb68HUUE7oiyNLR5AG9fioqS1NaYzxz4Ha
5RuLmMsnqNdMMcBFSzyRpUYhJj2yfti0TU6mca3WAp+8eoAH4fBX//c7t4jQ+CCjyzGL2SnqR4uo
dMGxRd62aQCcU6wJtc1DUMYA/P34aw5XdQ9PXllHozCwhD9bc+901U9k8p52xJgQj0VzX3g1cC+4
aPS7kAZzmTj8mgb2RTYe879HgdkzUV47blppbbRPrUBUHW2AnbYMhm5zPWBh00RZ9mhzPU7YDA3E
pAClWZULni8r819fHsfUXYt5VHt8gDgKx6S1eIzZD/ttSZKRS07WWkxIF+h0wLmTjEpf3V5y0Q1+
J+xSIC7ULrfUw7uhasDP3jMIAwTDuZ3u3sEY8q+WOAZqHFs6Mlt/JULGNdu/d0ZZJ7OkL431WzUk
68YH7IvMNZ1Un68NIhr2NThe9sM9kenXnjwqHx2UBHeF8xXLvn6pTOMzUa1vc9JwU18dNEu2e2Xg
KDTWYOVC5fu10EmQcJtYxLwW/XZ006SYiXEsM24DuB5dl7HRWOZv16qdTWSOOOZkXuGS4axwpsw3
z+21uqoxZjRONrJnQ8qwFvIpHs56MOdUZN/4Y913i3F4IZhrHyZWkCBB0tIQlFKnPDJ6PoU0esPv
4A2oqB9FdEpF+3pcSOXeV+leXi/oP80/yg1Y7TfR2xZqN0VmdVis2MHv86vx1JxBHjwJET1a1/hI
aYbm9AXOP5BVPJhGqyEuwdpTarJ/LXqhbE9emszVXGuSF1Ss0HJ7SnzSZOI/WJQS4g/R1MvrDAU8
gHi/juF+x6VtFzEV/5p8WlNEqT77ggDt42cJhRxJLBvgSlrh5aDmiJdnBfkbkMLzNNEu+MlvMS12
VBsFu0cj7K1sgi5r2GweoCitxMRv1uy5Uf1TZDnxmkWIMc4ZWo/EdQ6GYUoJe8XdcDEWidpGImVi
V7QwHL7545lxpwysSSzIV/YfdULS6l1Z+dWPevsaFBZMgBZPhhDRB5aBbNCggmtW3As++VfifmUH
GQtgr5Nwsy4exiDQcfNe5lVfnbYCUcACGGtHqTmHT5KhbrcOf21kfV2c5u5mv57Lo+TJCjKr01/Q
XCsFeLSisrpts8e4kuAq1gYW4T2X1BIzsxnvdBh3QvD+Yi9wMKuR3Z08ao7Cncsl4+/PLyiHWr3m
xJPD4FpUrDw/AlBQast6XHZjKQYojUqytKsMEzAfEiv8DAckIo1uGBUp8/sHjBkkzCdWdu6DHG4V
njy25dSeMv0Tn4Yhii9D+7jkxAtTTbghST7TbDfwIYc3Ks6Z8D6ogf1DPVbNp76WQHezvwhGXmwg
IIsaUFB2HVJFtpE71Ld16CsH23p8dHz5232XCraNM2hxJEgtuyuhaSHZ5fL/jqdOLU+zCYo+0wYD
gJjDNB+K6kwJ6ZKZJCM7fKXVn/MNTz4uUuW/fq66PApPQDPiYwsPMQEscNUII0J/FeW9dd+u7o3R
iVinZXn4hXO99BG3W33aILj69jczo9GxGtVdNTWnQ7bPx38saXSpnpyjOpl8ghDBGgYkld1NLf/0
4ts3kZFt+jJeg3ScS1FYlXSZglhRFKOYi8Di7oV+m/w2IhAMinzsfyaRlzLb8e6b2o5UNYIoCLrk
Dz++c9WfOoIF/yyAGATD1NE6M7IQXOAvwf4f4TdwhJeoGHeR6pPyw7QrfJ3kjLzXefrEv8hM0V5Y
N2cDdfPhdMrNg353aC3oG+gpEqPSXN9Cnavn86blyba+wMD/wwHOxM+lo47o+OXhlfkHu4mTGhQ6
/KiWs33r4S5i8sbL3SlKE7GKhbnSzy7dYo1R5dl/WyTtMm4DF6j6O8m4RnumVXXQbwzJavj0gVJI
jFn+6xACvdoBEhJ4XreCaB8S7Vjz3Skd+i68drlaLPQhQCFCRp9054pHK03MIbILKTz8r7B93aG1
jwnHDIOgNh0UgOGZ4FyobUoodzjGhPaOCX43j0pMfaeuz3Lbtv04eIcfTF8G8Lpp3yPJzhRJGH9o
MzJsEZRrbFzaU+urley+xyrh6fpnawfTMtLKvlfx/p0aABTUV8za4QQP3WZTuPuuV63XNr18uaE+
aB0YuSKNpaEky8YICdqCnNXMsyt7Wlv509V8l4cj+khEUcjYI9gQ8DbRgCnUkc+Nz/xUtRAFaPZc
c9zFyej0aomdPHbYH8HAPNV01V1dZ5TL0qPLKMCPBZvtG6gDyH2qU5Dvj6K+4p9NnDsg4y0s3xYt
M6JJroaDZP3v9w20z+1QNh2XqUYr3bETWYDxh2GHeaFa0hv7KMjqpsGD049mVj+pZJctBgv06pQk
CgMji5XkSUfsQnAqqehdiCpWX1qrFpTi0L8WNh8xFej73gAo0+L2ppyE9VpitpzBxr4skQU4SIYY
ltQKEWWSrrre8xqinJ4LsUySAC5R20A/VJs5qzzcygqwLj+WDQups13trkvQEWWu1swmj9UV2yGU
RZKe8oQNsWuqUw4Day4m8ynKQsTGXpv2jimxMO+9n9SAfTtiMHOLVz3ZYTL2Y8OnS30DnRVw6PKo
4dpHZI4JQ2JJcnm38/GooE+mJA+Hg5a89UqTPU/PZi4BQ4B78XzB/bMLXIsiP1nGTEiObEGkPW9a
y7UNiGTuefHRkwSnwkWFKk97ZJ+pkMzx1sWsvnj71altnC1TaCN3+8cAGc2vmS/IVfRaE74Wn/bU
rhpGQOa4zdApUATsbKjkARuayLH64dDg5jBRmWjwN/Hmz9FW9ph4IS8EiTTtiVa81aNAr04U9TIf
+VIiuvZBVBKrDTh/ePedlZBRbaQzjAHtqPPy5bEG2v2lTeBq0nMYzOAwqpdmoH+T+fKlvrJ6HRzl
r9m4rquf3uus+9e7v/ERXSMv30p3Y9h9jQ7bOb/Yz9cLFmob+JEgplJMzqF5It+KCkGXCcxf3Aix
qMXUVwsRjPEG8US1XcHMiSi59jNcWUlXqkR6b9K1w97FQxIAHwAupE2Y9BUPA8A/hrZCHOydK9Rc
rXYTVzLtqq9YWzJcNawZnHBEneq/GLQxEZ1sRiTOwm4XdadvwnE84JoGb2lZa602Pfdhh+naFvfK
ulEou5QwaRSqojqicGG2IewwDjOh08B/+lhYuRqW5x1gmMBLBbWut2TTEntbdoBVWotOMkJ8uXVX
04AF0+ad3Damts74kSR8+145YAv10FVFYkOQqQYcLLvL9V3n/kzHi9RvXKRZUz0XDOdCng9RWz+6
1h3kWtqL5V/ElWvp4VT9kdFpDj23jVExq3uTvd/WCHWltONyNA4iilWZBZpPd+v+gJlEME2D4Hlf
So8Pl1lGDqmhkCUKVhyD5AIReZmlrhrTagETImknLbr7oNSL0xDqIK97WOydVwZGF9pUn31BzcI8
A5rtDCu/jh5e21M360rknGRK0wq9Fknl1KSNhBGhcnOzza1Yb8yInjoQNkpLfLvvUERx2eYxJQPn
eTzi5dlpyeOXm+G3AhuzgKHSmFXUvNpIxlxIN3B2962iwoJLwTXil8/6jkGRxq65mWZtso5XNXNa
/3sLJAUoBJ1HexpM+EPsj0PQ2YryU0/9vE52MbVNXa/YKwyP8RG2oktYJaRIjhWUKVtYMqnin3TE
6lgxog4hjIXJnrKP4TBEG5EEC2stp/ezIyLVVQfx68gFLNTTiUzPRGwURbIjtum6sKJuymxbx7UX
ouR/5FoUBmzijT/nBFZ2RHze9d98J8gvxKIHTsb7q7Oo0/LEQwnEYos80XMTrUhteMz14nWjFZWG
by5OoFEhRk7tHDp3X62ZgvMDhrpbHXLG7prFpNpdehJKUM8WKck1kxyoCFaqN4G5+ddRPPZwWIez
AybldCnKFjADG/xq/oUeSaVyjOWPTmxwug8FXwNWNA9VtLcBLj9aHZUFi1mC8EX5EllzgVKU85Q5
D9OcrUlC7xxoi2waBeU1SJBpHYhp118yGbMIp55P5XMJJpFp0CXNyQdMcxL/VQiLS1QH+6RiRtWu
ElS9/bakLiitdhjOOjY9rhcr+vy9txdVsCMbU3EpfvWnrvMdT7cKe5p5/Tc8dD9bVjeFuHoHc5C9
GWyU9umXedwKufD9SAlmwmXCp3NoBPHnU0NV76ERhy7ZY0T0QNl8D/Gkosrp3piHAa6igul3JfJL
5Id8kJE7XSKagbo/hxEmbTWIVlRTF9jDUCBTeKOtZfwFn1oFdQvihuigjjzAn0HjhBn///hk6Bxs
kBnbNMHwQR/TlCmJMeHeCcdjLDqQO/5Q/+f9ytulPFxBUnE83+1RyH2P/5duKZfMmhRwCNbmkvOK
3KgW/7zIjSilDabdmlSpcIRm+Pr63x8YM5DRMIv2viLdeLK+8AeHlIAeZFVn7GcAdkRhR7PWQJU6
aaLA0aQGAuIHFVCDzh8cmS9E1xluvBqF9M3f8Uq5rp4U+p6AV+J03Ufs0khZNfaTltevAU3QmAma
FMjZwGYLCmNOqESw3XZQlFD43UzgigOzXWepMu8YCg17LqRf9UTH1BqrOcbP8H2cC3eo/J68XIK8
PE//tysAJj/+MjfQD6gbgn//LcITClRs4EEfYaLxg6qcYNWFxm2n8I7jodQHwlmhSSevCOJYhbL/
wc0IGId2a9WOCL6WU/soyfXtdFpyl8LJ/b9XDLqp+vLLMnQ99kp3cCFA4XbGnrtBRRgxb1h3jCRw
/8sxwH7Md7vylNBJkoHQFl42mFTOGYvab8GFrSygjOxyqFKGesupxUCzGcP2C+CAf1INd7Rj3H4b
AvfEDYVIAvw1ZDtpVI12PiOExlPL4+DCc/Iy37Bxc0CudCScEPMSAhzZBihAMM30irmG5fPo9rUh
8h8WacMvkoEDbido8hPRC/8K8kyxNix98Yw0WVsXuPTO0prcPVGSuDYv1j98Iw6UOelZtsUO1iAX
wJwGLUGY0o0VgjI4KFvR/O0I3uVvtPuUGA3ZuLM9Som2V4WukzwvJxrPCVUOPuv+dD/cQsUaeKJi
egL7Ix0y38Hu9uPx7UD0f5oZX9IbWYpiS9BMpg7Tmte9XaEKSl+WoGJu/LLFlyCemQN/3KBvW7N/
wRdb2LtDhSXlMHEJbSpkf68c2fXtuIvWZJdpsbStLoyQ3jPviW5g7wv9MNmzB+XmsxUyPIQBJWKQ
enl5+s13+K+9mhBlt6ROqRH2mio0n5dU3OhbIfzHnZ3Xeb9meHPeVfbBun1x81bR3YAfcsCUi/w0
YIvuZurbwXF1dgnu8Q3ujDkjyRhX44lS4QDdmSMiOTKO1TRuba1ogmYGBd8B0/j2B8Cw2NFQQDvS
LkuKIY/mNKG8i4Wl9jjkAjpjevUdgpue/58twZ5owAEwTZ4Vium950GtxKBmu2OZCBP/Ph99esbN
eYh39fDzIqKjfuhuoHgl56sVQ/o8JqaESZBNQNfVe1G8mc3RfCxC9NrUjurDCU1Cbyajo0q0XJyk
idSlfZuc0k6/mkBfffGWEQEAanlK8Xz0wT5TpaU/kbBH/9pkMQJIiZSqCTVDgDz1mVp5/lV1/KRG
I/J/csVaomcdK0OR6s4vi7mlRO3WHNPugNa/0MiVShQP6ORsCrv5nrjNisY9FFcrU6P1chwGPGV9
/EB6i4o7SDI7gxkMhxicLflXTiTNqGVsUpaDAUeRqQWD7u+sj4fAm1TtdN2NXINW39/WKJ3EqfdZ
CJt4sdw2ORa/RoxcTDcDiA00BYM1BKGRbpia8QVPo5HVs/G47P/sw0Ytp+Zslx2XP3Em10rTjECV
RpQn1bUlMh4k2fp8eGa5Vrhi3y3LZ8WNQzorAwPJmLlX14GHChOr85FRqXbpfcPA7xF2PnYfhVBf
UupSKnCHt4YifnHbAh8lPiBOvQOcPhciN+Xv059JYeIhwVJeXNbODBj+MBPzIVtirfVDwWXXFSHB
ZfkQXXTIviz5M/5SGXY+4lJwP5w4v1v6CrNdjSpItxEGZLTUiQZT+Yn1cVl6ujxzriWNf+BZR5II
jqbp21gF4eLIDp5UrgGc4oZLwf59gWUww4bnTcm9f3EA6VQ929zAo6g8mCbnwaZ2I2U4DRppfKhU
EgxxQhUexRmx/GjMCJeT/WpdwwZmjIsyMzI4v2fxRpXg+1+2wsxkUmjYNiKHa/4lpfbZo4sCOh+2
N5Io8Sn7rqQbBBWnxS8x3a7zdGpohwN4jXBwbY3oissA+GNfl1/7fgEQ1Mi5M/WCbz5wYqvfdCAL
L9jhm29amZdXCgTEKzeTEGg+bL5cwCGg8d4IYwvc3moeFMBF9dOB8t1N0wydb1V1vqTXC1moPxCo
fuNQfoIqCdQJr/nJquYDXKQSB8/DJXw6zGAvd4Tft+JhgeCnO60IEjyjzJr4NB3kDahNtnscXmMm
LZ8ks5ZckeWMTWNoDbJgLdN8NrS083SjmrJkFklPTdeG/zOdLugsYhWAeF411a4G9/cojiFkecid
bwnH1pTwKMsoY1ghh0Aphy0BIKLjJoaYjYL9efnisvrgaNJt1Pze2ZZsDTBeOZeSFO6prIBwD99V
fsI0r3riAFEOUunY7kSYPDIO4Krq67yHiyzL4QH6vvR0VNUKVsczVju4hTxRLm5AoSz4NMK7W+Jv
309SvsQ0qVhMrGIVFj5EJsMunwmlYxHbeLLI+GGLYesJAsN9lYpxk1VYkTYHbwSgTuijtP+6cYmU
yEFOQMJFYUbffClcQsMq/cHirieaQrtE+yhb+bUzvadlzSvy19aEC5ij8i6AD3C2/nhLDzsLIHxS
u4CohuU1BfTSHzwdjzrV29HNb0hBTftSh4ZmRcqm6irBbr6tw/nUDXfi+7AI8R9YqEFmoH9QqW/7
qolRMRKRWHCc1EmUlWSN4tavpL4ndMkp3RlTb+QKiKm1NVih/6p/wOxNnja5tox15O82XGq1O60W
/ku3lOkb7jwUqdvKjUcYUGkLQQ1Y29jZGPts8a4vN7zAPIGksL1ERtsOyoMt8M0i8Lp1BMzpJKrh
knWagk6X1O5nn2d6ba2hZE0u95MGHKQgrW3YB5jkeaEhQMXLr1vhM2Yw3XC7rhOmQfvK2cAVVUEQ
znaRDEO+DeANqo9uT4J1rCIJXZ1ixM67pYXLn2rlLXp4hAUFHrE/Zd1fu0LWtUZZUfplMXig+wAd
o6CXfFd1XiCYjDdTwyVfPawNnxzCEvfygIvqesfEaiWWPwGHO8pTLs0psuS/I86bfO1uY/Z3LU+0
CpYqkBDGegytzyM/V/4kkx8CCPjbgRRgJJ/eeyx//KYbjChYCJmVXyVs5KFQvqbvMqVRcfMNHXh1
3QSHAr06mtPlWr54dP0wynD5vxPuNwJYsaPgp1JKQXhXBF3kSxdsnaXjROTymyeNnrumLvobIEVd
gjI1uzObrA4r+FU+blVS8HCavfayNuIus3lSIpF8MX2Pk2pSRfj3W7bJX4QZ9tjZea6FizPRf1a7
MC9avQCV0m6VetnTS2CzWV0Nzp4acPaIzONrCll/GUzYa18UUv2luSziJtaSCcjliJ0/6HVViF+K
mrbi/GfsHADRA5HQWov7TWm6esiyNqC+Vot1nN93C7lrGW7Ov9IZFqtEexqrTe7ELNTReme58mU9
a/plXJVfxs/oc7qbki6tU+ToHw4gA7+OnBRtzbNAwdzuHudcs+Q4QD5Rztrty06WNAIm/ErS1mQ5
5RKpAKYdh1HpMn6svu8ENSd+Sa2+d2JF4/P1NPD6J5VTwNxlZKGisF7uvJlhZfmWKzfL4tL0+PIa
CXR5ubw1LuBEbhXM6lyuzrCeAc5GkZO0/IvS/gkptiD0D0PrNctUmtSGDIoohWRXPDsMKS18kwvz
DSicthjrpvrKojSlXTC/RAcywCfHdxSpd+ISXeaan10gmqzuQRSQghTueNKi9EA4eBR4JbPqW8Eu
Ra+gzL5Ioh2xAETgxsMKH2wDcsT7toc0ZWQ/nZfbfOHPIt+ib2eDROY3R75DjRiWq4t+YoRv0Tqc
7h7097c+l6WBOzgLWcerG8ijKkyQeK3bc6JMfCnx9pGn+XpDerdouJyRcgqa9Md4BCJh5gycpBAV
ZM8hSJACvl9Grl5kNO3ILw3cMhE/iAdAOLkUmP8VSAYacWL67+mTx1zRRK+F2BB/EK+8I2bYOY9e
L8TUlPj8gliK0DnOBD+LHntDhWxM+JgTxy4xzj71MP6itVG+dYgpUmklEjtswusbCyj29MEj7/6D
E2MLkHlLUgc449V3BVUf+iqyvWD4oMz9hXw8zH1Gcsn07VTcFO3iZBsAPKAqq74XYe1SI3p6K1RF
A6ccj4tLzzZH85xutEA0BoX5TP3zz7WX8IlYRM6w7XQtq3zUZw/ON1zqrLYI5McBb+RyS3+04bka
RGst8RC4wkNXk6/s0dkWkRY2OqCHfZKpDfRtkWEND4WeILAFPaju2tV6SGd8vqV4rfAvBbTyWm+H
ppnORT5IYecLuu43sAUxz5HD1GaXFWv2fdQJPtdkO3xloeDtv1B1n4KnEpFSAXX1VBJY0hMkson7
uVZ9rXajmWl6MjtZ77niJjTKd3cvHVtD6gFxyWBV+E6v3K6jxKK2AGHd1/jyXA3zlCjdCrvtPMih
wTlWM0eI/3xcW1slYa/uiVySjvg99p2TMwk9gInDh1kyrB4Kt1C5PCK5kXjqKit5L7NeST/J7GxD
2PvxdDNuqyxclJZWneox13JM3aDMEQXzEj9tPeiIKuoX4mKOFyrHdcL4ctPCpsW0E/nsWkJBMzta
kr/K+Ooopo7Y+lBBhEUohKV14rGytEpYgoBc2LXsEp+0yETNglp0Kfr+m+5nLThfMcXnxmQI8stJ
M/zeJ3pjj2HgAL/aV9wCduholwZJQkKeGhIuZtcnzBGydK4M0ozkd4sQpMh5avdZRCnz/UmW3SAl
lcuHV/7UdwPTxRX8nXe1NugcZx2yJEY8vj9nLG5SpIU6T769O97VmqPJwAM3KU5aYVBM+gkKhi0R
WhWxZzSGLr3DKfGmuRdtTp1skU0+iwLsswWFbRk1BEiF7sWWmD8Gnsd6v/mSpvV6e1/6z7RpcCzO
r696WapZhwE/nDBRi8WIKSGj79B5apvRj4kYaZwnLQc9qQWl4Rfb4IhNQVnUocK25aEEzJVCFjMt
ZRWM4WKZGEXnDxwmP7vFfqsvyVDuIFNpxgyy//tYrvtxPWSBXYei+waLP8P0k9gkU4BD0BQA3jlN
z4XuRBz5mbghccQrUrSW8yzHj3sVXRdql1Enyztsly3Esrzb/3ET2+buOQJQK/0RRrO0OxvSNYa1
IVlUxs3RBJDtOIKd3aizbBbjRvg0Cijw9xyPiDM7rhKaNDypF1HrDIZF8j5lr8Hh6bN5pZCilyRA
gocweDWcHmEV32s8ydliOXmiFiqLNQjjT5AR8DDoph6eUKwmCTKuApc0yE2sozDKK+E0QnyZPL8I
+c7cja97yUJLvLy2oldnxT9+rshp5UNFnfZRTh6FIjQuH+L9EQmT56eaGqtbV9HcpGGysk0/fZmR
QXf52luybLnXPpbkd3+yk5VJ3Ne3t+R4IYBmM6OG5wJdfBsjiHjsX237Vp+I+DwSEF9tprTqB9Rg
UaIvcRHQu8p8w8El1VNMougB+vzrzht+kmMJN8kw41f5phtkVLENXUZARa+3Gocy/NQIjBPfHApj
PcSDD+WgfmY5yV/huxSUe9uPzbYcO9MctAMNk5plNNt4Sd30kkOxCbt9upxHDEqpg8961pstglmN
vGhvO5odWyohxoPtC7RVqBUzlmbCRq1+Q+pxcPbrYDKDhKoRZrPbZq7LgShqsEDC+mP1vxNVEa9t
Vwt3bKGpG9TEKXyxCHENMCmPwLH1+PZ8CX9ZDHx0cBcFY1ukaWpq9GY8NXVwb9GuaWwHCjgPlRXl
uDYLz3boJx1fFQoReni/9ji0SwbIixINIYag6LpSobHIlydQ6EJzlIa1VpONm+L32f1eXQrhApNV
7P20sM2gr9Ea2m8QE8mp1HAgz7ZQad3j7kCMG2Y4/NputrI1F2dKZshcsD3xAsT19KkgGnquRBps
qzi9HrDkF3QbAr2O/GuHk+RVdvSQ3ESCLJmgDi4fV5hh1evNjrCwhjoqPvCM3PAEOd3BtM5f77ML
A3N8CAu8v23aYiz20nczEFw6J5YXSWuajAX9lwxdlAS00nNYTttNItP/RByWU9PtxOIdbpTtog8L
Ji+KlljjScq/FyQaFmAGexZatYHjA/dFAmn5etYG4/+ieZmyKTdeQN/qaKqePyr9ia6Ce/nfVDBT
xrY7MOLdPsOV64PKf/puJaane9R9wiqEj+ewsrTVJqhQ6v42wbSsvgG4Us/5sA3CaOqIp3kdgrYW
EHugoEVPR6ENhWQGI/D8yLf7khuPVFQ/ORf66Epm9GjhW74uQG/hSWVFGG3Om3osKfb7W3yOVtus
TlihjuTJXqzrvPiM8I5n7xGFTOjBB2VwzAsu5WSZR/yeswgMUQJEixRudy3BajQKfOQNltaEBbLA
+Wg2mlj+cRpBUVCr+vqbEt1GMele1jLUg3uolfEc1rs6uTSkr1GcFWsYgacnEDhK0rV3xCH88s9g
VV7TT8GkH2lLjXoGW57vUfh+PRAIf4/MHW9p0j8N+NHIZ102a5r3keTIivMkluD9QqdSobFpppOt
wFWFzKeKPjV7gizItr381oXD6lfVy3+vcpU1+cDb1U8z5V5CLO7Jp7/h8X3q2EmHtpo+/i6lLnbU
Yw1YPQGix8qAaatopaGJYba4w3N02IU49r6IODtiTMRFgZf1lrVmVmMsjApgg+29g5E6AzSZc5em
oJaCdnGUG8ucZW8GmSg9T5wGk7LZQsL/2RXZzNTcwzRa5zAZDy6jIwLlNrgCT3kXa1k8MYZcAvKj
1dvn3A9OFx4hWXW7x6vgW69qrux1IV/bebftwXSz8VhZU7C9R6FlPYIKCLpRj3/yTjXaBDG4oQ1A
Jp6tlB2H6KO3zNVjuJaHim0HhCX1pl0yfnV8yv+HZ6iX8+Pos0v+qxQGJ1TYGQpi6XPhi0SheXom
TnLOcU+S1ASoA2wRkRi8jmx9fe/0iyq7HO58jMRljBkhE/BInw2gV3L/D2moUoHxEvXeZEYJ8Cco
sWBrQdZRKL1AFPv6C2jFmEsFOuPohlbAotU5wZFo9TM9310yMkzUJELVd9jrwMvVzAl2u8g3Wrvd
OsgiR0+ca4H8LeoLrRcrRt98XrF/PFD+EIlX6L4mPw9c9xlSxXqbZnlNL+P0140eDCZaYdcKBdHK
3oxRklrJXDy+bVVwUr5jWnF3/ax4aapxe73xD/Z9RdC2niIoK2IIMpXjX/Rnzq4TeCC0EpVOsvQW
I+eoNjwpZBx755q7bvr2gjv3UzfT30effVbPYSXAshoXpdWEQCz5Zx0z10ojVq2fFeEoz6a/VSv9
6VJzyGZ9kHtAs0AIQghFYV/xyh8oKQOYn2lGHJfdtqdG/949dhJaiSQpeDQXWPYAIMxgYsBCVbsS
euKh8Aqx13KcZcI6cfYq4DAudYUfsebJJhVxhDqxO23DCxzwP5p9dqhEhEQ2ftyW+v5LDLv9rJY0
8ZyNmSRNyhCSiNLJUTyNjzNJo0vpnH7DcEpGRM2GNhAO3NhJ+zd3NsDAr9Pb1+Ve0XAWKP7XQHaq
+NfYt758jz3r8mbINWWDfXyfit3V+SvH2KM/auELml9r0MtGnrCg46d+uxYOdhmjWOd79dfY755f
U3Lq6eZypyXt4GmArDYR3685OnUlrkfaz4qEKvozRIgfgQep2cNFfqoheEddrkoM1BH19ymgldmp
3vMp7wZsCcGLBekSUa091IuLxjS+wqXGBHtKk8fxBlH5HKkR4gwW4H9nLbHqM1x5ZrxXK7Opyfag
p53hDuqD099clcDYvWpN2YbBxYpt9b1Eg3u7yTAsRLEtOoZiX5/1NpUbOD9O6pklBPQkoarIob3e
773WvYELRHAk0cHV+EuDhUk8MPBczabLwAyq7tUeLBWOnoMs237tAEl2QOzJROoIUoF2F8I6dFHs
IkG4OOzp3TtvSfKCcDzyI3VYcNykZm8KWULxVUtG9okFmzNsE4jL4U2yip16X4Dr8i6ohCvl8/uj
tl20mx1l9UCwnoX0akF5dIYXGkd86F8ukJgQidaHtxrJkNFYI/BYEyjEL1RsHUY7z97t1S6bdzUu
kcsoL0rrW7ZaBOX4sH/6Iq+Yd4Fy9PgE8ulw0LDrQ3YuExUBOE9N2hsK/dKFC4gPWL5Kx3Iysua+
2GtwXH6M6paWf3kVRSxoI+Or79MWPQmMxT0TvVL07tLOEV7pcBx7F0jfT9Vhr6LnQUG9Bz67zLxX
9WDPJ2X8cNm+fl5021dd/5Q33p4MAM68m25V1MkE4fnxbh0LutkshGgFmxdsOwhpYdzQExqjtOWV
frrXGp3zfYeqc+dJXaRCtOgH5lqiKC8yhmxdJBw1/KXCMH9nh8gQSrsQ6/MNj/Krd0behTcF8KUo
m/QkTTkMRPXcbhiWh01Y/PqB8PQWzlMQYsy5lnr3ML5GOC2mIbF/REjAchQuDedqWYTdpGRJ3/4A
fy4kWDSnyM9QTGu4zHtA3LOh+/LmpA5C6TIs7avwLW9n2RtHDrY+V1SR4gUbnkqFCtEtSyEBpuCx
rt2ALOZV0l+VBDF3qU8R8aN4mpLtyQZm5g4pl1rfXJMgz07VRQi0/mzT/5X+e8hNoAIsns2+aHLb
SBFJqdwyOaSgT/FeEkIY5nG0SIEx4tTua/iRs5rWhPIm0hLxecx2QW8phTvfuy++kbgxAGJ/hOhh
eHT29gMPWto3ygKiBwxTUHhQIxs8wDX9LLNXgSOzhLPk/BreEZGsfQOW1nW7pnT2wIP1cRMPxyWJ
09K0lMHTK6UrZTZoHXXYYobM1RnqaBKnxaY0QC28aUVC/yz7UStXMf9ctrScgH2ayPjt7v5mwTHA
adDN/WjJfpVpUEQeKSu6Evz7I7QN7XtGixKo/+KFrn406PFHLgLedd5TFL9rxTfwoA8/SxInRZQb
xff4B2nh0S57sATAv0fCP5kiQCXLxEOn9zycrjkYZ5ZXhd7nnGBjUKSegKSwfPltdg3Rjqtx4gDj
Lef2Hg/Qi3Fimk5Kz7+mRGa4N8ubohYM24fJS7DgJgWuAQw38tFt+/DbdZwZ9RlwWUsq8SGbJvn2
rEhdek1g8Fz7UIqL2TK3L5J/HUMh31jvpcr2eUr1G+3JrcGhQRZz7rxhuDDTFttAjdUVnLKSJDmd
xb4+LklscUtGNHluloqZSDi1ShozcHI0L31ROyt+f7KBaeHzNjE/rZeaz9FjAGWcMOG3ejSOGkws
JG9H+6HWe0M0M/s6fSS2IcV0qqwJqNR5RyWhIkqtNfHqPoH9nOOfkB+wSKtLxvgi7qSvFbRGtGOX
mXZnNXfST3TXCSKr1hY4TUExeMhPbwO56pfS9bvrMoZCVXTXXIYAC/lcahcanwmLvU4H5MmZ+IBd
vXl2skypTWj+pNmjiDfQ0Kz8wI8X3FaTh8U7fHwHquP0Nun7A8lFlJuM/dgBs3zGFY9sxvM1POQ7
OJpjcZSuARQ80jg36BS0O8+AvLkRyb0OM8qUlWsVh3xr6s2vWHaCkS2ISHE9whPiUta/F8Jrq9ng
6gwb6jFX5VJ+SaG3e7+MuU1OtCd0QWTGFTAs4bLni4ucXEGksKzTR8AlEWbUX6eIPyMydqeLyZwM
WStWtSEKCOHf+hVzWeSnjRss+WplGOk4yp8pEkZNDQ/FZK81dOTpfBsw/PaAncNTlhQRaxxQq78+
K/lUfS3zRgP/e1zlzxC6tqwi7E6BGwnu6DRH9475gx8cvb2RxoMZOf0HpR7GXXbFmYXEN9ASk8EA
6F8BitcPVsMldIS+DWDnFYdOSue63oYrNl9baKydTHz+MBURg9fIKWLaJunqFRNTHEX02UY3sSL+
RQC8F99jpU9SCqgROUEDSK3uyx1zSInztB9FzkibUuvq0397VoiljmqMshcRykELwRepRRyvK5aN
X5HoPDHIbi13xbGFjgus1EntYJ6Fn2bzzVhkXfgaQH20qaFRolzNvu8wRiwB55UR+YqP5/7aM2IA
tnFYp4c+UttFJOJvHf+irKuuosXyr3Q3wuyT6KRqoefh888Nfn+NI529jGvSLe2x1PP1hG01JIvW
P5D13WKFNUaOqZqtx5+uA6H1FHhyBVcIxl5J4sY3jkccRe5cDywKyYMTYpYEepMHxJl/t68VwAql
HRz+iWEjZGQ9d67NLEahiSz2SBPCCSrncM4bNu9gkgjnk8zJbQ4FOw/wQwvnxiQfSa44BD2kay35
FPafeHkI9Pg5W3aoPvYKwgfYYp1XdovsBoPxwJaYEOIU6ZtkG/Wh5VGwMgnHWWrESYNEF1UZxgEY
eViNBjoVAjt1UV/2r5L9T2shGl/MVIAbCfNLOCk3ARCNj+Oo4W9gVqSXmloNxtCMs4JWxwPXPPhw
xoA96Qj9tjYU2To4KIrwIp75R+v7XpDQOYs8qYEFstLrRMPOb98lpxPQRk6jUiB+Lv3XNCEV7SoS
1ItayfvFduyks0j2qjQEQFl4ktXKB9WldeHlgpJWLzz8tW4XvE637gpz3JjwMzTFYsGl6xieBf+p
f8mMXsJ43OwsBJvZL0A37LO2izYE8gO1EczOSEtAj3ATeAvPPBAspzYZPOtyLMvIyjoWjNzgFlT6
dxKSIPsBFXI3ClicyNp7n3XyRGpkLM5AFnPkqxzDfWo+ct6ZOKW29g7E/4uoQ6twa571nZH4kP/u
Gsg4iPZfBx5hx8IAN9VHeQExaaUnPP7fY1x/d45qRgZ11B6r9fuFMT46aXyKO8NqaiGbPFBN/gZf
oAqtoNhzgNplmElVY2C5yAb5Lx4cZZlwflHXGKpiS6Mn1ZbfUMBek4xOb8HqygkL2VbB6nFQjyUD
4Gfq3mAbDEcK7juhukLS0A46A4XJLbgzJPtHsVX+FkLCs9VU215qA2aYZZ3qhIxTXJ3z7WpzaocR
/jErro2MpoGP5nVDC+NcHjVljcI+bzrOeUI3RXcPZwfZZI+fjLxAiG261IWkV+h3DkEHTJ59do5h
stXWmoM48pBVH6Fat31gMlogY+15gA5OH3hlyTTEsjZRRgbPNqNDrZA8YtCLhBRsQNcKByshnwMd
8tUUJ2ESgR5Qn0mrvA5EPG+Ej/hzIRIHDKFH5nlyQUx2N2wq+VcZLmi4R653h4HcY37CUSmfog1z
bJFavtTqtrkXXwwVEuuuFvYhQ6B69H9kGkSaYGmjZ59804Ojj5sV5wE1hbKO65u4+cjDQg5vS3Nc
uz71VPkLc7pO+wGW6RZfFO6l1OZQmwRsO2T+xucUONI4uqyba69PMqxzDI3qNuteP2xzepgSpVxv
poZrkmNA1qZw/CGhnbxTxuMVp38gKBGoT0A2T4f5giEl4gYwLzdZtCGMx7CvVbOs9Soc4WmA/x4B
osa1kwaSsbjcaKYeuGmuV9VcGqXqyZskB1GSUyAYOnRB/8rmacR0X73vrEWHdLdAfxf4N20eGI/B
XZrmpmP7Wf1sGMIokU4+if6R0OSRA1FAQhQr2gE65dTcD07ky5ipAFXr2+Q/c/+SsJNbrIXgFnn0
1XQk9BBX67tM59GrYpQ1y6MJ/d2do9QKc80Mnfdlv9V8z2sDnEfEpUbwa36fFcMVRXT1ZHDjQ1VZ
GA2y56tD0igezIcL3nK1d0t5Ptetz+X0MM4FOgGDZPlv0Xq6PR+e6KQC+kpNGswHuO2DdKd0JAuD
7N/lK1EH3ioR8EklUQxAkbt208WBMvEMRLRHl9DDDPiTbQiz4nHkSlrz4vEgMcaMf2BHea+OKxgl
uwzp4CuGeWDvrFXW7l74izf8q0YjcCdjfh3c5UEC0GRPsylS8dCtxJTC94WaqLMiunWkPnWVEJ6o
1g48XtMGFjc7BD4ki0fvfcgkHDhjLEdyfMsLNhmM5W+0d68IyzatptFLiMBX4fNVb9R2B51zprOu
WqrIjeA/80T+qIdt9daYHFsQS07CGYnpULZBreH1+tsuFSQOQCkMKDfw8+ZkASIyYOhQRCom/RC5
yvCI+ov/eD48H/gnm9JxnPhZEBj30KpzGM1veEpePexbdWanuN505v/nWmsIzieV7Ru1KkKVdGu/
aEkKhFYntCZ482qNGAMPZWOGyZcGVTNDgpOO/t4sJmS4UFTHX3Po3Z+1n9odQwVRYUS5EGSJfreU
vnpuyM5gn7TBgTdsIygzsvLgwQxQ+E8FsQJbM91AtVKlohyo9KjhkFU7IDzoxg/4nMK9mX7Bp2qJ
yzwqzJpm2sz9Nw3iG6NnzVk7yMuQALn/5dvWArtMO3af4saxNa8wDRDsv51uUInZ0ZdHfyYaITFJ
INJBu2xmSUEwVqK002ilrlomNEN0WpyQ/p6BKDodMjWr0Od41SwDiGQ9rDFDl//TT3gXv7y9sTLL
di/TgAXsUhFq+yD+prvV+ZexCom6+Httnnix6Dy6ydl3HTaEG6feXDwgXHxhGtrghlvSf7CeE60Y
ECl5vTt3vDZxyg9bhk45oNXUa+IwNr144FGIHMvS7ykOJty6ywngninMFDd7rL3Qy06EBaQN9b+4
BXGJbIHYCfugMFwhNCRps0DwuMPRlvTRmehh7SifaXasarY5RJQ4oPNjTfleiX9bXLyHQ8wkXURO
3DEQZKvUHR3HJOAHKEXGCfk/TMeQ+L0nbZwoLWLQ7HEVIrqUaL3hpbztdPXp57xJ2bB7GEKkv+Mx
JUm6ggbzwzoK3rRi5113FBLcDE+A1UdQrJsbugyUxVwpuaQFSlFTLMQXnRdVXNxAhhD8rHEitmQ0
nIWcK15FbNHzeD426DBTHqT1r06IPTD+KUre1i0tEsa7A5IVsNsixX8+Hipu1L9wmkXsB8HLsZOG
ujxQSBqekv0ivVChEx2+a2qeopegINMLP0rUqS5oD/GacqthVRBcx6T1/7+DfiqVzI/jlsMF1XMa
82nCc8jKcUWgWyaL4wPoU6fbp4eDshuAd39NNp4BQqw7da2rCo1pJUpeKGi/jKVfd9HX58kZxYc0
ZZJXbFFYM/A98Tsf1zo54y0nokjXCjCF96SfREYj6uClP57khQXG4ICQj/MGlVds1YFipdFu38Ty
CT5dGXcBdcFoc1q4BNfyCwQ3iIctnEjbt55Yoo4BSU/ssLCh2N9Dt003ugwhuWyHvDU/cmB3vE91
ZY72OECpQg6XFzAlYAbFRoTrG7dCupNoazerruWW2uQv/pRThRegVz9cD0h/khFDJsEgemEecdKJ
+q3vkDYSrfYew9QugEGCG9k1NTpYPQfrBxX/9IShUgjTyQHOYGSAixD3MmI/kdPgaNA72vWvmOj0
hr7NuDT8Cixfaz57C1drMKBaP0ImNi1bz9sPm2iT+1ExDRZ3i0dRDHqUiPjRk/0Dqy5orzN1WdgD
RWgEdYGajsq2g3AnLDdAIYkgy+GMi9ix0ato4b3zFZ3Sy0zJbmwi9Yy7ytYdvMUgKWqMKll4eULQ
LWH++WXEFNqOGYPX5srNY4uvGJkY39ZOC6KanDsS276vqtYEv9qoHLghnyk1un43GGasCYHGuYNN
l7pywW6osrMwE8QgjcyJ4DmKfqd9wG3Fo3slpFm5Bu6JsUXC3vjuW+tOHVMLNgJ9z7thzxUJXlWF
sc8Yc0mHERAA2caYzGCoJmqgW/NmsLjIg5mPCVuqtUPGtw2cIepMYbL8wond2HgxPWJ4RfikPRQj
3dwlNnLv02ckDyGGMXppXarqFRHFlrioRjpNoZBo8SHSnGlllQG7/n/jb0wHVenAvPpjLZ0adR+Z
WFofWA4pEIT5wAVherJvRRnK6mi11hUed8YWg00uHK3+BC+WL7ZhkGG8sRR+hWbLDI+6A/towKPg
UlVh4sx240RK7R2yTXpgfWBw5aJC8+FotPU7ldlnlRrQUPPpBCAPWRvgNPp6tEKoqxrcgWBexjaR
jEyh5dKTTyF7JE5x3HiFQKWpNg83mXKUbagyMbJLUgAkYEoA3of4gnzDAbLdsIh6CYnIJlqlzx8/
j6C8088P02KWTg5ybIrUNlj0xmIBzKtM1fJsvftnxZl6ZFLBTkQk7G5reZ8OLEk0YMJ39rqVTiHE
27EYutAbTbZai1MevpmPxTBBIsBBBh/QSHSb2FdpdUExejBJUWibooM+XoI76ZfjWBhZM1rabbnn
HaHDl+wSnwSEmSGwwxfqiPZiCCFkWSt3g5ayHHLmvn32Dbk7zYwwa1QTPMIqLLjRMokT/11gbc02
beYO174vwAwsoaWpgfYzHYaFaUiGDlwMAYP40EcqN1HqhqO59vNS3zmrVkNpX+H3T0x+e/5Ra9cI
RQr9gkxFyJy9WQuPquMPueGTeSXXqXSDLiWBDLyxP0Ycvr9Z28ui5lG+OrrSIT6KNHg3K7woP50Y
0TNrvj6ZwnmQ47PARFtbwgyXgT1RJKhXGDUJjEgIFf+xkWLFLhiqrfMuLM0Pz2NEeI85TYySxWql
mEC2KX0bUALUrosa3RZSBfcJw17kj/97sxOpP9CuA0r6iN2kfCM8gyy5KiE633DkYxzqsjd6/4tt
xSpuwPP+y/u4AcaesdchM1ImtXdTdhXA5IpTow56CRgS03hjrnzMsfqtuhpwRfVYWDPlCgRLkh/8
o0am+jBt58eeSRepy2RZjLzpTI4M/P8HLKSOXqFduXbcLriwh34sSl6PRT+bEufH5yQIIo+qGhd5
jeFL3YD/5S4PwGBspo/Tq9uVIJ5qbmx2TKCf83XW5eX0CocLlz2zks53zbZmUtAbQHNSU12uuP31
nXrwTcrYPapzo3q22wFnlFMfQfBApUxEpJiHZHhAElUj8JkcSkhzR8aTpGj8vCQ+8Uoxs2Vg7YcP
2ho0QrD6lbJDOqxFw2QV2IAYzTB6hSc4AP/3IO0l62wMxas9k0fVoEaWDOhn3RKg8342/BkudSrt
FFlZ8gHuQ3z46tXuG1aFT3C7+0owZ8STsFGvRehXrwwttT2MSerAFr/e//PubrNmR0sMBjKbrQ0J
EpkvMJnpdWGyo6TQgJH/n1OLEA3w1Rjp9v12eUT99UPtpgTyA6EVAXM1Qp2UjmSgSwlWCOdI8Oov
9dmcDY4jasiBW3Xg+Ejccq2vuSMXIeFtUPzdkdVb+g+ZE+4t2bHEgvdQsqU1MhRn/XsTwJlhTthD
1Ts/h2vcS2wifboo2MaFeODn1OSCyBzzDtfGYKVg7880nzQFe7feQ/ehqA1Q4z3M/8w/U8CZ2bcR
0NGWKXP2TFrby++E7y8KaXOIN1OnBsbBj7QuzYth/9wIJgRcbWMaSSR3dnZ1Gc0Abj6pL7Hdbeb4
RGLVC8PF0epc6l01Tm3+o9PMhEraiHsUj2Cej17HmFLlH+cb4OxfgvJUjirpJ3hYeYNR+4YD3ogz
8gng+eUkI5scPZj1C6DA7e4V2atsfmD/kValsnAJRKoWHgSfcViszl9a3JvtTHkVzjdFSwvKkH4p
cd2HjHepTTzHag5EFdT2Ta9ni5aDcQAMmnT2sDPCg2F39uKIVesyfmR9MydRIwI1F3qmLUR6O/6P
2A+zzkASgo6tonzRWGBABt5nUeS3p6zoaXgMo5d4VBCTEDGcgXj80UphelOOy4j+xIgjyFLka0b7
tk8fnd1pAHuNc8Nec2B9PV3uhtaQWJmoMV93irWB/YIlffajxgwgDsMEsyx2h70h9kNf2BqZOOGV
VflDv2cjjHjkWYdA67D1AoEpYxTZWm8cpc+w90AEoV0MOZgAaDmzfPv2tg79MsYIAyEYXEUEQMr6
NZpTdZA4934xhMcyjx12I7hgMPSjpMasohcaGL/AZvIleZZ1pI+l5AhkLSODcrK7I5L/lN1U1EIP
lzw91bsAxvB8O8Qz5q+vb3NpuJYmBoRmPGA16x3f4Gzl1Dio0vpxzQ0rEu4xv4BqnxnukaRMHlpB
epIih6KBrpSYUHVaWoauHLHT00CjPvyunVDLkI6X1c8W94G3g47OhtxAG1F+9hyYD3uz+bno70wI
3DNYpxxtzMp6eGhxrrM03Ez0QJ3fBxi2Cemv0RqR1kkhufN55DrXSVsPA6j0DdU79U1cCPeZ19Ml
CUx37+ZW56M41ZxalM5lStheC8JZlgSFzS4GEg4nnk2zYx000qxaYP2af/+wf+rUSf1H/4k8woTQ
T9PZ7E9h503UfZx2wX9xFiI8Gsll10bmTFtCVzA1ElxkSGarhN7ucMXgjgizOPczmC/vZqa4p86p
T09tZlTF+/v8qfXHLftuRzizLw5hpPL4SHNfAWE0wFGCHn22rkD+eER47SGPhIFLlvUtmTVxzvz8
ttEGDrvjO3B9zoM2hKl7FSOtWPiZPB4CHwIMMiSKZExYnv4x2pOajAFtNEtqUvN8Ivo7Xs9erCNL
g5qasYHqEI4Wq5nJgNHHB9nt5Vmvr9BM4f+V/eobJszTfQURZRMebZ4PZsVRLqb2mRdXkQ/4l1DN
AiSCJbB4B0SeOWAdFESZ3DQNRWiBetSKQDI5fX6grLJg6dovnNCSAOp20Hr1PbjQ5FEouDPMTFhC
3P+o0K/4dg3TCy4gDCkyu12egBEqsOwqR0RkeJVFT5zTwjJs5svtk7irpp0ZfJ5hPBLVNDqwhBJp
jkejthc3tK6oqj/kKIbVmv/czOtiONoxNcIS7xUpQE13ewQvhjcuHHed6TbJGrizZQQ44bIESxcS
2D7G7wuJwSjwhkHgL3WX6NBy2wmySyQUprwvM9e2KrW40kDWwJ4LsOewtj+tXV7Kh0s5T9nuIcmE
R8NgSIpylGkWJV+JzxHAIeHZ1jXdtLQYTqJan1o/IcbWA1Q4pNBcTwA6h7emvKlp2UMl1qz9NZkS
R5hoj+Kp8chenCEGnTXZxZcvdz5wDb/wF9Hho0ddfA1R94fQXkM4rF0FiZwedLBaMyjcBP7Tt3uv
Qf53LExB/8wmcIa2F71lnlhIqdtFa0t0ggqSH6PcCXpL99ufqj451hX2NtngdSkqNgcMupINp56X
tf1SgZyWTAIR581q7WPU7UECAa9gxelOat42GkuDoiv1S1yHxvYAtZIi/Doi34KPiA6Qp+1+1BCT
vaZSgSf2iY6jw9aKn+sSoqXNdtHNtV150sjUxmEPn4r/8bSWe4Gjy4QtIq75pNwIxXTKBjOGf7lo
RNK+DwFnnTzLeM46dZ46exg6g3anM66S/AaWs9P9ULJ0FYj/1jRIQoxvAlkJdDljVjamylRHUY8o
rgCir0aUOSRzolK+5BbunW7ShI6G4780kHU6ZbLAeZP1dms12V0VIgqTz1JPrhuZRme2qUESYoLJ
wHfZsoklVSuwEjC6db7vQDKjQf2QZ/xwCI28YLyXuc5LbCTcgbJO/artkFgxIdcXtMelpcYOlxjd
TrhrT66kYpe+vjzIqsnFm4NCLqbXNL3ZfSoafoVjj9SDsDoSjDkmUjcpPWiz+hy3PkfjbIrrwz8+
P45YvevTfgOcmjoP/DfLE+Ul4GSu90ovAk1YcNIm+NgPg5QkYJidrbp0krj6C06Iyi9roesObgKk
mtrU/NlEKL9LVMZKzsJpp6LYFozKxm82F1enHYykCIGNZgTbY9PdsJEtA9nNZ3LWfFCd6Qp1aBl3
kt1b6G9wjAmkNxK2ux4+GocKrVnwJfZjoaPcO9TARhRaQX9+Z7CogkC3nH5LgBESnrysEDMbxjYz
bbd+T4QemQ+cxatCCdVtvnAjKq5hikM559OVXggppNRjuUmTO98mg7v4bEM5UFkGGC72U9Lh0yuY
JZp58Gzud3hJKDX5gFZICA+GrZ3PfAXLl6re2t/62WOWigtX+MbWWEwCB54QXFgq6NJaS0XbuXS/
UIAG5SU3UXxxVxrnpUYVVrz4iVpVTvB7o1GeEqFzywyDdWtqu3zl16/hHsZkJpHswKkbkM3bKNW7
btarBc5xNgw78yNw77/bqT4m8GsoGNF0SIdNUEjICVZOrOqr/9RCXs66R8jj9FyKhdFxRR5EeXRT
+iWQDh3FfXmIN9OhIA8O4SPMkOf9UWQ85nrxgjbxqFVKjetehcGFZddFJw9S16eFnMBBjGqi0JoR
HMNYE58uYzPXveTHXXmHudAAdtyIvtvpJieNjPgIgVWsLJDj/3BrM3ClgJuLJPaJyy8/b7BBihTq
STi58+iMY0FTrOW3uTV9gnXRRRY9zY1SA5tq+0r/PP4OGnzJhGV/KCNofMTuaELZuatsUxQ2zBaM
yB+KlOpwui+2UiKUWFnqMKk+reOVpAeJK2NgSOQdMoO7y9yGWQcGB2f4bfB+q8492b6CWiKPJ6Ae
bEFqOorvYXXM6kPGaROm7DfDg6ITyd7GNSPjEMFBKiQsipFLK+bcVX97XmL9ZqBBGlJFTRhImcGs
5N4QnhbBcgYtYEfPrr9KkNXwTsl+TQVt14zjrIs+ey4aVvF/ZY6akBjUOH5GdfpDZupVdQ0tW0pC
sctOooYZ485TnZ0R7/zM5kd1w4727jEWTShpm2WG7w16RAzQmMSlxcZ2Rr6s2qQOFTSNSrB1CIyr
hsxUeuMAXEm2EzkDIM+hYuJNaM+RObMnkg4J28FyvNwTMLOd6YbsoZCVlBVFPz3IL5LpCXCKyMM1
AOYxb18jqPeIqI/cVdyJN064Jp/jgmYdKuDzhqw6tl5e5+IQOr6emx0y5N4ZhhAVzjdE+w2/18IH
lZjHc2NxVKN2K52OW5HrwegkpxBHy7CSM6cb63Z0g03HXEWbKwa2paWMG1mlNsOzAlz1ZfNeXmew
rQt+iDZMBwVLwc65uVT+dqBXJSxNIoGrZqIfxaqb5JPj/Tx3Omxoa8gX5DAUoCL5l0S2Id6Urh9b
Cgl+5QKUqNYulgzHWlsX1/Wt+3ct2oihC1urq91jkkVt5YSRSK4kI5cB1Ex/RKVkXZw11tOCkVZD
/Vne9+TGSiZcFkch2NVgQiH8DFqy7hTRBEtS6SraMDb/JaOOtO7cB6x9yYjtH9L/oLynVdEwnHm+
EbeRfUlvmV8WB+T4YeKyPIU9eL9uRtrMNCxacYE8XXV9n/MiPyxdivZlmTfOGErVmrdbD82oGtz+
lm9Pzr48oFOVLi/1ZNKmpGSnIMwbg2GkzJ8vof7YGDg2KctNw5zrZ6smP32wvr22cJOGXcmidaDG
xPyNMuUPvCu9SyqdbxIJaAYrnpMajWGFDJRJ74VoVjzgyAtDNmnp4YVWOtxY837SBNLKbFMNlO7F
4RzuJtxJgSaHqlvAvAWVJ2pu4jJEf+TULy6eK289Lyf4Ingf18CgiV09LmuwPjWzojx/EKT+/4UY
RmBSRgHvwpitXRm/SQr5hI9btP98uY1FNXcYbMRL0Bd2JQIzxtTKuWsSlrjal+TwGlDASVKi2t9D
U509ROXVbmjLYZXluZ5eL8Gm1B5SsglAEB4MbyBwprKWPYrw/MXIKHTzuAQpf2FCePXbvgzxfrCH
SwdjClmyYjtyQC5j3xxwpMgHRrFG+9yrcInTw54fwb1z2LdxZYzdXOgKi8ahL24UZpoFH4Zlv3DT
fJ37P9NOOC16GUGms/3BL0+j33lRqviD1KfiqdcnulqHgJBZBRlroLG/9MbzQXavGpoA9nrMvsIO
r7uRPyoSS6n4EROzq3yhxdaZfiA5/k20W1tRyLC5Fjuct8fUbQGp9YqAO+/ckUv6n/ZT2v/qvyap
ax6cCYmrqUNUZn1RHanS0vy7bV7l8a5loHh+/FDnplUCVUKeM3wOrBoOjLOntLEPKdYVxGujbycl
7Ja4YRsvgEQO7utwOUGI9OaWbvSNMKiirioVM4awz8AvBZbLZZZ/WasJF2EC0TzpMNzWtbfzv/Yf
Hhyc8KpyNUFh1oQ9kP6YpUvEAATjByFdxBQ9pYaAL++Fg3CffkeXeSP+U7HwAh7HP1+8CnS1ERwg
N8zqiQhaXdQAYs7k16/4qDYdGs773RD+ncApX40UmqTiqQVjsq7ynxwENMklZSMy+/UZVM1Oh9cQ
M8SFamzsIQ5SheOMye01sKgXDcOrrczzGP6d6J+1/grJ+WUNKZKjVQGef+ZmR4KAq1nxtF2OK2Uu
UhacpVtTpjQnQn3giNqdPACGFO91cWZEetGCZPo6jdPnsmwPgWPafOBygKtqm45U0gIz5wtRf8Ni
RLzxDkb9pTslbDCWjECRku/+JNCeu3sJtbW+YlyZ+Yg3PMdu1XrwfehTyLcpUyWQGTWJqSfLnNeq
6zpegWst2YEyNo56qeKWtA0pYCGJJPWBI+xELgy22iip9OGXp1gH6PCYHAHdT9XYktW2ypjeWNGd
WB+LriqEMuJe0YF1EuPRGqFhbAC8UtXIpJkzuzYR165qnInC+pGzON5+IdC0vXiOxghUZFTZEwyM
f0yZ5th/JU6XSrE0MZ9RcG/MuyDlseGqcDPHolspLALvlKgKXzOKPj50F6Wc3INBXg3u45HoKa8m
0FRnd0RFb4LFgSAsdlkLfFOyzcOzVkkUkqiSGqqpJ/BAai59hdJpQcDa96uhm5iY+zk12gmDWSqm
dTcahp3duFTq5yUdsBgcLkZYQ2kfZV7A2SMzwh0rqhVx9lUigfQrMD87tyOh6z5ZJAZuWDrI+LVA
/nOSt76XwG0PI+/qKOliddj8qa6GnHA9Vsm5DvjhiM0qZ0nOBBeVTdzeTMtNTfXPqpgMySY1ayMs
ncs++jAKNOgonPs+5HwfVcL7d4c8htTxFNxYFG84N7jLVrFSHRsQ4eAE+a0JFNVneaTJeWPEIl/G
XzjyxNR6L48kINNmNgOHLrmwkv5B38PxLFLfXLQEMcBlhKYSbJOaUfnHggi5w4UGMkEV0ztpUcvN
j7kN5LWyewijRo5/3mRS3Tbf4mtiLTqutJufxOF16v877fTt0VUqFyRV64JOAyFAaeJirC6unLqE
4T/c2k4T5O+y7ffiCw3ceERoZyjtYuCCSszuabOOpSE07nKGBIGLvgfbbWvW9A5y9kdYHst5mlt1
wWLaFxDI1a+GFAJ0yLtDLN3TVfHJH1WXopRcUssaXOKHxIylKIdGQYb0Wln9gEw/nOGDRCs2N8D0
sSYKXtbnd8PidC9A74ixVHWpCHoEpTMAH+pD2VD+KeMKQcRYl+GpknMmYylEDyZE6McCYE+k4pWO
V67XMtZDu3dKwVsGadlUCluWBF44fq25r/SKoH0DR0/12Uk8pGlrxe+DOaeU6EwltncKcp6EXiZf
9pJjbJqbfsk+fk3kSk6PR/OOqyNrbqoXYNUlYTGJFE1RHy483Rci39GLnFr6rOcLn9lB/dSuVJWc
7IQVMQXWCnutZsG5IAYMBI7rLxtkekWx2VfQgdMW1xF9NfCerWQIIXcHOacd1nh8KKlCcL1NN0lr
c2m1TnaXUi8gwypW5pWo7+rqqNCc7yhX23j8jL6zg3oUcP1Atrj1bvKKr/ZQjm5lS5myarJt1ZbZ
RUSVj5RcaXsHE3YeHxnc5p0o9RkJMi1VZbCsbO0TlEtO2m6BQVN7IfJf5kWOOiGvBlrH9KNKBubH
aKNHPZD9BxkoWARdTXJBinjojpQTmw7hmt9ThiznKxdICt5lvFCs23zwBM64jMvE1HW8m6zvfunq
QX1qYXHsw3rgZJC2LrQcIaXYDD8gwCY1QPiYbVJPAZ5DWh9FmtLUltF/+Tpqb9ktjzmYfNBzxAJw
MMRjT0FXBYM8hK5agLHYhevR+bDv1Bjh9lOeMAQsOCbiVjz/fiQ4eLd+giNbDqZIpdOJ3ikUEKkX
KxPQahyB23dkE50X24TGBz3G0glMgpHakRVLcuOnlOVKvN0LwFbfg4PFOABNRYgrVQ60ZYe9Rxwv
Pzc6dzrsIyej7bQZBJY39tP431jX/22JSTreGeFcu1xgsjY+9DH1DxYhfh3Nh6l/IeYJxdHv4PyH
sYADtQ2XKt/ohI7tNmJhlXGbq4sfeIopazygMa+9HQ8l+SElZyVIC2jRXci/+pX8pTfCK0gDXfpq
i+CeYMkSioxdJpkHyFwKYuGKMZtBGbE+HAXbjR7qToOvpe+XBnskzVp3QoQcMLfPKj4qQfo+c/gt
UwrDEJUuz5FB+tPu5tAAoVxEEBwYTZRZMsAywvnZLLV8c3vKSzTWDLVi4oWj2h720ZVVG7doPJol
z3Bbk2e127uoXBHGZ1v+eKlQrQNv55oq+ViDh939cK37/2k5+HfL1L1wDI4PJ6943R2BkYJe9KDU
Y27ZCK2dah6nDBrsBYJuCMEBMT2WR6iYG54Joo2xDvAbaz0T/T3ny2WeYWf8yTdeOvFM2AanwCaz
ePw/a3tJJYhBUCG9agiLC38qo9n/rKLyVIuKFgcrLO+E9ZyrLMpLEw6NPZoXO+4zBnK9MDV8niq0
xUMlJVNfKhBtVICzIjnhh3gFZEFk/EhOsbGEvL3Dw3wy6T7RD6KN3tJ0BhIEM4aWcQBDPISC2tOP
eclTyTLQJAIJvqnrNpQ6yQTVthMC9qgWmI2nAfmo0uImFQN8/NdrWbX0eyVN/SB4W6fTh1CAT+EU
UTHd6YjO5Tp/Qt1RR/NWbdSDFtFwgaON4ACQEYcuRkPSDLEmfLiR8EXFszDKtYgmvJ+fGrIzwjpM
Mh+kGSfcRzu/SxU4Mo0gzzNZdspEv8c8OoySe/WGozkzNl8ilM1xvXQ3D3MGkMk2H96t8kp8cO66
Wd4V6PLIQjeStMeL/K+X7mkLRu5tWp2xwqh44lln9EA6vDeuFZxeZDOPMQjKVOejQp5ixeNU3DBX
J58F+AQMndbg+ytB71/J++PqgvbrgXR8sMkcuWjkKhfEeJCCT4oczZBC/Y3dHKUZ+27vSXeTUtjd
FI53lxU36nqo8dzdW0yxekYN33R/+og1+nnck9j7ZsLlIcAw8J+Z9CEPmDktUd4N1HxXxb6q+MpI
lO3R7XtkwQlM/n0fl2rEYIZFwqh0x6dREqL1rrZCvUL1DxSMtf04ZDGtlRLWq2vFh0Cb9qAa1fRI
nElYb4uGXnQkxaqGPH1qGB4xgDr5IDj+0LfkA8BszlAUlrKEJdyoJcaMxTfkbPGJKoR77zsCTnCn
jtk8YboznubArT+tbGMsaM2mHgr51wHJrCrznXpnAHxROsgfT3CkE3aoXZswy/Y4GZEfoLk0QQKb
HWuBYuL0uZDBdLYy/2ISeSo/ZBlV3STAMvmDAyOAAJtCXk0T9VlvvwWy2NhxcvvFQ4ceiBJ+pxEM
tnggOaOoUjngAK07PgaLBEZPoKhIpDTu1MrqbFVZTEQP/ph6pfXwPYZAIDmIQtFGWgStt693shnu
SP+M7+YM9GsgVmVAU9QfqtiLzOgGE8dHXHmcLJm+gtrrS4pUfFazrUw05NOkoZm/rI7p67/ekPI8
ghHyCpRBlhRa0rFYXkCHiIbk+lk632BsWQH+EAFNPsFGhnHM6EI1Vf5YSy3WCD5PTt7jqWbJkGF3
e0Y+P2MoYqhhyT32/aW4/G0Dkf0pgftW4nqFd5mDxkoCiJOU6Dh7acyHxxuizxlTCop6vX33oBmM
wl49iCcpN4O+cRBPfKhRlpNvtk2qfNzPSk/9NKEkoBdYzi7DBxLg7glh672lyeC1Tt8vQOnPWa4W
UIOGhsqkyM7Jied0iyDriNudrnoYxgRc/i4Y6+EDCNdyXW/9L9dG1JepM8pJ38oAFruUPhnmiHbB
5vyZ6bxDi5WI5PgXNRwSX1Y3fKdsi27i8BI8w9QFQSywHIn/I6QqlFlqUXehUERsa3Fw/b6Gx05Y
rP/lHc9NiSDUgcLYVXJABeZHH0p/sFnBXR+RufpyuBmI+Dgv+KJtE24LbN0a8RYIMrqwhNFWPrSz
r1BfhPCYt6qxH43W2/rRennuh5WDtAQNN9xIaMrZSSVSwTaOJFInyE/UhhO9rYVYiI7dhSYmg5DF
H5Rw/1ARJT86W+Vq6Ol0mNyvXb8+XEsOFPq5FwIls4OGy2pRm2P3T1CwcS3z/8VVGMH94tB8d/Lk
atFH7ST5zz6QT80XokVSlgVlBgMu9WGxggFQYbp2U5BsoaJ5rAGM6mcajGZHZWh6vAbRrvGWM2uu
zlzYesdxcAnISSxqXJpp5MDCBZMRhcE0d2dLjah6TJNcHphfbHPWh86XKB9xFEROl3Zhj9i/Hy0q
8MmwVm1rPv7ludroBmXLbbxYs9AH5cIzqJhTkk4IkwOHRbaqVrNDph6SSH/j8cUfPvfDLJad2Usw
cHBjSemAZP4dy03Qpg5uzqMz/+pUjneQIzo8RhyBTwmFPGwfv5uv/osE2sSwOk6Ial+cEm/17zqA
6MDOhMK1EfnUF83esYZ1ml6MmPSRp2Y1inMV7dH9+rQqg7xjatuDZZkdyWk95Gru/dVlwQWeyJUl
/wUyPB5Fpfd3IGQ3koYFACm4eW3mHvnTHGPx1HsV2Qrhijy9RWkrZxtCFiBKCCuLOGB0kfwdy+25
T8U87vDBPJTBIBq+24xn/hsXnvl9Ey9+Zan6TgHe8BvxfuV5E6yzF2zFcUNBgSLSsOFWoV5gtRuk
H4+syXN+EdXO9LxCfwwy+ZIV3BFXZzCneGr2Oi9FqkixBP2R2AeNkcXd16PG9XSTtlQeW3fDYKMj
Qd+K4A4jt0k2g8vuC+GxmcKoaHxEFlZNgbWfTMhelGNnEhPLAKOEZYaKRTgwy7VFSZKaxJ1TTT8L
XioHObGkT6xrJtzBSHDuJvuvLgfdiliqmEX2Mr4G8aol7ld3FPIRNzBpzxhVIw9PHyTn3GcNYxeb
xax7aRpkJdEG1nAAhfSdc8ANa8wpHJb9LsYZGtmEvt3adGPCMS33YnUUJBrZ0/dwFvULUPd3VuC9
V8EPg0QSdO9GMBovqokMru1E+yc+YCvyXe0woLEiGOFsQMuxtzEkn2JPZ7TOwa55H/7CmNLvRf0F
gbZFUmdjqvrUpwDKYLBAtq2VVLIw/N9A79vuibyjBTKoVG3NaswFgq4JBEykf0chaf3zzCi48XXt
63ZRoJDyvLtuE/gmVNHeB/2kwlEgJlUbQPfplYS/bDsrJt1D7OkJtgEJKm2kRo3qr9VnGuwfxqmr
+u7dEI34LuaMETitq2RbCEm/3/Aoqa+cNrgh/kTccq2kX2X5woFI3JxcIfWfiytyml9+N/9BxTGI
8PU1axc1L9rE+6N6GpLSlXnsMxSjfON95FdCZ1VaEF3VbPhhpMZUBaRNkefMuyqk846RCdwGiNrS
ph873DPbiPa9FHj2VaoLNjQDtFdVPq4pcNru8InJFSfAyFnzjuNQ5nTSzG9kohtYntGgQ0Q98EED
Y+zZQJ1UU6MkbDkxmLZIx4hb3gc527HlAbkIiNRBhLEjXR4BxPSFYITmmZ+qfEvUxCMD/4GMRW7G
NJ563eLUT4F+rpFQIkMwaHE2rKCe/o6NgdxFWgQv2tzIzzoi1XsvLRamEVp5/LB+yEfhpaftYwkZ
bqlErJdogNKgayGdwAQHQdIVh0hQ4utdaoSyKRA5B4lzRcduF3fJItgfSjXoDTwYw77h2tcSHhHa
lRsHJmEYFq6mdXyqhqNxfHjHlR1Mr+SMDvRy4agCN/HaG97fpjyUNZqHK0gX+44f6h5v3w2qVKid
QPUkcpbtEVleaBEClCM5B37pklq7vSfi00MO0NKYwAR7i8q3as8/2QKl/+rnI8sZzl47u4b3mXr8
8f+TzHJ/OtVl0Ak6kT2J4v4CBahacG7B3xg26OQGL3tQ6bHTiLKEujlQi7dA3vCvFXITVfu5iKlV
fPYwkwjMwf3PffgryrK4lGZMOXs+DLU3evzbZFSOorCcdfiBG4psmVMKHz+NpsfP2wOlFI6ccOKO
YaDOkI1aVd+9m3bi9BjWfOU/E/oskIqskCfhuzOmMilA/9QYRZbCHpaR+qoyp6roJBLm8RTHU/Ux
TAPt2ODJ8uaroVD3opSYQ/iNYSGasaBX3eUQp4Rbz60BZ7KCHsWIv2VGNw3t2nG3fErfbbopKct0
IbMSrP6iuJu1hoCChhlyJC2xrZem/vSAQZqGAMayLmgKTdmA6JUhpW7symc6t4EiAU6+pNIT8GfC
HxVWM+blpFoHWM7/sOEYAjgquDVw8c25K8ctiS3RNiBmDSo3GImVq0NHCFnOd1dObxBbrpLHAqmy
4PfeHoq/rerpHHk3zr018kCzm1OsFU2cjtWyHvXTZo6Noy9T2rCSUvaComS36C8ECsDdk39+PjWj
535pCYWqaFQkRwos2PHuVwiB/UUUnhrZ8C64t7NHOjJn1nGqbS2rzLXc2ZOiGVwmlg+P3oINBrwp
aOkvRYiyYKvJ2/vXMULhfa8FU92AuWiTEiSzS9GyPul5JWYVr8/N5ki0JyLT/Smqa3BK542eYH8a
5IorGZVCv/EZgAYga3pTnNLKslFzHV/9wdVNC5newQcEZUuOPgMOIaDVIc8JrOl++d3U8BaO8XWV
TNB+0/14/LiyWguV7KD8d0O8WyMuMgCaK0AEQZ8EyBiD6zofRl4mmycIDM26s5+KUQ7AEU682UUV
jlom50IHqn0WjvxStL+dVTbtnbPIeLzO+UKnSrqPZhRLm5SEBQN535shNSgiNanZHJJjNRNkEC2y
gjlgEVwL2jjxr2bvOyQKxaYxKiTiRESTAOaxlfAmmOFB5uAAIex+7JzUT50vQzSQZcx38OWuXSXP
uZEr3LY21Nc/Moq0YN2wCqzJJAhGWfY2PHlip96XQqRZYuZdmY9FcHsUD/bqRtQ+VVxH/55rS7ke
V3nqY7rRDdBaxoOthWkDkT1i9Djk8N63H4+/M87v6TRvnrpW1x19/IchIlpepr6YdrANWxBF3Zp+
h64kWwDMMj+U4jdd2RU3J/LWebYuc/mr7Oi1u4sMISX5KxWG0zDztlV8qZWLp10uRiulc9tC/fol
PUuvO1XpztWzMwzTPhi/ZjZHr7spnhYknpW5bujhDZULq0NvhtsMM18Sp7sqhO6UJ8qKbVstJZwH
G/8Og/f1Z/kJZTWoF6G2twJjaflfDvqLoKX0ftKjloM0sj9ovtEPvedSVOvC+JusBHcqslQ25KOF
h7xMWYt5cPQhB5r1SZb/8HPnNnumLvonTLl/ftczWiYob7RM26Rt1PjFKnQjj5FdOetbhPh3NGQ9
pmOnhFuCzRGidpg0rcgNcyMK5rY4zbdU95O32YRxTHaTb894zMnSN1RRc1HnaKGmTObnXCZbzbeu
tBJrlsCpgl2H1CtCrzzLWTplAZ/9mOy64t5qIZ2vtlwtO1zaEdDW2fsU0dcIPVr4909pSOcfXVkb
/ZhplvENcCyVfAXSo55OAAx89VKe5squH6hVfLO3Ja/ydP9NJLFKrAvzI3Qv3daz0Ls9f5Y4UoF0
4IY7f5vSeKD2sr1Z4PpFypBpSHqFlmxPggXNWZgD5MZ1Y36CEkJcifN7dGQiMAj3Mw5+RGKib0en
Ai7X1uFlyT+kpopHa5tz83blCm2D/4ogB0ZBdH/wn1qXb1b4xGFlpTzQSXtffukCAGikkIR1bTNU
HaGoBoetq9NFVnAb4a//mz7NBiMcx8HR4nH9Fguh18RfH8yaDqYRIGVgenhdzivRgiKfcOUPVXa9
kjgWjkUf7nGv2RH8UXzfTs8iPmOGAr2XA4gK7ktC5O9LeorPng149e6ZNbCSG1dONuyQSn5yc88E
FuYxSW8BkiU9+h1G2zYdwLJdvmaoF86T96EBrc/TMNMKXY0CHvTaIqPfAYSdOyVG2GRnTkhr0/Q3
HFkvt3XHJFhsxtcYFH6C7jsv8piiu01VPuj8occTJSeFdPTZ6h/aztPG0dB1V1L4bDe73MTnU8Ye
uH9gykqWsxKylL5sz9i7EzaYqjptwIJtmBca8qlsuPIrxHDRlejw8V5/oNFS/ArbfCl2dJVGaYZ0
1SdzVR59lZoIC0RtrqPMrvsCgt7fv/nc0VdyybDWWVBIS5X2SDJKJfZ8tjvm1jZVh9lonzK6OQOD
lHy2FdSpTz4qDzN7J7eLHVlNSGaXt00jXtlf5L7jS1gLXr6n+eIOmw1Jip1Lc9Rx+msuNbMnpKa9
58Y1CBuAD0qX7Ehj7cAtGaB5YPyMXovL9h6QB8ky2WkD2oZ1wYpRLgpROzYoGQIQnsJxrN+1ZHbo
7jCaVB3Ag91MX8PDzpHp8Bspg8kXFJWfqwjqbAKoYBFWuoVsuWlA5BT8CgbYo19m/W80dRquDPrE
rFGkqxjjDIytEsklOYe9tQGEjhpNkboav3FJeSFeDBjpTjZSAPnkrNI5T53X/1Vq9lxdTaLm9GB8
dfzEZ9zvqR05vAWYK+QcHBoJM3inz2cpc6oeh16BKG3z1K/EsdJr+OgXFRcbawdpPgPjE0ktuaQW
34pE7bBKA3+0n7z40+Qg9vNRjarHza7pkG+IZNhgrS1FWIMPlXbie8+LoGk9W5XYW83jtjsgQNxZ
hAcToKsJqgcwwzpa/HSOOw8WdhL6WZWZDQMUQMF/JZhhOJXVCxFrjATuP7bCl0cfyDnHf/NF/+8e
o4PPFJ92hRM4y2uWRrODH3XTumIbpyWMcpRfYgw3JS26cPBpzyTyy+vhxd12NGBBXeNn/PxFvZH/
YuKKVey56h5veC3sbwAhzQCsB9YVg4ikJtAsarwYNbgNwdu5GfeaBbr9xDjzvd9kf8buMoKXBxis
+0UQF74+VdcL0Vp10DQEUVAh3fOp52gZZs6KNheB2Nf1Osm6Q8VbzJVjy+nBouLEj1poLU8VFrW8
vayA2XhZZbyjcWIeyM2ZwRkihZXbLt3GjSYOrXFSa/2x86T172bMsSWzkl1p1alxdCY01nozBlBQ
JpALmjCHE9kxwJcs2DuEOg4UBGfeKFG1AQlx0eGIODZSAPGbv0Cgdfdz+nwbLJpaApssbLgJudr5
uvywt913xoTq55m/TlAA9HzfstUFvsA+n+fzGcNmC6oXO7Q7Elgkpvdb7NtmoFHLPF2jrEUUaqvS
xjR/GRqbIVgnanWkyQZbs6vkXKXMpJGTZWdHe1DpiL/kRVdTX56d7j1FyVfYQI1JdrPVYsGYUnAz
5hcPUN5tfRhHuZJ6TfRLnWaPTo4Oh/IcafoC1EBc3m+R6fbPon7p/88wGLVTNC5yLCFhuDzCIm/G
+k4K+uCA6IMwCgxf+KsmjfjymQXHEbHWBtIwAD/XrEZOZYoct5a6QGSToh2BMyLolBLD4aBIosfN
xdoPsp1534g0DEE/JyNkjvTtPhxECbw5J0PNno91KtTabgYRAu8FJyD/MtQumeC1P1jGBPRlkGtX
Hc96+EFaQZlWbD9ZYJ+oOdlGa+mQKAZWgg/Dn4Q2t4Iy4FDWbZHYrVS1faLlVqDSThi79u1mmYmE
kis8iM8SNHiu32gi5eYDRZdbt6zN1yKATfjNHyPGUJaoAQv/E6iGtTIQrSs9Gun2TlenW73mxb4W
2KeczPu5RVcg+lqqiorxS4MYh2pQZJa/gygw8ciCpM0vml9uPkSbCIcbRGZA1u4aI1nDyOSUmE8N
qmYVJY90guyam3wGXXKIRssbQnCWukS0pEIrjMRtUCGCYpbFuz7phJHn3HdGLua2Sc3gUltIgKxh
Yn91d926OBLC+sIFcZH0iSVXNHhfNT7kbg7BUCyBrOMhTQfDlNHgksjbCqS9ecgPSUTVpBV6YBju
GxupzkqA1DovIVnoPLjE7iUQjvnPaprHAkpbYLWm2rwjrOOEvvjWQg0N1xM+fMJVvBe1uKtMWKDe
lx87xT+fMoYNQrRbs7C5uWo5qeEWYHOXWzIV79PxA9yySfjny+xM/gPRb6ZXN64c9qgmFpnWw4zF
4RSP/1sbMfWUm3qSa1YfT1Mg7yAl899WUvANLo6YpS4aS8B6iC7YaGBVMDZF9SPZZHwSp+G2FMJK
KFTvUk7ON4Ctc8Ktkad6rqlSfKmMx+HBj+eMKeUxMogj/hjbUZf7vH7wrRqbFP7Q0wp0YDehc9U/
SnGFEQxKCUEmBJ9lQuzEqrsKIZ6I54rBYTZ/oz4oopoBu8Z7iBrwZu8BPBML3+3OI/hNMbHQr6Sg
JfaODJVI5FtgoeEvBMlaTjuy/7iVOQkuP+7XbIDIoSpo60QpKtrrPImaSURrOvHSYdAwXSL12p0+
cpvjhEriOptESWNdL6v2Ue9ed7tJ8hVz6GJ6TFvZQp1C00yfeeLG4ZeSM1+Qq9uybSXMSkVQSmhC
d793wwdy+4pGuerm+JrJQ6NBxivTpUWhRe+dD7FQmm7ZsE9MptmrrWIXNFgVe63mCwG4QLO/NR8L
QYM0/V/k1pjhgwuhWFFM1DiUE5VPuQqiRSVGe79Zg0s1IdmrWOJ+1MG5uO8GJTIHxdPb3TE4GNbZ
ENl8okqEY+qcKW2GJp3SxfIh4nZ2pk7/ovVVNczy72zQ0xCddNBoIYWmKkt5LPLl9mkkP6030nPy
kGevePqfTLitAH0zG8qV6+iV7jJz9oZur5Gi6yQ1dcprseBlqdae5pPjK+63eWAmLBEaHiAUsQrz
zqadCN8SjOpWbNjmnw/hzptTn35xq5/IYm9kocbGhigC8iip8lv9woDQd/5NMvAb+WhtpKjZPLyI
klxT+6HXdtZ+WMX0W3N7nYebwh8YBZ2Ra8gxu22o/z56QqJHV3qa2xaGvakUWcqxbVPBADhvmkIx
KwU2wiOK0W5pi2CD75RL2FAPoia7b3z7T8jVL+e74aUJnr2RfFitVYP3AVwcvvpuQSNjChNqs9M8
oigeaEMlui0inE2F977E5nrS8SCqSYt2szk4nOelA7hdoLsgEdGwQ7qYcVFcE3vrSrGp2pblGMU+
WYUruUbC0U2zGRATrDbH75xjq4EWE/VP4vO8aJzAfe/2BXMinHlIyglcgItc/SPZz8EkZ7xco1lu
sh2nw7lKcRnlRYHgF1FS22Uuk4qDjqe3cPsHZ1X6wUVjhVZb07MBEbNI7SAUNHl1QmBIvLQRjF0N
LMtEpz+ZkQ/p8qdYLGjatM31sk3pzsgkJCKsblHX7xPS75O8gngVj30DC7w5ZTdjFCu0mkMoGb7T
ME08dqkAr0bnfE8AS6UCuy3LOtAAQGBnX1KDcsFUQSdqTie16IziluQyqS9kKH8E18onV3er7y9S
MqLh0TZImKAnfOOohUrHsuQTYeJv1Jnr9gf15QFFF3rcPLYjfJJDkAzlDZ+QpTndOkqhs1E2f5JJ
MyAIK4xZG8oAR2FVe8ztCv3PS9TjU4/btEXoJCs8EX9D8Vnhq7fkG96P+Uen6IoNDiCdtZvf1p3J
IXVsWRWDUmN0FPTwpeMhEN29kObCd09RYyllSB8XTiQpW/RsOGlKVZQLkIcObd1JntxNHrSIyyCI
QGiY4Gbcth7ArhHzERnUXAPyJiQcclvS/R0pmKrDBIbC35aEdBk0oSOtXOcHhE2nhx9GsXulzRN0
f72oxcoHRp7fUonbX+xKK2DDhiivAOdvs9ecpbMT4fb88ghKxlaWw2AsQPGTWKkzYSq/EYGIXtZ3
Kh2+CAfAYBbCwqWeVGnOvgFpjs0f9sf6MNq0BOF0X7rQi9q3N7AnAOH+Y5D4Nh0ynU5L3w6WylrJ
r5/60NmcEBrzbJaoxVRhUdmPpyrElFSFQydk94eGttNhvq1tvSHXmtwR5VvUxd6Q3u+rCwNZkMGl
RrmfvAZljW9GWCbCYqZbAjponlGk7DtUUrGNBQXnE0OovcyUcLCqPmzp8rmtqAidWoSwimQITUjA
wd3/MO6veKS6a7gduvbipW+wNzuZHtTRdaIyGo22+Ar6C3LA9f1OjHeLMcqs2GmVFm8K2bmEoJfl
0zWyqKZZ/lRG+9eRb9tlRP30L1mNzWzThymCQwy/04EcqSN4PhNtCYEvDE/SMAHpnB6r/BZPVRMo
zYLeUQXu/jupyXfhTNBZ4JJH8t/BsKAWjFrq5ZtPlemPMSjUPHZccKh/SFXtg12dIXiM1HuUcD+Y
aDTr4V2PjULic20HZJuzsb0EMsp23fpDPS6/z0+HCGLztqpqXj2NIbSS+KyWb0y/mDH9NtCyIDtU
qUZs5d7TH3V3tMzSZURk5nDuf3Fw2x61ENfohVpIiIYn8BVDO9ucc2VvR3Ok5bm4DyU9EvI/IPEn
kvsHm8LJYijd266HSTQkw3CihABIXziBydxdevUAGpv5nI6/UUxhdpVvo+7c8jwMgQBA9zpMZ4Gn
OXqR/YcFCj12dUxizSMmeAjl+ZyE0wSBGwnEwS5jGWDs2n91+q/b0nRM2UZjvQl/QhJpLIRBIHha
K5ip75miztjYZHI5n66jzM8v68VtBgu+TkfWwfeVQlmsDD0MMT+4vtO7Vkara4LHjHP7obs+Fye0
m4tAw/RfghUhRuftKKtq/WpHSe0+LzEUMFfY/wL01T7H8LfjdcNOEHyTAyGRjePMv0/rQcEhqV13
uLoiuFctIFn5k5OA/C5xk/YEHw3hMtxfumgAgV8po+hlB+meMwkE0Q3qm2f2lL27H5oJ+01ajn2v
RjYzVa5TttWxFXPqwLuZqXn5pxM9mKPygYq3hT45bCVgIhgfzkljGoWbkJY2Tg9VnSmaPp29ve34
rAf0ALMPR/m7dVU3bj6MTILtohD2IBepxboak5P/LJpRphSc0CCzjfZEYR1sxpUfbG/ErIuB/bCR
9+Shforvk23XjiX9CfM1rKaPIQc4jK7vVuXluiVu9oX93BYzjA3maTlVbnUYpvgcJnaknJyc34hc
A5ZjGbzQDYweu4X3INod/bt2rCqT/0/aFSHS+5EuOJYB7haWTKwuP2g4pIA/v2wYDDZQzF51nSeC
v3KJUXJgglz1DZzbeM373A2WU59nPtHBY6+3KQ1diOm0u9lgsuwDjiaK4StBSTJ339ZlAvqw3CJq
Mj6qe2HSZnRDLFOUM4B9GcokEkG9nHOenXZwj96xDRDqu4+dvifPw/nJBKZulyQkHALzR4UjGk+q
Us54ErL+Vzv+iUn/IXznY2Kn0jyQE5X4zz4Mtp+vv/DrS2cD+d1D1mlFMyzi7sI/SF6Rp6av1tLg
WBSfuqdoIfi8m22rOmu5uMwQKs1n6LpqdrWt9ZVLjM4vw2rBWM7APL0WIP6o96G6wE3cYvQ7IBZE
2PflhMaypxTs1/tXwbWAGna4UhFhabB4NUShBfCVnhs0p8uXXawjmLAsceOn1aqIoveem0fYWNZ3
psygpvgLgRtodW0di66Oaxc5h2R2j3lnmDMJ4f818o1XJqbrfcDpCPSTwMJIognPutpvDLz10FaJ
MZvxzwMizLe41rClEVFE62AcnzijJhu2RCuCkrLsChxMPGSPwizeAH08Pn9k3iFtW+IGRcj4i5+H
R/cf3WMYTGzn+062vhUrodOMPk+YyT02UDdNOzmq6Jh0y5FvoIEet3UvEEnYh0Ga8Vdfeo6DrhkS
M1Cfn3y4uKD21z19TghVZVGY0CvvyucOpvtEFvVSVZdL//++5m1xkPBCxzkmE6lVOvbfY6eG2fWa
Zo+IYZJLLwizfEWHEXPKtTe7b/yTLAlUwfpK299fEtSUqBuT2zGA/4YsLEIl78iU65ygHPAkNjME
fKjSBfW1/LGfqm1vQr5RY3gWtU/O9BIHvpXEQak5twgnRONHhjKjWvB5K//BxsZUAebpWGzMK7kj
p8l+XSMyRxn2MhWnHEjm5Aca9WwiMzg9JjqkKc8TPI2JxLwjeShamxDINVHm9/i7ZZwNSGaXzMWq
mg8ByqjlowyCN5PusXKvcBbuU7LZlVis8flkJjLlzPGHINEyp6ssLWlnfadhCqPRmZ1IAlZx7PfC
Ukn05dsjRN+ezqjUqtnTPVYYckItjGcEnhCX6rLuZWQYWujGNcJ4FVNvSb07aEBDXu4eBpK7IG5H
mNC7/1wmniLYK2mhK2Nfm+T/ttUKX3+k8gsb4VLqgJIlYVGkeLR0tTxpG1G7s32ooYESHSvU96jF
oljzdewOzZ3i3klHG57OfMBCIK7wu71GQ3zyNqRnI8uMi5bjHU4SolQREzF/dR1aKGAcPlj4GY5z
T1pnGGUU9hA6QvVVofhJ5mAndGwyaaG5e+LeH8qzeJaoZopRaWx+MyGoMQpcUP3eZSztbURNG/yr
CZ9fP3VtPqTYzyCRtratcVaGC0/RILuO7vQ4H3aX+EtI1mWoHCA77DdTGPfgcnMUqYBG4BqbKP/c
H0a/WgbOns8ogRmwnEKjdyXW/kYeTbW2B9PNEREDplpWKET4SOfgMwD4H+JqQ5G/wTZSQyfHqIqM
RGhgXzo93gtP/I0lUjZnQdslDGSfNeMjQFHK5wuyX+67GiB+WW/saj3X8O0HYPNdGUfxuXijqyoD
R+gDA9dmY87Fb6qM/qCz9CByo3VvloY+BLPee9YRwHkuaXtQ/y3OParFKkQu1M748mFauVi4g1Ys
Kl/SHA0VX0wSqfep87CKm0DRzreR4uJKOadyWoFoBkzu6jjO0wzLCifw0u/i+DPo5t1fPBhDLyK5
saZpIyOgjsFMP2m2YKMNzEOgq9b43d3w6Xt822RwHYFQlT4OqSrHM0fRB3BmCdQvJXxuTkWBCSK6
lr7U6rpL8hHPsmALXbNfQuU1/p0wOLGW3eKuRnizjx8RUwCnutH2iR0drjqBv7XUCwOSHhSVZAtH
phYt6gBJWdQdbYwdpIcpIC3aB0ijVaLl/UTqVV3pjcOH4B0BGIHW1Ngn/eHBPLHTkGSI+UTiNyji
cRMDq2oDersc3fNywi15zBjcv7bRIW1VluCdj9/hbF28xaOdEhnOaxfn0TZVoJxxf4RjDL0F5Xs8
LslbWaqwZ1SPWppnv8nH8WCE/wpN7Sue5yWHl67fbJpc1jYyinCtX4PmVscuymHF3MA3i4O7Df2H
9sZYaM838F+qWAcrQr6mSxNSL3y8DvYLD956B4r3Uzvlh69FJDqLHRz5lnV00m2XpX2iyS9kvpjm
0tgNTpNhr483x3gJAVeHxf50LHFut4L/GctFM7HalgNAhC8/pPM5YcBcTeYcBibXuZf9s0A6jA4t
2pmkU1ZpDdLywCnpwy3OktG4qMwi1aVbEXLOnSPTD0r7xuCFQFtj4sA9W/lZdm0P8mp7CFpz9VfT
BHj83bNT+Ze0DyqJ+4d6IL+ImlMBPsXLbuoz9jaIS3AWMeffRj8l8vKfIUmMUyVd9glbakFHMM6a
Ui/Q8f7ijiMdFSklgpkBT95HdcYG8afwdeRVYLrEzVgbX6Pdvmtcxb7mkDPx9f/vEhqtldZ+TeA7
paVoicbTX8INDm/lYbEgqpMoLx4msk4JdFls1q5+iBvwFlOjLiJGkpuQu3CkDKb1bbLgjjOtWJSe
8xx07qZWb4tGbEMrEKptFI6QhFefuavBxAXXVBJhE0U7Ib4VMJUkuxsGGwx1Dn5H5i9x3Qlq8dl1
MxtD+z9+k1MSDYliI9gHaLBCxF/FNO4OOZw4ImRmC08Ala67YgxzG4qxa0rzdOeT+dPi1Fb82Wpz
qfCPJpIvq8YQM1jgvBW2Pcf7cP7vaOrF4pSJZysitMBIVRyHAbXx5lA+I2XTqka+E8ZCqK+GvqJw
5kHqCsr7caVVvZcppymSZNNat6oZnZQSuv6a/lQeJ2N/hahNYpC3LdAhjRXxo3gK9XUcgRmxxTjH
dHkPXOSiQpSwVq4JDNc5KXqPpBQ8sO3qQD2P1NfTWc5VcmZkXQWqa+0wraih50VcL/FC1wvfDxY3
C0PVlhaikEd6Yeb5sFdVO4+JhoBin4uMPtNspqsMCBpmCLtYBGwX52yf0FvE7Y1tIAzE1k/wDHOi
RFT2X/Ycno7p359NktCrH5abbLy2dn6PRvoe8hUQQtaJ5HL3yopGOoMbwsh4bz0P2kQgUK61ltSi
cyuqV+RiwBh7KbAN5kB0Dc5U7HnXDQD11L5gB8b3z7LRgDfYEu8Y/3snntPW3xq+CvA/gqCObFLO
Xtdk6RMUGrSVyWZvoJnIiAzgEVkHX4azm4paq5KgoWnoPigwFaUdHRhkK754uNk+G0Emtw+DdMt8
+xS7//1SmNPG9X4/b02ih/61wkL2AJ5GS+H928wIE48MU3mAlVh9b9d5zX6t/uC2qXPu4bkMcE0D
uBXsnKcjYlpxllq52sAx8i/UBgDTlTJfPmMNDBaDaWyvGZYdc9XKeywEMjXtPlPajOBFUPdHzvCi
bTG1MBJ9AUfMUCv+J53UJYMbWcaLMZg7Jl2kzhb7pkTmjOIcT09QI6j64my4kyqL5WQ9ZecmCu0X
f/ihIb13R8KchfS/gYj958kG9mwmcBXUTHtL85q80BSMRfLuG4HolJ3KCU+Z2cLHxign1UxTqyMH
rvAWv/wjBDTsntc3c4GurYahbaubuCL/AgVbhbzdpq1zIziEB1CPOJiXAxuxSskqveLbmkL0Ez5h
pv/8X7h6swwKTN7yc8QGXoeR8b+tJywPK8pJHUyxWZmgtmeAPwVvBSb5ZPXRPbpd5UIrJRcFAnni
UMnl0WGeKXZ3nExVRqIq6Ewi1y9/+Qu543gnXG9hhvIzCWKv4jEy4qfHlsySdKG4LaoNrM/f7e76
Dz9QFnwc1CGv6zRm4E8M3RHDPBpT2xljHHTt54/vn3OY1R0/mz2yVB1tIKBZgNHLnfpJFrU62Bwh
CBfUjgr+OosLtQ7IDqPs34q+WWi5BXdXzooOC+xFD7HdeUC0QeIi7Hx8NZvs9onFPNeoq7flE9Gf
GBjHU8jh78SHXyo6QT4Aqwa2YvJHHs+Nz/Dvg67TWZQ5IBuNQjQgWI8jfJmFaVSatS0J60pBan4J
mpu756jaJXraMNNGtefguy38yzk+CqjvD6we8TWI2aBHTv9AvzC49nTEASYaz/jTxReihSKFyTfy
HfNTK3+TWku05EYEVhKKXVYRu93lJ81TmpR6pqHggGYok9AKKGhGXUPkCtgD5Xo4bwHs6F/jthwe
nEMowNhFsbzs5hIw+ADvHi12GH7z5Ise3TI/P5NDJlOC8f5X3/MCC9WN0w74SnERbyBkx1BODoEf
SFjR0vdI4Feau+p+NHEcMRmlTiIZtfpLIxjuDelZpL3kENkcO+dutOH9nQxV+b3sa7qqXV08/yPP
JEucqqbsAoFiv4MAgaO3PDFbU7fsKDIm8oDy2w2WeNeZkVu76nyfgZXUdz+8L9uKV05DfEIDXcOS
LwSoQeZ6kOwP9dxNrfYQl5x+LrpwjmhVCVKaWc6DQ7SjhnbHHr6vIWb1RRlm2ArTB/yyV9nWW7sJ
YbGiX/IqEZ9iEKfFhmIfOrkJAwLgVHQCyKOYwhB0NsUGx4sbcG5B6lGKHRNWCim/edEwsgft6Yxj
0b7FV7WVB8JuSKM5CkCSkQJlg5Q44X91gefriaPH2yeNqDjU5QwN7laTXkP3WrOV8O0igbJ/m7+G
pHoT/V9cSMjrolsTK6OBUKQs9LjSxnC0w/OpiidxctnxGmay1cMN6RZy7MMrek+6MFB7WCjqbD+T
zYFc7NlqAWgDH4QLaJy+a1yteYYRhdyoe0fcciFVP5SEsAcv+vk+ToGI8p1Le+q4+jRCe36/2+3x
VJnlXGd8hCpcsX6qyC8OhEnD79DGpcXVNDX9BVmlf8ALPeuVNzHcRrzaGSDFNcI9tL+BApdsmk5Y
lMdhkc5ycCQCr9A2wLLYSLAF34dgCoLP2GkjJyTcqru7POdmq8voMUkzh7FTEYI3OAkWA9ttky2G
IkwZMfBYovDn4Ep1T9BxhJm9ZCnE7l5mrcwNPR6DjwKPxaYK3Q2bqJcZytquYy4bHB7iqVnbRn0a
d6G+91p3s698f4vvCRzhCEbTZeuAJKwopKyLPsBTY1B8COHKXHV+5peyrjnoXiXRmIFMXOknLyW2
m55dKTzV0DbI6LmLL+SX4iqauDZCxzR7xGnO2kvQygjxwOLzxTj42oLG5l8+4Lb+W6F0HeINL8Fn
QAoiz+Wp8Zfz9GFrMOh59q4f8kzLmLaYkeo0iunHMkV2Wh5cFBD4m2hd1lBpVKFgUh+N1prJFqMq
cUfdde6r5D+zez5XIVC0+Hr2KfjJNDv3F8tjErhT5PFZiNKusMU1rrBdpTWgDShMgN90KgwY1kfI
MDBMQ0H3RWz85M6mfIlnAbMMidygSld6UlNQh7cH/uMigQmqcy/E9QxI/oGLw63sIl8uGTDKtJCI
Mf4IegtykNP5Qkr2Mes72dvLnbW1VvKas5SvHlN29iU+/ot3dcFVg1PZz+3KMQDTk75vtWiBrwTj
zUix6W260WNGCwr1lWJc97piFCIeBBZTA0L0FrcayN+kHgzJ8hym1MgG3+rolZqOhb2LaXa6jCFV
L9Dc6g/0XMBPlAltp6SQcy+oGuwTej8TxoniNlWm6w0NBcn6Kn5GRi829K8GNdrj3EeC6HYiMgDG
eAG3QMNH8mfPqdFCGWF6rDMOvcOhdTkLGu2PELrZBx6Z1H4qBiGLSWyj2C6UWBU9mWLQaJRGre8a
vI9+O4/kOK165OQ1Xn4X+WNlElarSwRD1B7qFTxJqtbFZyksKLu2ID2jUb61AmjvD7wiTP4TVbo8
GhFLYWnGwo4AAr6Gs7HhDCAIHMKMRmznhjJlRIVIneIDeMD86Jn0O/hn6J+Mzqv0J8HCCML3D8CB
b5nPVtXQ9Q10UnGrQwpDPLhAnHzM3UL9K6nGmX0J2yGJIrlPTNPyL1wokJjLPbnJYGdXCvarhmEa
KDvJBykHmFWhaEjk7nRiVzExv3YE4e/KnGU50ccLsn/5oITC/Kg6sTagW8ydm1594A8rmFJ43aJM
jgK/jIqi1v66U0Bx8pkXPiZYv1TT+5fuyqezgrkwbhd7KqOnNRJsUJGoPoA06OddePWSY9qlmYop
/FoXXkOwUeEKrYdD9RoR7asXQbqb3APG+9Yvt0rCdyDS3Rt2IY2dp23EdwtSBdMnSAtfn1lGZmYb
7TCfbuOFXfos5oaP9eI2HzP/8WNRQtx/QduyV77FM+lWyAqdsmp9ps9ro17jPw2/jvRrzrVgcjF7
MvieJNVrs6J4zDVuUOEdCgFgia0r5sPjeY+af7hOxV8d6E6BvAin0YMwRCUnK8EbH8AgtsPWJJ4U
WQzSfongJ4+iGuO2fYEJvWVxHEJw7urxQ77904XkzuUBYmKrHxbwjNro7+XPelogbT371A0Od1Pf
bzAtbUedVSxMJIMeQ+m4aZZWo6iqO/safPFQW0Bs7TInOJ8wPM9IC6YEdctBBDXJHfCHqm8RmE/M
rcXnJKpNUnk/MV78MDR8PkuJibeJtFFM6vGl7GmQCV/PdsH1OSPaqgbrKIEMtaWFXEkeGwPGdgxv
iQIydBOnpX5YPDVLLb9fUXLdai67g0vF4CCQOVjZ4ubHBhfTaoDUeHM8EOLgY1bgJBTyaCoK87Aw
oaosz11q5KqJHQ5i8eq8241bgN6xY3fx6g3e2ZLWFfrppN8hSKUJV23fN0L5UXHjEDFwyU7lkplr
yyKvcfYkd3kGBdVm1cuKju7CxEfcBU1TrU1yShxk7fttJBK4A25x5weFH5aqsqceq2DE8zs8R4vl
rRfTJ7vetRNrbOVasKjmRQWK2qs7IVuCGQ04nhvSz78zj0niTn8JeyBGHpWgapkF1EOgxtK/yPqE
l8td3nk6Q+ooXklAdtp8wbmRziCniQsz8m/1IdQKvrJv5+jl+QN/Y0uPPMPTrLUuavQzBUamx3mP
wrVR34LeDIP0HXC6rkDUNwJnLIqxC5JCT747yjDohvZj4WAJW6z0+XkM2Q6r+/FcgrU7CaI1Vkb7
INUwJfNPxVjYmgCpIn/l2Uv8vxHx3ji+xbwVmQSluvSMsff7bKl+N2W00FKBmMK9O8o/qXlJg88y
MmKIAjU0BHPd2G8OcVJM8kMbGN8lv+beu4SGhbU7uK8tOz06tAGLj/hbVz41ZiPzPjIl1XDlTq7+
b1JIKHxPookQp7ULookLhGz9k6hEuySTqYj1e5V7ClT8AYVROtYGCDlrgBwx5Uc+DgY7cTXjTKnq
fQk/6lXUxRKXP1rW3vk0ioIVJdnSjw20Faptq64PQRsfKXXH+wwxNt1QyysolXK4pLh8nABz/gq6
Ay2xk38Bv+39mT3EKh23N/YhZuRtBNQgzq1PKq7Gax/H37SCw1ZY+CTeMju20YXMYXD8zu0JqMAn
ouCvB5HsrGst1uWYz2/JG1aYeNTysIhcWOjjNGh7U6DzSu2etnReJCTDDQPesoeLanS+SOoZK2N3
rf6tkGcJtth3ispEJHQblkJsoU/7kbTlxumLUPDQrTvjQ6fmdRyMxAXiuxeL6AF4e9ZqalCqTLhC
Ud/zLQBVloKtYEI1T+aKAl3z9ZlpyB45/C7uFFCqGPtnJiuL++U+8yTtE9sdokS6ZdPyv0aXJHks
yeykQjLZb0ZqUt8CwYapwsJU87sQyIo/C6lT+ltPQtIH254Rfks+3vjP/7ke1z4LhQajxm0Yh0gr
AqpYq7YIrYVTzJonH7+pqQ09YAOZ54E2+sPSNFtl65rbPT1aB3KQidhILvmoaDl5BtXYY1D/ccEb
xh4MOeSV+gHVap2GxQJZUCeDoftOmN5GbMnyZfmlxSd1QSX6ix2x95lfc8vlYSDYqe/AKB4oAR9k
RZ3U6wkZywIX/0fskZ4nMkHSRMV2eCUsJ5DOmK4/iTEN58AqaZVL1vgd+0KT/uBTpgIjHMspFexR
7dfaM1Yw09jptLqp7c0060MUvDDUgQZXUuyGc1Yjl0y+jFAxJe4+0bu8q9BjJJZefshf0L909Fcc
1llJNxchafXwPr7WdUR5jUU3xYWNCr3zC9RkvtbP3J5F/5+riOTssytHKarogaaVGUv2ifO6RWhj
4Zt6Ob7540aXItSDKrB/ZZ1gcskEAuJHUDC2OmYJJlGLxICjNDbZx2T/MHtHWNGoEMjQKLpXcGti
XjUxrKiuXe8UYZBkEiOQFD6Qmt4/1Yu4POIuUCfDKrbtqiKbp5FV3Ge6ToCuNCanWWKNOAj1avpW
uBvHOUj0Fa+V37UB2TxEgnr5hBlAnSC33ew1lGBQi9e0iDJEWVCwDJOZpTTsjqYcGG6iSQWVJQTv
Bot4PNxVIp7VH3FYLQ7yNF5AIq84LJ0cIxm5gTfckKEFoWjkll3HHJWEpAm/03MFI7bwOjpy2kGY
ym9yxkTg1tber1goJtEYgFM0ATozQoSvAMSHfIP29VR958AFBVD9SWMEBEF3HVvSihhPcfnuMb1M
6DdyaLuob8lAfn3eekoBuChX57kIorHEfC5YE8Ht+iVoaMP+mpOHBXR2phZ5iLgGaOP+EThzrJsw
fB9fzTZAOJMnG4WCEZWgBG4sYAR2/3PM5njuTRx/ZRL1cD+1MQyzWq1J4L+xqbcy/DzPz9yjz5F7
VQCARcItCpV2vP0btz2IBsRDgHZMA9sKd+QLGeHiqaBw9oEDHBtWA+4WGRhs8O2L9TeIG8rIHKR8
Q5NpHpnW0diR+/ryYRk41Gkbcs2Z/WEUIYAZ8YO2jTy/j/Y7uK/Y59uT7zOdwPpt2m1eVmpAA7lT
B4yVcOePZYJHOHfa8EXdpGUPGLUZiJJmRRMnh/lP+r986qbcjfD1zqLNG7lM5ix4bEzFmExeNvLg
S0Cq1bqqer5OH2g833xUMkUqGjt9oq6aJJwQf7cFr5rZ4OGcNy+Lt7h+aETvtTQ+Zkp3GJmqQ8gH
u8QqjK5kDVNKyxhurPN42qeHNyBstFwjoaolOQAPqX0gYrYBnIZF1xTEN+mFhBAHSPoQptlHILKv
bjDzFh92niCfHwwbuWJOIUqSFfTSftjqxJjTdW+R3EXO7HSiaHIfTSG/D6sAix6sF7yygLWQ5Axj
46ZvU5N4D0H4DcXzIhdWmsLltKI/M8Lq9UZjDalsRQkLinAOKRZveIF58BoBY+LQK8N2K3CV2TBB
T8WNRs5Hm5s5RDIwONOXMDj5AoEk3kuFMvrtvJh4Eie/IlpOdKZkptkJ7XmQM+Qhet5MUC6KWUEx
BGf54vvR8jLKJMQkiXe5Re8oE+a0Hv1kBjON8fq9jwO0LLnD7aTM7y3HWEcuoe47rx49KLc6d1gK
Pv7f5mm+TzWnFH+0T822zGsb83wWQBao7U8bTTCOmLqTVegtqBm37LUJvqJtE7J5tGtcmk49Z/98
AU/OjS8Qo1OdH+w/vkxOtLc1PKRjBAZO1CAKwgG9zjAcpKXt+rUXr+dIg0/zWmhw+0+Qhe9GilLc
ZhRGfUEBk0a9P0y5x67OD+GPXJDBelAAHw79s1Vqv8jcymQP6vJe6Cv5dPhjuog4bBdYAoBNZKR2
8RMvBZHcRdc47YIN8pGzjMH9F1b62yx5FbolzAnI76Emzcw9uGo4f2e7JGNKbuL/ohpgXURG9Ltz
tENNnfd/AhPH26BzIo2aoLXeJw3Sk5KDAwLfu2j9Ejy9psT2uybd8vCicGxRANnXscxyxGTfVmqe
ojapsbSLUNsWvR2JITV7EiE+nZknWZ4663hMXe50mDGphJoWuZ9Z9iXKpWOCWEVrJTwbq78bWB2e
Yqd6L7jv+f8JY6jTQ/j4VtRlpdADC+I8Y9CpbSx6mkhdnI6nPaLrjkioMYwxq599utQ59rxrMAMD
fequAnyFBrVC9yqtXfftyvbJjC8rBMKO4EtUS29zLATONC2FF474K8oLKtgcl+HvOg3xl1feBktH
fBj68mbyZ2SeZ74IXFeTUWkVYCdhaK8EabsmuDtdUeYVt2joSgmFegIe857T4AoHfsvz1A3MmXfK
l6rwpuz3XAax+OD+cmTEDK0TwpMHJss4qDGPZ4MX4K6JE1VBLkzVgPAYWplaRVM/v4yFaGdl0Ck2
loTHRvsiGr3uWzllOpmrtGHgVN0ZcIzIx7xW0xWmN3GlgKYENYmpAgFi7TwzILUN7dDumlYeGFH+
ibhktIua87D7UVcSYEE2/k4XMluHQd7/nJEg/2J+D46YYTvW4jtncSohVzcR9f39XbboSifflYLK
JjJr/oAPSjlb8acBdnhlVCItrfaPAGHZLYU6ISP0qSw3N42ydB0oH0qCrDuWI9BuWjUjXkpea0NC
z657alwWuFfqfKpeduN2oNGw0gvVDiGJub6vF2WdSOcq7QpaHVBbqvujuEBdlfb1Zu1cwJzLyxVA
EKJePeKcddov8aezsVy+hmdVYxx35OHp6nGO7nVB/v5ONYK+3OIt8/7h6iNvf4qKpnnmbJiPi+5U
88dQKizhYtlrC2hKL6Ot4FKxEY2SMLN57tNdaLlVjcoQsD4wpyluQV0yVXFDmZWQAgeyOBiF54QA
63CVr0XBgqB1AMGF1Mc9FYnGcZX062A7m7pcp6JYZ5Y5yofcaQ4SGvX19YnoCz10RIZodNMtsO6Q
0zIWuqcF61oeX7ZKLN6eZSQWt4lGGWZru+kxAvo3CHDvk4lr6guF5T9ccbuOkAz2H0vFpyvuUNgp
8DHJEffrZHFRwGtAPZtIkUwyELgUmo6oYQETgwKcufTYcEszr4YjPTvH54LzQebT8Q21Dq+nIzSd
6ohfjQr59pbaEko4DTUQLzkAaNDskPV28gKv0DoJ5YgXpSgNAW3O2Es2cY0mxa6xHodgpwsJw6hZ
HMpXDaCEq8YQWsMOiYFQjcQSUlae5DSeoODLl1CQKQAj2AAEsA8QxERzlM+KD+VOrMcm4YMQmyQr
x7rqy9ifUoHuaisd2RLh+ryZhhFPIhc/coRWweUlWlds5+NatYXhpkVVoEO6bxaDPBSEJOfd9JNd
CSdXUtlYpqreKAjqANHDu1sFZo33QI7DffDWg8tDse9eWx3nvEdXbRyDAqe328cD8e3nZED62eag
8wLX39dSGc2lWZUwdzfp2bDKAnk2Or/HtZYx7G5x3Y/Fg+W2JiOodroBq5HNmJZglRRjKBJ9218j
rqayMfYTGSoOn+HZ897bwTjsAfFO/T9RLZo68beCu3WE+O+CzW5sCUOcS2pfHdoR0ZQl0qCf0be9
H4LrVPrbvFlf3xNX2CAcmchmaYyzh4WCnMOib/CRwow32uNktjC659t51hxOF9GW5PZPaa+McuY6
tjl7sCuqexBpzIQsntEUqBZ7wCctak4pTUGiJbTB+Ygfrote4+cAzOrN/ICqZz6U8gETb+J54A4h
oozG+OgAW1x9Lw05wf32gQVq61XZJPYwKmwrWS8o88bbYNGgM6CLbPOjp2XV7pHYTd7ZkSK6Ue+1
H/NF3FoSv4phJYG6lDpI0DDUnefISjFNmvEcrj31KayjsMV8bqAgU0VRgHW1X/IsDGcY25uOjJwm
5XpX/xNM/Uso18EXaFURyuj/iRQd2A2thrdvY5H5Dg5ZK6lB+RtaD30bukwagW9h69RoBc+9WM2g
mcKK9HCSiK0b6llTEdR81UTG1PIrTXPFuVSXlIQJsd6JrpfkFatbbQeRd3EIdkdBTyCsDXaOAXrN
PBic19t1vAfmZM90e6oMShPkwkSqrZ/3zyXnUEM4cZvZQ2CKVddytkB3zeeV31oS/SlPx5+tXdlz
9qfaE2qgENFtjosxQ67BgPQhx9n/yenlHa/JDqaotNXuwmZDQK1KEU/YUjChi4GOemePh9PaZ57f
fk/JBdAFXHrEuo/oWYUE+U7M3UTBG2R7vwabhR2cBQdp4Ur7U7OGmkNMN3mkiGkU4vqfwE8KSwIs
GOiox7RyVbXge1sHB/YtAfSmhnzNmNAcI4dOYnRonJVSwoyQUwbGxf/Xfy8S6Ncl15n+MaTTP7U0
BoFTSVOFJxwC9mbiUbxuFSupsvylfmLjn6IpfKylK5SBJ+iGpAbQcvGEO6alQjpmEz6dgJX/kfrs
p57KW2NPrJpecBoRJ6P/2Iy+Bp/JEL2dYXvyLVnLvZWIQVkHVYezMYt576nVqLKQaIt3nBthFhun
YVeynS27xG7V20OWJ0yu59CDGXxycmjGsIkawYCPAUFFQAvfYDqe1j0C9mtaCp78DYWiERaVeGLl
bg7P2/iOlX8ziUbfeeJMGuAacpalio1387bzKGNDIU4bPNcX3htegfhl5Lg3d2dukcnWwAVBMdRF
+8zHzrzx9obfWUMGxlOU1KG9v5HJIV/hz5yUIq682+IpbTGt7FRVK5JVIVL6MPtd1pOhAVGR+wNI
OTHyZWNiMA1VVzcc17wXuX+3XXAtqK5c09g1P8dXQsuwjEG7+02by1gtQTJqeuw91vNxRIV+WV+l
kxTqUAEqbHvnyy5TQ9rELUL+cN+qQ9GQahzejnBw3PpqR4Dp6TD9Ey539ENkUtZ3CnIBQNcBQgWX
1NlO8S66ETec+VVf58x4LziRzGPqGySb33V5bBL1Kj3+qlpAs8MC11SUP3MovOftbqfP8JAgpD9D
cqI+2KtPcKTO3X8uev8m+IXoE2p5Er9gjDeR4HeMCtqpVUBAxbDP2LfJk29Pu0/YUDzuIL9HKtDm
KvR9n5TZfDcRvIkOKJVKISwuKDeGVIWxgp/prknylMIIjLgCOA//EvOp/TeNyUzMkPU29ZEXfdv+
O4T8bxiEPX1r7KCWnGibAuVJUE+ebKy0e1Yf8XwjObPMHCuiMo/L01kJ8sdtO/zGuFECIsiUjLt4
fTy+cQq9QC2n8KicsSdgQfpNq95zbh2C8+NCdPPUGotKXu/KxwWVR/ZjVcvjkDPUQgc8J4PQUNII
mm0g7OKC9JrmjzZwMpym1NCEhJrG5JFFmMk1MzRLc3vgAgCuOwO+vvC5Fnj2x2LB2v6vouxhPZZ3
qencVDuC+v3fyml5FHOAXlQwX3V4ZaD8XqYe2GF/CQzO3B9dlyC5DGHNduR13pVSiBNMJ7Wvw2qk
xmq2sYAdJZWbI94i01dJSA/WQ27ND4wGJ7fuBI3cCqjqOCorQBjKvezcMHjB7qOkgMV4O7mi/BmU
LsMnefqmBKKsvF9+D9y0EGLfIsPlfJIMT4vFiJqvyhshrph3/KrsXAx0hv2KprukZMZXYvQ9jlum
VB0GtDMWQeTTEQ42rRh54nv9qx+wb2NFMO/GF71p0nEflMw1c1njjZ25ezZht2gEu9oAV54fEz8X
8vX5JUcUNkMvXfONnBWCSaGDaCG4xIn8Ac5oyCkwEYFs/VssN6NaNA3FZVy38KF3eDVaxHQRE3ig
1ekePoM+30QpnxNKGFl+xouCwOTxSuH8PPP2X4xC38g6BLZNqC5bP9BTQnZra/3E9HcuG/KeaH1+
LwW/PEe/0FTw2iC+o7vTjjXLXD3PSJ/V9wYp63fnXrpZbwobcwal5+MN4lGnRDmwNkxwtoAcXyh4
1/78oI88G08FNIEuOe6zRFZpUFWrZ4VYxNkUOXCUg2/Paq/wWN3x3cVY9SCKK9PYAht72JVfbP/n
R4/r1FS11ty/90QMyOuKaRuIiWyzlA9KOWzfCnZKHdvs0/VL4zdDz1WSUty7dKqXMu0a3JXhKAa1
rtlcBK4SNDm6+7Sw0XSei2oC6WcCezeL2ZrcOeDHkga6yDqgUMLYMewJFfB5DSAYddbdkjXPJCs9
PT4A1HaeArE/WBFyUgU1PXuU+sMBGE+McuDnaEv9o5j9iezlk6SoSPgPoFT2k3o03r4ksqEntUAc
y6Y+pVWL2XF7yp7e48EHdpGW+CGh4ZOJAN3IXWk32Z1UO6WNW38O+s9kCgmqpRSvSKmiwSdpuVeN
ELDKKUx2DhCFTfUqHOapmnRYkN7ZxmvBitEDf4OSvtHfVpM5bmKu9BT0W8/aOnIz1OzNl8U5lskc
K0N82griXbvKWeIHKaSqOElWnNQ0NrHBaAYin5CfK5QotbBI4wcTDMBLZg3hZX0GebZdAqNvXKLt
4ujJdA+rfy3lxWDjLvONtYD1WAETk8lz/UcTKCH1EmGVxUjOPyUIY4ZSW04RplwvTicu6TvJBVe9
TOoZ9Ko/p+Cauq6LFiWI9QEle935cDcxe7gwV9Uo3J9s12aYDcQj49LaPePi97O38Os6Q7LE/HDs
vIJz9EQgBCKC2DC4n69CoPC7Ba5rDLXM+/c517/WGxNBC2iSkgm9YXhgHrhdG7oMRmHKfU8z4Vpv
ouNuY9g9OPcViufFY8Kn/i+q3m5x4j0fh7VDO7hbjMVSEC7kqubmSZHeFTa2dadRTvvulp3c6S6y
KJvT0nuGon0zr9A0lAc/g+tZiVWmgfXsMtc84zyQ3Hc0+VfLMvtEXpRfDbOeq+mjMoBJ0VX+MqQW
dIOomNgirYpO+RxEBSiQczQrcab7FcIZAFDwoZhoxzfwq5IFDZu3UO6Z1Q5m1SI3VaAMHkUYqeVn
cBoe2D25ytIeA7PDSrUAlAur9l/8Aw8SotlDjnGWXkQ/xrVPRFE9HF4aoBmPcAykFAds/x+zTj9K
QwZc7Y4OPSw2D0UkTUX/YYqm3TA4Ht5n2CrHr2l1OKdIK25Ht0GRGYnkaoKvYWsPSy9lys2tRB7W
XcEv+9N7zMncvwBLEMfQDqKcqYJN5/s6ksniuNg+uDOI0WsFmeC29UzmuXpeRSYlK9boDkF+q8y9
UVpy8GAbryRkQoBknfOX3Ote8Rw9/PrTQkpa5uBKI8W8mL9IfFQJRklZWCr0mVrnJZa0hAgqVHyz
tFpcCRRNSJrRWe2Q1oH+iSU6sKuiLuWJSjgfRQYxvQOeyGERGpid421RhAE5CsCG3keH7Ze+NsxU
ARfVwRXWOFY/FjJZRMFAbNNTw7PWNbQEhee3hGmz+iRM740VA7lkaKRNZDqR+4OC+ZNmc/jgS8rY
IDOqnGlR93qvdx3CxpnXuPyV7iB17uATuXRw0eUyjmPAVUKtOIYUXzQFuwV2qHrTEbVsfZaX7/xh
/vPF5fFE5Wockj+cK3E9mnq18Avy7V3TG8KLUe4xw4tW1Fj1Snr5bCPOihnkZUm45PXaofVBSeLD
7eHG9RzWyO0wHxejamBB0gVkdHHkw0ip0XhddcUMjm4JMa1N2PZEJi/M9J+RC96zj6iyP6Q/Oa1s
KdG0VIKJpJNU025Iq0Azqj8Mqeh3J7iUFf9x5O030B2+ahiBfXXLN8jQq3PfyuAYvgdKUQFo4Qex
7tQItbpP0KfIeo9NtTeBhMpyLA/o0lfdgHI9PFYMHXCaWsQqG7L19bTyxznKQbpwSCYQ9Yw/oQ4W
v9Lmjvh+84DGgeMrK5sAd5YMQAE095cpCGqLMG5acr58tT6ZN0lRHzqzvPAEvPsuBCRq4nXn94us
muuj7+UmzGFq8BKouK3+G9k5ewu/JqEIrGuQzuvcGuomriZbie+lq1YOGEVoqBUvRN0RqvR300ix
DuMEMPl2TMCB5AxVCW1HtG7pepsQ2yhCIK6yqprTjDoR5ZbN6mEaibeGH1QWLdPLpO9a1VW5JlHF
ywcqwi5ODekY/k75i0FK++ODKYpVmms6si9ZhTIKdzd4c1gPEUUhZb4vX0aj9kc/U7fosseWxQNQ
TZaF9PJ/QvyQN95KhuXKViX+UCwWhK6N84rbeDspoHSOYfhXiF2ZBNDQPBFKNFRONDXjaw3aYaq4
SIOKXFWV0GCx9qCP7zsvooPtGL1to9REyY4IjiPHczyAzfT99EbUwSyh+Fwyqcold7zBzXtXdbPU
P/voWB3XWgg0SxpEW8DTEwAOq1sre+veI47lI8UZ5aNTcn8IS7xIKwMgoR0XOfaKIv1cdQZYs66h
WveukD5J3MZUeUYbpLQ3kEVzSvlItvPlSNKKJzoFRFihnbSYkTxvb4h0XAa6dOKqJ6x89aLWH3MZ
H6PEsh0m8WK9+zYjrRhJDFot6NadyOMiLkNKIiTepw+8mbJhtMcEKLlGKEF8Z+H1nD0e5Uok1Y5R
ULj59BUa02FhQOiKFSAmVpfMBYUFwcIK6wd4dRZQtECwYcImtMwlicNDg2YIcoyKKCOxme/XMyR/
2dJ7yQDtOM0+TIZyoP9BQsLTa+x9jJ1d9eXYP0d7H+sgcLer2FhQMT/LOcelfX7C6bVkUW97n0uX
VOqlUWDtqn9uDLDagQ5Hkoy/gVpgb8/WwJE5PqRk3+f3Wexpplo6aonytsHZD+iKjEw3Z47a5rtd
xKu2kPxigFsnMzpSrLQRaDbkZs1dxvOGHtBTEMYOERB1gDN3+AQ0T6YzSZzVUf+AYeJIr4KHqmbS
OcmjzcdejlamY4ykJRcDqLH3szY5m5tpZl1/BnjMCOexHIrUkOgCfFuwpjgHcmMJqXQmBQmsTZXD
oharXQMpJg21r94PKUnApo7SoHkAtKo4ld1s/8gIEIRQxUVUOLxgyJR24ex1Os/4q+Jaim3L67vt
1pgz86cQ39XUd3fP8GsdVau0nPCInzQcx3DWFDc576ac3UpJPgxTqLMLzOY8RBw75K8VhLTeyaIr
VOPDSD5JbfANNLoPXPw9NovVUvZR73+ihPn6+NdrC+frvQZM2MLae+4JHw87RPpp07eaEozBWNit
dzgbPlD40omCnu1SPv9Liah/dIxGrIq5KDtsPkCzi4xFidUKGdCXL+qJmYnnfAK6MPAThe9ZIP34
2wO9fqoQtmzQQmCUVyUgXkgynOEqBIlEQqC6GH9xn6GjMNj9RIf+LiPd0s/QNC8meqcN9fZ504N4
bCJVlwS656TpBwHzuNgmikIubp1aaHpVYTtSi9Xm5aW8aqiGrYzoyDcpzTVOVhCY9T652nk40P+0
OCGkJjlVAgzCSnkd2Q7BSJoofLZAf885aBlKBecJVVMtKR0Q+Jjc8d28QNdK0l1SHVj3+09VKKZE
MaotP84IzU1bP1isF3QfgGf9ZvKjzFZHNqu+hKNo6EH0PYxCwYwpZ2G+ofuUhjbqdWhYSJ60t289
h7Jmh6FvsMdoPeMO+aMLqdvlfm0NWP77dXwsdfwrRiJQfFq+qc7KrZ5rjPs1VesUU5pDC37rwSAl
eNwYFGo0qNRPa8r8VN7MSfp73q7Bo9IAb4SjTQjCZUKIyAdi1jZKk0pnZCuC80uNAqH2cOAbdOqW
Ss7/2SwxG0aPCC3krqDHk1PqLorjRrzzVDpr8buAr11NLFy1Ps6a58wJV1rvAHgC4LhySb3gvFpc
uk/SzVWSI17qXtiB5TKNhr1QRkNnfnDDRwcMOOXI/nOPQ1VoamfkndC4rHju6vJyNDocWcM4mhgP
Mf8nf+FsFHpafYKlx28LZgYgcnHO6apPApG2OiWkP39qGa7MTLb1unEKmc8DSIP42YFZ53xgTCwY
8gSvd/Wa7GjFGkrMHmppvYJSUEcyJ5Z3twykljhDq4CzHNRPbBgcDSr5NLbxkrcXd5Ulh+3VbY33
f59mbHMBDJs0VqhJsgSjdoZ4sfqVy2/Aydte9avbTGHMyBWuiML29ZLFw+1Rx8Lh+jFay43v5QFI
sTrZKNAF3k3HbBTc9f76zU2+5N8Wu8KRU4CVk8ytWh5Mqgv5bGqgZoQJOntq17oIOsqycP6uwsuZ
nV2KypdzQr7Z5a91lGNFwpY0Fqwsecl7MJ7vz/ae0kIvId9A6wfprzDv0FWO4A5mp2aaKWseGZeN
wAWcKmsdEOl16VyyYSVQmMBZqFFqtBmMhAJjuzQUTYqBXtUCEEoTDW8RYF16L901S8aIQz3r36Mf
wM75ptRFI0N750jioRLlz8t/iP8c56NaOtfRF6H+/Of6tgZ5lHvrvQoouppbERsmo74iCaqD8qtr
uTqkZsfYrH0EcBYnzDWGi0+bcksYfv4kADVM1SRzip4oCsW8yEnTUSu1UmmMnQdZwTr7YMh+Pw3L
bkXhGyrmbGNaP81HpRyRPBvmVqKgWvmCBXov8KZYss6fWBdf/1Xx+R1hqgeFhB/ZKfa8LWzqCT1p
Odno0dvjqAoMqoMoiQEWTH/9vUUfl5psL/JlBTmDVW8LjHJiF+M56eutTJsBC6TcqcAHqNmtjcwM
qymEw4y34CYj0AKCjihrDvsesw0PXrE7YxHTifm8zi80yCk9cZ838sfsuTWJY7ASeORNkNXCaGVR
oLEOPBM00m5QX0n4+DNIFqwHHR/Dxv3+xMT2ykVUGMWTQRF+hBWeggGq8COQh5nWVNb8HSiku90+
38toedN/aevLM/P8bi4A02RKe/QWx+fVcNaPcLC+UUghVfJtbq3dyO0K9g2nuXes3oVKGjdCaZ6T
HkGojRHYHdJbrds82K8Dv4oD6pk94yN/Ccv+2hRyrIQ7+HNlj1onhqZIecUBtcNG3IZi/kOBoEKn
SQXT0Lz2Ak5PM5P8u1lcJGwdnaIh1aUQVCDOmI0231MYDX1pHTuAIlaTogKSYK33TaWmTqzST/JJ
yDMa4HjwP6JY0akk5fwIi80pDlx9Te7vVwJBc1qnmESyjojx/VFtA+V9h3/QERzLIi9jcdCamLUk
31T3iPEdiukysZEgC6Wn87EGPjYlMjNlVt3xpQw1e7i/1197F00Ua1qfO2+rXyb7bFIfabk8/+b8
Wb4wZfsIHkkWJsAMPKtIqaobiNaVENfEiWCyrP3Wr8oifAkF7eo+kz9cv6MtWteEAsSozszfFEla
jjTPG4yC34e8zYhkixB+VgZVfUWRCuxMGgIup6/7vYK+dMYe57phIAxkQtB7cOUrIaOUUvBONt7o
0lhCHIXHFZu2recyqR7Mz/Q6zRny6Rmcq6U4XxdCr2g+SWq4gMwivoMRUCMYQ8HPhNQcyQGWmqIJ
AeMq6cfQ0SbsKvEwupPl0UkKJOCazKF6RFwpTwtL6Ws8wsENfNx0E2vNePjwsiLKJm9Z9JS7CZ/B
TkJxf4q+Md9tiZGpzUlhsMcwFTf29Hl7li+6ugHFhr4ofH/aVgFVYj5RJke2LmvV6pNgpSls7p0y
lhnNWCwwff84omR4NXMLhpE4PPY3y+tSM8aC35j1EThEetWz7qKEXj28aUsfVhKt/hvJlqbC8iba
cKvDCxj7E7GuPWrpKA9+tX0oJlUS0mL7dAqBvJ8LHxa7geaANSnF8DtQQUSUB3cyfqT4yDV1vJFL
LgFSE9bPMicqR/rOn1PI2ikvlvdxz2yqIkKU3dtg1vif6sxTi6nn/yYjePCKZgICltlsENk/Wfwx
/2UBX4v5EsIZVU5Xa2llAi/onpeCn8h4G5F2hHvZXs/qwqQlTuJhmIqTslGsoG86iHZ6Z6kJdiQz
ga0Egf+Ky5Ut1hCudRMaI2NZeP9UelHuursi49UNGcGYmdDVsxxp2zIbIC4STHpDY9NVrTBr3HR5
BT4jCW7Q+u+shUhyjjYHcjeFkzpLc4KIG1P46E0NkEe5xN3jjWsXj7a8mm9bBCpXYyzfFGh7NTfE
tk4QvsPhQIHmbrvxzmB5zcYtJQdZBUIps0RpM9KbPZ7u1Ezbvki8aWeCW6npBbELa1rB7J2cFYCr
noZ5LhjJyaQrKDDh1VXB4EN9h8wXgt4161mua79JQL0cq/nA002azayzDl4Hcv76Zx1TeyQypx/h
yWM2g5fVYoL2rIX7t3jK0BzmdW9Pyql/ljsE88Z71XnRkAi4/QewSUFcBjYRaNtmnoIkG79HPxsH
CNfiwgB71PNaHupyV7sTO+nQecdZ6P529wmEfOU7jCHpC1Q8jBjKhYST29+xb3FclEsB92xmg1iI
gbKbJjiwiCRDric4b1NMWoRjVsjRA2xs5KIksgwaq0i/BkmJNlcTXgQI2ip3DpRgCLUCTHYjx8rN
GEyhRb8umJk+0eQ8PU4khbgLp5MGe/FJgvpJ6wrHhi6W6u8cc3LlMiGkoKyncrdyAWlgAM04sGoO
joHboQ08o5/FZI8jkl4GDs4Zi9k8JnObZTjcyNZ11N1Scsadb/9yGjaiVw/22ffi86egGKJ/rGmq
o2oYwmcaFHbf9UOS7PRUfoJOa+6jass6q7znumtYYW1YcMlbYt8XfCca3Tsq9G3QRIOO/3cuHbPy
v1MrQ8MB17tngu3XDE3bhz/4bzS87ehnLt3SALhKCOfrmn3LRSjMSxd6UTyY4yoLBvxA9TqP4Tri
hIWhKmUEh0j3USUj6Fous6M5yfPuW5ieZ8Kj2tk0Fhkfsaqq7KViv+CviS1NgY5QyBFMY7DBvaLj
SRfbc5TR1b46on0vo/hRzwvTccQZbfLqP8tR7VkBdF1imPCpjD8bMFt2u70U+IwRn9Dqo0eGjVYJ
4BEmY3LscNm5cjVE9Wc40bxnq7AsBeRJPoMtUw4gmve9x9V0NPy1LAoNC1fDXcemOgFOoVEGCOMK
LjHSkNRsf/QuKg5GcwVwubNIs6OAUaVqhQiQ2Pyq2FEnzi4l5rYLrwWbdEOWMBI1jJmf2mSdQJL2
jE7G0ZPskH39zZpUsEKWa6a1rim6PMJsDIukQmZYQfgJxoBXrdfNhR1hE2m2ETPhIUOiDrS/5JfA
6VZSpXc5qC2rK0CeLl90TeOrleBDdBuxxyz3scsA3CYq/1yQ69H6JdStm8utvLhOpDS6u+0dhAdK
m38GQrIuQmxzMzRtY0KXsIgDoES7awVsZY7o6xbCLSdIenK987UnME5MzL+VMkDhqDOLdJEM5I26
7Psoi1jWdfdQ1q2CXENtrIatbRavp/wH983gfnMjzBkgscATylJ1YDqejPOIFqLAB+tHbHb52mLW
ocLFmWXUrQKZTMn9LTcw6VZpRKIVZJAjTKLk2k+UPyFT8MpyQ0P2Qygm1uKcaxebYI4bDGGhGNhO
GW4FStHIt01d8VYwEkzpZKVI1uARUm87pG4OLkBlvuhkNtnJcLw/L7hlohYrWoNClnv+UbSBCA9P
PeIb5qB5aILgxLJBPWOb3P/y2e9NXILji3ZNtEhw/XGdzw90aYeAgPAtzUcHSRxo9Irk44uA/8+Q
VfCU1BJZOZT2HI5e3ma1Ez0gdWj8NzUQRAYVsPW24/bT/GUh3tKUWk3cU0HRM5KDMDdXLIwJIlXa
poV3LSuQFc4vF87Xo21J7uqpGz9mYkOl7LB6iSpgCh2zkCkJ40ke1J1n3Bv2GDEgeDwkVlSD9wfB
rjAqaPTTBXH9ftQRQvd7irt6D5gaF1P9ueVG/gv2digLINKhtC0dOhV6S1fEN3GWZbQUwghamhNS
l6LJ4OD/KrIYMbOxzTDti+Lv4P+X7hpoRG1irApj4pgbq7wNUd4nQuSUxpRDvatSbt8rGyQ3S+iM
0OKTZIMyv8cMGl6ZAptHmFyGOq9Mkfezkx43/K/pUMfapiUU3iuqghyTpB/19OjOCg0knlyJVxgK
/5OnoAs9z268XfvRsf63yhqtFdNMNI8jTHn1XNJkYbBgNcs+Ba0gOc4k0iHQd1HmuXB/yd0oKFqz
fhRbrRqp7ZWvMLZYtAK7gCABXR4qbm083GdQedC1GbO7YgoshAzyzo6XMm2CjZNizb883EpbQh0N
xhjddE+qDb8SLemhLRpAzWeYH8x2HjvchX/yyrA524DNwLrp4HFgdWa9xICMnTi5Rbo7ersFJaJ5
O1rWf+5fXmLAs5qAoTZtWlRBkVkWLuHdsAUCabNTmXaub4cNJhWAvkPmYQzPH9FpAWKxRgrMsi0e
uh5fCaPh61DD7lV7Vw1yY105izZOxxe2QXLdJxW997tz2k0ZfeABRs2v9LSX42yhQs4WvV8f3WIw
MUY+q10r2Pq5Tp0CZk6Crbq6v11xa/JugJAjFozuKJYkQ9SbZceKqsU3LwFaJuzp3BjaIDr7FwqA
6pHc+L/UtNv/PkER47lW+dRJA+nM8HWgX9WunmvdEjhro6DCKVP85mWBksAqX4q8LD0BC6kgiouv
RzWU0R46M3qGjDctpckMR05viVOGz3vlB9ht5RNe70iXn4uz/ucY+OffM56b+zug1t0wOv69RfZW
MWbK66jgDYVIMMHm5ftW0t+VdMNTrfSFH8rBvwjSphJDL8o/MIiEoGinwpopK4x6XVi8XWKMDs4a
f6FW+2PAz+4zFQ4CeZHEvDaQCD6UH3UpeQ188QQMCRFSC67uaA1ViceATz4Wkvmg/Q2KSyTYbZB3
tLkC9VlRT+gfLRaqJtzQr4ZmZF619gZjThY7zKLm0YnFWEUSPK+Q68nc33tqIeTnFVnuNAuXF5i1
Rd7uNPHe6P01FGUnG5KR4dA3QIvtEKdVReXh+Ym1gUx7rbGPmdoIwHx9cpNr8wedXM+UbtBTTakj
MuRcs6nVUDHtDrB9bZ26gUllv4mqEHp/Yfc085lvG/TWr7UeteGBCmjhiT5f4dZv6CFwo00lQcSX
7H9dYapv4aRSuiG6vRE0n9Zs90a28jr99D5RIjpe0rhMCBUQe6zgbrqPsxGB/EZLowx8lgHj/s9W
9kJEiRWpAbQDvou4bY+5RG9HfK0rv8sLpZ2m6MVdH8WbPyKScPW3C1XzWW+03uYZgYX1HtIV5YHy
Kd+RhuoIBVtBZ9Qk/FphSGLMBrNBYI4ZVsKMnRDmwDgb853NFJt9S6cgok5NK8Rnf+3A/9xe/JSV
Kd26Wb3aiUVM1ai6Ku9iFCKP2RoItY605S3z0OH5+PbAVVxTupuz5rWXy8r/H3HsbB9/qxxr1rER
wPNAT3lXBq1Mw6cpsa5BKc0EzAYIy4pM4I4u/ChqcDQy10pWRCt+2HeuvniIONz0+7v/HKF2k3VJ
wfcRM/UqTvsXFchEsBPMsiDhEDnIn2iNR40/d3v3hu5YtU46/8fRpQ344SaciKX52T0WCmlOmdxr
PUqlVwbWo1rcsFR4rM3piAxDFqqgvBrvruLdevUqn8QJW25iwgCKiN7VvSS7JadA173VHAcmNJCa
2SFALzfkimCsaYXbITBdK9Uuo8I8AzWawm9DjN8aBZgLkc0irwm5z78HoCqoSwt32haCM/fZyKH2
LRGN5p7hXMpueuMS2P4ZkzWcvxuYw7BcTxPUmJzKYOG3HjGaAcTRsVzUmij9nLyxFCwmZfX52i1g
+Fli4TlwLNV4DWNs0vhcFLW+rkP6cmD0xyVkuz25kOQ8VCOIuBjUV3lPIHVSC41006/g3oC/L4rZ
wcj+pWIlLJilPDw99mbP73A0vGDtbdlxHthW8jRAMOBJZcHYMrxBShtCJsSZGg1DtVYHkoDgbkhJ
6RIPGZyWnZ0sq2wLQ7EwOl7OIxgxbEfpBNgTIxxddSu1NKAWethAc83K05YPhaLWw1a03hdymFeI
nhIUEZRKP4sYHs82oNMntmnoXCjxNo0HF4aRMrdX4rLBgweaYuOspW8RYU+cWu/lTMPWnVIOXLUK
3FNtEL8BPqFHkPU7Tu1suklEi+fx/g44G7TCY4wDkwUU0Ex1ho9yR6xJtMp+NtJWJXmx7MensMxB
h01d2oeh5rT9T1LpaEfZoRpdlItBCsd0thp7PRF3SbW1fuvCsXAZ3xiI6lT4Hdl7cq3TeNe0mJSY
kJo4YRuihaR7C4EujT7UFwPYrKH9cr8KhJbwVUs+Y5Xqang/eoH5w+oUuwTJe7P1KDhshP97xxbG
8NUDbgiJs4i7I85mTHL1m29vWQJmRU9bQsqNd7gv+veH2UpI8IreeYu5KDcd+jZ6rI3MHfbbdGCU
1lnAgrjBDWJz3vxPAlFCr+8KRjQEjf6QjSkdbOTUnoihMqXkcDZBn4bTQp3DT5KdV+9HOrSlrqi9
XyJbK8sr1/Lfs5sWNQAlA6dAINNJ63xW3zA7SoOVYpT3raXB9wtamPc4tX2EANFdww8v9SodEjkl
lu4ces/lfCzJmnFg3J9nUijtP/+rdktRRGw/aTzgYRBw4woo58ea0xUc1UDf+10UV3RoNoSgb0h8
ejioxatDQTwAj72jHqLEfCXwxpa42GjFwMHFayXj58CCZySSupBjBijizr3zyW3kCZV8mL1BEByk
+TFWYKboKHr/IR2pZRQrfdjHUAS4SxOnkV8yf1gjCsQl9cWUyf++agAEHgXDiERNFftFh8uRRMgF
dzZGs6ZQ4960xMlMD+DoWWt1+u3EWPzRp9zp9VINuJsUdDreghm0atJ9hE2JGB9/FtU0lWHAAuJJ
b32QADEFyVlNs2Hu8XeuNr7dFJVgjbNVixmaWNEtAZXyr9IMOsu+8PWol8mnaAH8rvUI472+K5I5
GoiTL2hUI9HF9LrfGHyi3ntbbvr7jmguzrTY0LUwtzMmPVaVFQG5Yy+GuRAolSEmMTaipc3J6Kld
U8HX27Xw8fRt2xDYiFr9m10N0FljSf9I4DHKHmcjiGqOEj+cRjTRsVzeocYTQNXIMTw4GaHyQMX2
pmzJOoNgyqT+QBXgoqpgv+RZL402p9LHbgYJ5/EPBUFLQ1uG5TT+GI0+pgnlYhiBLTbQLB5v2EFC
2XgzEKpB/lTC7iYFGuUeaLzPOO1HgvS9mBpXGIhh7S0HVvn0jYmb9K2MAmO2qddwjSRV6kkJL/C4
3i46KwNK4T60Q4x4WgJyW2XNLpvvwT9/JUBsKXapron67DK+LDETPwwvuN0UhKNuyqeMBzIFuZXM
wIME/p7azuqe0LQYqLbnejiJktOQhVh/PcrfEK7V8HWbfoXkrgafZ2T0iLlMiF0+lhLMfxgBpz4V
rcu9DqqTvxIRhPi43UWNNHBY6FRShzyu99JWprJY5Rc2Dhfz4RPI8MhHRmqFgOEkD1FVb/Styx9e
yJvdnRiqabOIf7wBw2GTh7okZPrM5ohbv0u8wuukhi6bV9BwGdtD7dzRX2zsvyiqR8icCNS30TBI
d4gLVvohWHS2aBk78W9h5o2Fx3b37wyPxRwEEgyM8KF5iEK4QFnNpJaKKfUfndrZK9LeeASHFbfI
/eDzg7CvPkO59skXJ8jL78RbPeLlcN1PaYFsrmVW/7cUFJaaGyiq6plXVQFrOdqdRfUz02FjG/Y2
ERedFJYzIKIuBqdFyTP+nuHsBcaUgsuEF9GMRGIoo4p9gnAAIeBuwsO5wE++Tp1gc4lKHBx/UmxD
Poyvttzw27Cjy5nDywAx28jP6NlH38p6os1LLPLCQ3dzFq+P45nnfhIgbPKePq2isB3zFFPDuIaB
87lRIrZ+FIAAa1TAwDmPK75DRoE+GIxJDCSV/FzO5pEWjdyYIeFd7Qc8m49zaGCwN0IiLd1v1Y2R
iEG4A9LE0EfXp6yAB9PH2Q7/13/eDzSVJGRtvpZ5nEjWUejqrhOAaiKnt9QdYfuJfYUchyLvXve9
qRelE8BO8vBiJrpIjRfVvxlDs9EbEPboh2vzhvJxJmO3uopUUvQDkvTfKI1EVvGFfU+tP0mwHXk7
VPpZWGaaXRCUEl17+2HpdUKHMLLMva0tn2y9BrmjfuQemP+zY+9NJHWJwXxLQa15zPoQi8gPlmXC
d2tCBj85AAiwRqzFF850e7bNRFaQzD7YuWAxuiqwoBe8xWWeDLocXzh9BxSqTB6v+zH/IzcODJ/L
uqOGxANeBTqTgjnud0K433yB1+I/4DkMazyUEutGx954bg0Zb9OwF+KePjPJh2KGFSfhzram9Euj
SCXCHATFW/rWQUXsBgDHhpDTPv+LZI7O2xqQczMNLxVellEIoGkrZcn+/s1ECFajmfnqTNO5kvrr
0Hp1WMo5M4MELuxkiX4+JUYgZAaDZjD6wOnVPA93/Kd8K35J+UyFEJ4hSMJlTsW+JZya7tknfCf7
sNhLHpKoRU//0qeSV5n0N6V+zwoKedcxpmrRjPMRwtLXpnCfaRBE5ZE0S4FlkPhltwVKpkn6J94k
90fLuW0QW04ZktR2VxgrBDjaNKQ0h9BsuQge4y7Y6ZUcwwyieVsfGSpPl9bqyKslwlWBUNl8T0Lr
Z48mTX+AjsfWcOxrlMDsg8et0/BhseU2BjCpOMfYRHimGQSy/cYqW6aQbmfgmLGX7vkfGCLgAIFz
M3MooJdxgMB2NW3ZEjuI0U+FQxToPSO+Vl7N0A/tNyoteGnz926S34T2NCVFu66X64hOASKdSqlO
aOOtIk4+7SDTarmYXgNqYyxoTRWENe/aI/SR2MHTZpV7/Mq/o6N/Bs1mgMPbr5jnZx6nq28RrTGn
ezhVXhhUZuknqEtUlhvj/4EHqFpLf/oucak66dHbCLcrrTpvE3a4/LFIHltpI04paU76990J4ckf
2cSzk0OtlQEJVsa7ZlM6U9Ao2LSa2TAZ4sgruTHnl3G8pl12r1Dgsu/IybMZQFOdgiHOs5/aCTKu
RQ6CePk0VdfrWoTsRmC3oCVyPCd23gDWzMqFeBXJTVe2VRLH9Gh0AQoaxWjpjY2PsmLG9uD2qha2
p64rWSSUEj5cVz2mU96MIeGX+qhOa4jruEwFJPI/wsMlvyyxyY2RuV8Jf3JOcSyUQ7WQzhN4ba15
+wL6P4IRnm4lnWmYiDdgC2HzfDpYyfnApggFm6qc/QzBuhudcVmA7KsY7VjMQ5B2DWhlHxJkLMaY
jmuOiSYLeHrcHp9WzO/Cx/kjbUOGagzS0mDS1qWlFn4QiLGigMSxkVhP0+MCiGaG1sh8Oln/xEaA
2ACEUcnCI5j4DHcdla235WKwX1Brgg+DuxIOjv0ghJHgikcawU+mCyhkO//dsJMe+JblU2vI3TKT
NAwpOqkYheYKOzCwMTfUmYlcWLQO1NkShhz6yRuSDmKF8L3Tur6haPJ56Qn9qCtApxesqmr3nNZf
u8Cub/HVbdoB/C9+MOuAk9pC9ZAM6EGY+nz6PQaei/qllIumAs6GCFSpmLnYal2y3j5pakR/vmjC
aFxdVlhr1OJ2jKqFIZidz88DBQ14hYg7URh6yo2TVQ/3Shl51yvyXHi9QZqjY7DlTRmlqINW3pN2
+t8XP6FVHmRiAYfigkAaqj2tIVUWK5XmpL9d+C2f1XeU/m/Xm/k7U3hfoMB/L/lsXK9gSz4lIqeY
gIuRAUsXtK3vMIr8tHgUKHSEsZdC+bmUapl3X7NRWWTaQYDxguY7lJe4qHK623fNVpp/xiZgiYcG
JxXvgOfBw0neG1wk+aM20yAn/A/0aaoNGkRi9hc9QJFHRE1FRDSMW+gMkSzewx/k+iph7wZhp6X3
qukGkmzHG0zNVKfqtmPjyno0UP9t11s8J0TXzKXqY/kw+2NbjYtJmXAnmjc+PBOazEqEOVyCuNsy
QEpGwIL2RQT7ddfYZtvSWmA+unV80FCEEcCzMQMWDbBt6BXF1VU5PdtcHOdKxaJY0q9ujZw/tkhB
TD11UHkCPk3a0sCTeEfycuxNR4MfYEiAPGmL7ysiNZ1fjaAu2HTQs62wFFIq8EgW/rZTXjg8JObq
/CWwgbn9GvtQDTa7Ii8qUrLdM/RlmGSFSX5rXiloRq9A3SEFiIJiXTfQE1M5bNhqOHxfxtgJ3aq2
XGltPcgJMMw3GYe27IyhhWVrNtGhpeNjBxn3aXhhImsnyq9br+FF0hLUI0QkNz7njNAbteeZfol8
TexTcnjnhLuoxpnijzDbP3Z1CoDikWctnU5Uu/qIkHvH3pa1B0zjOiluRAZJ13FkhDeFnlZC0m/P
Dao/bls8mDTOhD2MeiaybFNQVkKivPvBJABzfy6VFtcUFaFHujpIS957y/rYam51arWdeZ9C0Wlv
BNh3Trx/vmdA2Hjp5DP1v9tgAb4bmLi1LWurboH+JoUY6VPWL7VizwGFBlWAiQtgiKm1xrrPrLcw
AmQV3jVhup6Oe+/EXn6IIO1pPNyPbCpcXZ3YQbGc8yDW0UJ0X38TPxtQd9NssClQT4CSFJCgQI/E
5z6k1Mtb7/AoN6OrOod7lPMRhWbTEOkmjHNe0wVXrXl4DjY8+c3cJNV9nab9PuGcitIvD5nlALpd
l911UCrY6yKZWTl7TMqfyFfMw6dLM8+Pq5RrJr91YoHuyzJz91D8nH4BXCY56qBtOcydg0rfHvYO
lzixe3DpyidPu6xXR4vf0B4uHOy8vT9PQ2b8yMdYMnacywbxUkKHvrgv1N9zBMMs2rj/ut8XypG1
NawCD22QqR6j4BUA/y5ZNgnrKL56oNionzxAQ1+PypvlFToi3tBNB2Ih/5C6XmpL3VHZUYIjKyk7
hZMk47qEYA2SEr+0c941k6sBdZte9ux2FuWY+p203HGPtHWvnlFpcPqluEfxgG6t3P+QYAkKJS7O
J6gHOmSm2raIi9Ob2yDNQN+5vxMlQsor/T9SJcS6RtqdIOmAscXwJFXdXV7pCTIe3RtTw21E7BU2
mqRI6adgUfZKS8hbDbAYtZWOB4MHmgIC6R3hZ7ygcQAonP/hG2E0qjzYs9ajgtTIOXll9C7N0IVZ
radDgl44t//8ImrhlSR3YyzhOJ8WNxqeRX4L/qYeREh89C2Rr/NGylVqukqtW43SOrgPP+75hrbA
wEzEBgLPMZ66/6qYP8ZiyaJxcP1CF0+PDtiiYZO3ZFULm/0cKNp10X3oIPHQLMdnYjriKyLvKum8
UNEnZJYfXEgTQuaQwMFtWS38DUsn8Ybry9j8AGMFEYNGZq7aV/WxmpXFNnpVWCSfnw4xL+NVyy6u
iPXUJnU8Td+FnFvuxbwxqg1YchMCOF7LrbaPbxChoVz4pykNHHeZzUm8DDZ/qGqHOr8oENeLb6Ja
WWee1c/ZFNzjxQZebGK83e5ot1/jTAUCTkEklJaQBbM2Qxxy7y2NpS0r4VQEEVZu6EYjvrB1HHHw
k/fC5UiVlFghAG24UOdExcrkAzxHaw+BaD1G3dbg20IlPzlVd+sPyx+AXMKFAYmumO3cEF5Pvw+u
MQOpDcDv+oUKIUMDvWR4LJ6ODMWe4Av0EvqWxxuoGSacNr/Z4kd+TMiZxcnKsKKk+fhdGnSzASTI
52esNbC8P2+Qxd5/EAZUzlO/HnKrqmPoZ+2LhL/mYiaYSi28T8XL7Gx+hrx0Iz3NqtOtzOi2qb4z
R+hS82j7q58sf4QpFYsvqkPPxPf9o9tru3kWDWb8ARa4LuewK50ShVbM3q4PVTAk+aO9kUWS5AdJ
8j7Ppp9fXFGuCUy1bz4GwD0U8WJhrW4leKAn2KXCNIFGrUl8p2rJS3Mi3nY1/j1OKGOBW5WO/X/4
rfRgggj3XKmtG0e9NX3EaHN6DZLU7xaALVFnZMVAvhyUswtTflDfusxFy0MSk6hIq96m5TTG/mZM
qguoacT4jTa+ZejSVHwN0P8xwwLrhhOyni+D0AacJAmLdFjD6AE6j5mGkZVPcymu5OcpvgHTOJLO
KiG9BrB0eLGe5RXkv5N5mvV6NkNnos+6zep8JDKHWYj3wa/4SdvHyeaVFnLYkKLSXnuG9AjIbzDL
7VVK0mFeHr/3IdcRP83C3CQV8x2zRc8RJG14RNSJNtCtmhiapFKYbtiT8GC2mfO0tDlazwSb+nnn
ELHe98c6vGGOjY9D6EpsiYZngFOds2JBZb34Id0G+o70SVQw9TIe3JaQCbiEKyd48kMIUheOlqhD
dxHAa3zg4C5cRoj/uOWoKx5HP8N7OohJX1XGvRc8SemfuPh3jsolupktKlJcuoHfrylU73MHgYU0
j23rIKZFTCLZ9AzhyLeV1DbHOvA+SSrg5ZFHd7qfpLLvTzG+G6cVIQOUJPDGcRWb6hBrGEHMhMq1
510rszcuJBqBaTTa3Fkfk0f9sWHjQQZVVtt99sFmF/LnJRlldSNSf3zdD1DCrHrM+zlzW19S+r4f
st1g9Tx9Ir5l9YOO/i6yHW9SsBzq4JonIYYi6Eq+lR0031o0sxvxGB3N2lgf8bkghfWU5sSpRs7I
1gwABfoaN7s0TCY0dejJV4AUMkq1h4p4g5YY0gbkFxV2AdvNJD80GGEGKDEjJQSphnEC0XOfd0Xb
rHvg3NsqZJiAQqxVQiubzDpqGQyaNEDe+4z2zk3sQYGZFdeiSdlkV/PScjT95Vv/sqgx4grBxfCe
Jj53xxF+omhu9xO+rwxkuiN/8fOfQ1E2VECNC9LpHU7PJoW3b8ItuqPN+SUvb/hOYK2n67GuURRn
P97b3A0jVGOK/+5vf1Qun3oaw7x3FjvH+W7Nn/eYIdUCx9Y4OxNm0boPGMjrqwXEJaziBM3sygBn
p5h7CA1dxqlq8x4mNZCTAnQptky4lIymcZlflIuhWZ8X2M6LiRoLY8Zmuc/OzVVFO0G+hhyuXPOp
1erYRSx3Dqe1Z3s1vIGAWKkDsNxbd7nrIrfpEY2Kqm3BdScEEL9QskB3lRWJUFFgqcQplCFC6jI1
Y68HONk2Fe3Jepactsi6AKsJhLiCmv7Cnz8yLYRkUZv3AUnPrGWCgXQzd8TTLz9iKyCM8LMjLWKm
Lj769aaJF7n2Onj/nRytOg3XnMJRTzhLcbx3zCu/XUEDiLrRYVnnaiUL8rtnXAZsKGKfV+yAIldY
s7FG8tk3192SSAROV/iq9KnixB4cZreMrzHo9Vb890pYe3cz5EO8/FN4K13eVExmjgQhefS3bbPc
tjDue24usSMnx+ovlXzWv2xMqpAmc3HO5aeS01lS7w5MEy7C6qVmS0UM3RLJiihDiTr7be7Sg1Gw
hJlUzLqAzDqBJvyy5+KF5zoRTAygKGLIF5RWK7zXvnKyhvY28hoeQ0ehBTCNwqisCgmOudP9MV7H
Q01hXG53ii2Ov3iYDXL0FhVHPxm6nkAfyAdS8e/bTSjuWeFOP86lIaT0mJxgDsLz0mQldKhzGu4m
AkwNr0s3t6EXRpY0Nx9PeedB6jwpWZhpf+zBkhBijjxFEuO+uWG8d7o2qn4afgnBYm/Jjhg7+kvg
8Y+6565gCCXt4Uu3a3Job3VdFMYraZppNg2UWETiZkf7B2i1c0U/dTf+oR9Ma0ohtqMqBLMapN8s
ruAP+4NMn9rV/focb1eQ1fMhUHWmu2ePtpf6k+8xGYFQGFc/vvJ4WJu7FOaB3CmCWnERM8uuAHnv
dFIMKKjY7rb1oxZXgLLfeVr0zbyzWIFfMbXEEvy+WEU2iaFE6btn7MWF8Z4IYMPk8xD3nNJ7q+6P
E1eSmn4HVnIpOxvXfOCGaC0sKnTsY2HRttQiGXwp4y6czaMizYKKEhDwn/7/rZwRjgTYqjwn0fS2
KlRlqI2BUoQjbkJBwGquvS8rIujdVa+1kw+MJWH6o2HMmvinMO1Pw7PJHPIqWw2XGMiFjZodRt9b
tiSTB0iloI9xBBJEYjKHTjbUqIs8RLfDbsyGBtocxOsfUjv8WuyzetFazPV6fycZMRt0jD/jH7zG
KoPTM0b4SKCf9LoKdGLuRIvD9PtDTUNij9cLQyc/K8HBl52Ns6R/krbX7ZSabUIid9n1KoGneOIY
jFbA32HJQt28vEChvGc1I6VLpDCoP0JMvsyh1Qgu0LuOqKm2tapQBfvMhrr5c4BzvfNZn9hJmZgm
XcGSuVTcue0jrk/mjZHPCLlOKLP5ZtIGjwy/s8iEcP5xXP8cQHGRflgh4B2Ijh1C9Gn2y1D0yC2s
AptXE95QSNYnK5lZzh1mADPlvRE+YgcChjS9Og2jnfb1qGzZAf7/l5lqIwmkG9M+eIbZY4W7DEu0
xUM58Gu0KSf7pN0GUIin/ZJLpstM4uu597a4NBqXQ2fFG6nmDFQQH51QIaZ7nAPZjVvyuLfOZsV5
5GgxJcPvF/4EYsdhih+DlTuxmc5zIANbYOEJuJyja3o0CxQJqY9ufjrspnawmdv3fVYFSacOJtZh
WcTk0k4m+SC5aVxWKKOL9HBIn8mmPoB7xnBw9qSkBAyae/IasOoGZX0RsQPbsT2/5dpGWL7zBMAH
QkY8EJuTToV95kudVLMDxG43xa2iwxfhwKVevPHQRjG/Hu345JEWlVufFNo0XlyCJlmQDxIsr5FL
YnG/IsAxSKi2rl2ErgKA6xXKWFv1b0yNwbs9dy1v5jlTbAoRQzdO/Jmz8zjkntR4Yo2Hq63oLuTB
VPIG+MgwxrJWqFcuRdlODrn3ihF05G5Pw8zbTJ9QnKcq6SDBLcyokSMtbshxROQXYSjoogVXovR1
oBZlxS6kCPH8FVbySzmhxWLH4TTxVOn7B0hYPb552W4Qu09zgxY1ha2lox/XNgVN738yo87eHMJv
KoEdHT63H9evGxakwKrYAGlYlv7Ome5/WRaqa3LBAX7kugJWvyKh/t+hEHjMeAdxCwShoQ5mVEXx
u/Q2LtPfDk0S9p+KWOLhtju8CbhLGezDe0kmOFglDKZAzcOjHVpt+YcjHBPdBk7hwH8kVdLXPy9x
MfXw3vWP3oKG19TtXhRkJdbpxrfj9TKhJWM7kNxQaUBEBvbdGXCw93eyBm1J2T9DabaMZM0TEb7Y
8itUEbNnG9int4OK5ksd5oe92zVwabH+/fdOgG5qED95kQ/yVfzSGVLj6c7G3YOOnkudQgV7hpEo
4Fw/drFa2/sClKsbGlVYRvEq391xX6d42KOtUItGLRIiE2DpKjwpfiUYgV+BwNpXb9CQwKJ4/W4Y
7/vBNUm6tUMrFyFVi0iOXaiRO+aK+4UBQnGRKiIRqBJvfYRKfjoktmQmrP+hDffcFZsi52g5fM3n
lo8qH9IT8mWr/l69KsFNeYsrF0CqMdbXjJu8w6gAVznK/rX+g7W95X79qZzepNvVoAwm699oy8G9
LtHATy1uHMEP0wBTjl0QQSsE9EF41f6Bblggmm73Atq2JnsPaQXmb/2NLDhQsSMFJOZC0Ssxmw5C
zFdVJMmYf/TCwZcsdo4rginl2EpjtHsXGlB4sITiGGiNEp8F4Mhx+5ffh6Fxp1nvCaB2vFyiUAMn
aNJIhOKCyIkXkG7/pPAk57ZK94DbnP24MD8jtRG3PK7b7wDan3nJcXdhuSLP1vi8CUNH1Osi38z7
7THrNrXfyhsd3P351cDMi1yoUJ3M/cem550HBfVEYsDg/5OcmUP719U/WciknkA1qHj2OpAswLJm
Fo/p4BXexQv3+EfzA3aSzh1krmc9UxWW83z0RW/QVhZZE9f5SopUcDfWtgpwBjNE8O5bUwgrVQTT
49fulpv0oInUY+lpVfDe+QUV06EigpXshG1MQnl4yaZFdRwSI3uW8U8dpPerZEMyysQ10ByL2Kky
BOCYhJTqq8FAEkcpb4KV+hKC2f+8OCMW7Rku++fkfrdMfG1BOS8t/SSqjv/D8Wm6HP8U+b7k6U6C
48Fju5Jy0+uxTx2pzdUHtUwKEOg1+2HJtVltF2c1OHNdVJYlL7/4MvlQv1g3BNAURJhWyhBp34VF
kJ+1Tid7qtw80/MD3WGUV1l5iftwD1FNLVrBNfJ+3OFqR7psO1ImDjOgNkWKto1TkXmSwQDEHDHU
qh3+Y+gDNjQhRegf2VytENFnmWYcQe4yh12ccBOW31SJqxD0quQRUwcLoZVTlB2PxhpFwcZK4rTp
0sW4aMJKuohRUsVvnpvHP53FFECY0r1i0+kqY2a6ykIE5nvuWUo2B2u8tz46exK266CA3/iLrfn/
zIIZxjTfguEQGcNuIgZ1FcCQLKBiKWoV93b3/2SN0pWyrNfS5MQMZr2MaleYz+jJ6qyOGo8LVqoH
V0Sj2Gg53a7MC+P13NAbNjXgGIwz9jgFNAwywC1ytoEuT1plEFLXXBUtWDXKnqZaBv+d//rOtCGI
b+Q/WPb3j0ewa+i0o8vtNsL9diexTSpZsea+fEIq2vpOiz028tJbZV0CaCPvULaJV91YgNcJzTQB
H1Wbb0A/sNzycj4VQc1+1z678AsA2qyrrPWh/Ed4ctiqAwFpJYJWr4qrJm3zqWKXG5EDiYU1Wjye
Zd1ecCxP8BBPsQPx+3n/4ATTyeB0h00Mlj5iv2lGYa/fwAmcYTJLsaYkE8fhlpsZXrrkGDsRBAJZ
hJhMuGyiVvfPqrTVODzQZMYK9cE8A1j4afVqyr1pDA+6lii7sKXQ44dbg5oIVmB5RS4Ia8/+oLWL
Utlmo+lhl6TZzQH37IS4njNewy45ZZj5Cw0B5lg1h/DzeNzXPk2IY8nuRKbvWotuomxlVlNsWQjy
nTuUtzYIaCv9pxrh8qMjnrOc1WuCawewuRCt+7A6UXhpul0zEzDrIVv1sCWVU4WbBXogqaG2g+cG
PSHEjcdw/yZRYf/RtPE2zKuz64yf6GQ65M3/KFvnMf7UOkkgtO7+iOx3abEXiV7VyzfWZJqKc7h7
UIAM6pZctUTh37PvY47h01sc4xPENzBOfOdKeKsTuVhooR04JgqDz5NRyPCY6Sb7BLnS2UKuRVP8
DmqnxI3/rXAQF8tHrRR2SxR3Yij8g1wqZamJDbxgJPfqBiO8PkMWpQob632KJGfhJ4aSaPi2fkBp
VwA2mTk8IFpB4ov3n/Vu4uBWjyHqbE2iisOmf5y2jeesU2gFqgWngXlmbZe+RbyE1tM8LHodVj0R
1+zw8OmgYTczs01pwyOfWoFElQQyH3ZFTPh9ejTPx/VO854rKmuEa/So/1sNUuTQFqvA8gz/2MNh
J9QJaHfFYs3H9eO1unlABIlPRHjJMSB2OsNQGPo0LgwnZGiHUx3UlmZt62XGTob6em6aM8L3QP4s
f5jqBfjsOCA7E8JTgiDjKA+MQEbWjE0SgAOkawToGtYWTvpdgc1bRWLDlMgE3Fiq8TtQKz4S4xZF
M9bA2qJkdWvwtFfUh0uta0fQ3D/AGxNnyQiFusg0HrM/lTdiuk39uUhDyOPOXDpiI5bnErOcMi/I
Rm7vH4SsSN1COFMo+0y7MF5FeQEfi2LWavP/5S6vvKEEL3uCrpX+nVyRiqNFhkrVopNSKV94gDWT
kQbsM3MxUX73fWmkQqHLZvRcDeTpvjEYzoL8c6Da1Ir9np6EvIQwRg16fdzqHKf0269HjhldYqR1
FnS7Ogla0C6TAjXL0wlUxdzjj2bh/A3gJ0mQCJzU5/RcMlLrNMBIR1NUZvzHQ2LqgK8802l1fyBg
q2yw0c+kWxZSVcFtGYKBhQJVzBZP/8BCoieSTXeCWwruNqfKJdbUaJptkBR8R5FtutSuwKQmtlA1
3FrtoQpJzC5KL94k5TvsHmb2jmToKOW/ol/ZzSKU1eqat3t3v/u53iFx9Nj+dirxnH7nV/5Y/8iE
Jpm1UmMXw5j0Da+kwh4cE/FeV7UofVxW2uS7rVvRX1BguOZryUrKy4wy41sYKsp34drTcF8RDooX
mVpsddyXme9AO8j1RFDzQ/S694RGJudn9dnEyDWXY4TLZzXGcmZaNTsiQdjq6dFWcZEDJRP9J2+0
vohQxMClzEqR4S8uVkPg+6yKKXTU8X4B0aztIP0/E+4TNJ+DvHMNpoFnE90f7uXx9+nh++Sw/pzI
GLkOVKjtt5OUJ6e67TBAmmbAz9KY5yCxinslz+JyHeasiVFfntB0Pyo1iS7m8ipjt/p/be0m5njq
UD971GQpLUFN4WjneDK7/6rINTLUT+v5gGO19HHcz6h5sMraGJeEy82sCiEgN6WU2Q1fPbEYLPtj
2p24ufeh/H5n++6i3FqNzshM3jE9rjKv9mMsXJP8a169nDG7/H4elqVVtZ0RrDB7x8+QkGL4MRxm
+Y1AE4FVylasI0MX2KvNMAjVbIqj5XtuwGJ1+PEUNV+053VJKVTJvXFzyKDWXUq5iZP9fFbK53Im
BcnzSOa6R5kiXvWm8xu80dlwwEWlzomZwWUgP3L5Bijwh8dzuQJ5hf0i8+ofgvNgdnr4aYiOqPIE
oG0HzStlm4ptg/jH4U4KBSZkbq4mn6MWrsi0BV46QfckwTgvGoC0YSD3PcZjUYTzVZ+pTOUl/9h0
aNuIU3C08N8jvNpQK8lzRKp4mV/2hQIhWkL2XKcH1dn+zShnNSBdiXBxcllhFpHg7/7OKRfkaNmH
lpJytOtZ7uruBhE9bpDD/XG9JLVHgffKti+NUHciozlkyDE24x6reAOLv7qojigvvadpNuEOq5Jn
b0AzJ3L6KpX+XlhnJBQ3EzvApHe3ResJt3JTVQl58S/GkgStYWD3WfPvnBp9j1uFBgIu8jXTKnOb
kDJQYTL2wx2fbQmobNjLQHh6oT91WOqRty6Plr5iLNBydwnuxTSU8gDXdpaBFwu7mjDEVjyUZQt6
IHZ4HtfyoF+rcotogU//VrckbIMqNZsOaB8IaMd9TjbsUC1GpdzN/dn0GgUhNBGwdVfwgD4ZzrQE
8lRVSELgWV/h+/XbxzBT0FzHVYwQKDZ1HIJlgpY00tAiTFLAtANEKrnkKPXoUnzNritzt+3q9s+t
KlB2LjJHx8q5jz6BPwEHYBb1OsRp7CNeC1Pc+wT69TjnkYDMLgENX8/m7fPajH3OHSHuXH0kMltC
I62ZUGt5ru3ppRjkH65uz1/ihwUpLvWKmEH2lspG+OweP17ymMwsE81saUvhVa3VCJgWRYPKOb8I
FOSWcKCOUrLv432vNDcbTqE/655yS7UFXxWmBFzAkVLbF9JNVwrYE9ZzyHeKqt9Cv/GC8JvLcL7i
rU2AWH7abWnZoxVjkecyc7WF6GxQKRQghvT6JZHW9JjzI0qp+8dCgQ8v01O7E7lXTW/EuPlZHO+3
Y68mvD/gtz1JyfCp40bhcbE3y1W1CAkjROfbX7TMW/Key0cnIyLmPsKxLKQfV4M0IUgZsDCCpjaV
b92hNBKBKkIgQdWB5duXT+2mvgaKFg8xdrOm0Am9vKLme5Z+WQZdlD+iE0OlreeieWCTB6B9k81d
DGWNoxebl6GJG1X5hA+p/374x5E9PNPdFX69DpWfWaU/oYTtfk+ykA4i9mcAUqksHFb52FgQJd22
6DOIs6r3Jmcug3gDGGCPzh9cE+jti0B4acTuvC25QVvvmngcEHeh7gKNsftom9UcsFHKVCNiu1UX
auK8AJAQqzS/g9oWkVAtV9m5ihL25OO87xf8BYjG8P65CFJm76QsD50PFnNWMbHxgsmvkXXzxT8+
BhY6Yi/DMoDHQ6VE4Xjl5JpeOunC+qYvT9YznI8Uw8KBifdZOZYvcNR/dyeN9OKhnbRX+6s9hFh4
MaMTwEFDS4T03aSYuwU5umwtxFdELKitgFME2U/PXTi0jFi/LorS5zSJkhJaBLhDjCqYswrmaW3z
6rnYlWpdWuT1IRL7tlojaDdMkvexZ6H+TF1dv3FysgEA8ho13B53FioBjFcbbqzAghukHVqoKHYQ
tER0awueNSBgSjJXlQSvHVpxBGDMzb+09g3bTL1Qyx6Wdisphab7+syTi2T4nDxj9T2lNjUAaviq
8QGlu4SyZUAaAFEvJWtjkkyW/0OshVkWJ9uu5SetVG9cL6DyalVjkuNUg3HFpCGUcYzg8BPzGhje
eMb6fn7HiEVLRjr1uI3HlMUDV1GN9suAryJNn9ZMGbUU3IOQdsypEgjZ/W0JgKqMqNhaAhHy92yq
fnp7AS1CfF4EvL1brZCHgH7OIsLWoFQwdydhL/C43+rjZNJPnkikQVASHzvVL3nDhW+W2344nr17
tNl5hQJcxWxWCC2GY5Y320RgkGr6I4bcRsa2+854RkAohAtRn5kXR3fAL+R9w1p4gBMDTnLJIc/4
OMko5N6PcX7A+Yjh/qJbHunoeFvmnAxwBVvoZfvpxdrxPg/Jn/gaxOCShtYk7m86+BimJYS0rFCX
tDvHvrNRMlsBVE7ADUa8yOrgv37GYckwQzmxL+ngynhD8EAtef9xO9Vt4ZA6FZ/VP81cCjFG+yFF
m1Z1lR1RL8OVRQTBaiAY5HcKWzAli/Jn0Vp2iaVD9/wgE+H69h0aGCLKDgon+vzhSI2AORwiap9r
AzUT3ynEG7cy2B/18Z143hXi3grdDuP64/ACnfuTeCyGA+495gQXtyFZYsCjoNA0yHsMw4CjMg1d
7ZxZRNJFNdg8aZ2Bdub/V5vtOb7JI2GbS+67w3le+HmCOcFG5EbYFbxixM2iyc+dMJnoCyj4vXc9
F4nRTel0LRMcjrrgn4XHyUsgqdQ7emNwa1ozGOY+rugWNV2zxidGLr2S54m1Ruo+VOLHYrfADhv6
+m4GIcJBHpuAt0oTCSMZHKGusJKZTpHlSxB7w3X6C1ITYrax5TI3hzPdLSq9MSPcDKCF3va3E6rT
wJJKpA13Y+mV5nDSL8bK34+ubGS2Y5q5Gm5/pzQOgbPkalbP/DZ5AY73Ac2MP5PV8RkXPTvTLNmG
gGpZroqHvsEb+fLMXud2ueee/cYOt38RcOIX0dXZfWM6Z0PLHCFHPOUfn/rX+VvPXdwu+uME/OZ5
SlialPRPUweJWH66q9UD6Pl6OEQvsa3heJ0i1IOmkq9IRvWoQgwAIU7x8KJ89oXfXTx5x8ccfJ9B
Qv+sJOBzrEQhs7QIENe3lHgSMzxMLiNJ1FOpb9fVd6ulWrAXJgXuZQtTw6+aMxHPtIxiC9TbyzC+
1ADGvfe0PwOAcVoFaFnPDe25clnnReyeGChM6cCJH2SlVac+Wt70JzkTuysG2W1bkJYEFLaagMEY
cqWl5c7Z6i+CJYGybQ7O/8yUF9EtTcHfnM8o8T3FubXYAFUkwGGYZRarObbLhnJyi4NwaKbJj+hZ
QTWDGe2ywYoNlyHJ1OvjovziMNTXFKY5btdZMxKNJZk/CmHJiG0Qhqd+BLmrITeTJyiO10SG1xAJ
/xVEVm/yCGa4M1F0d2KkufUZDEI8bOQW37NlnriUxWXwGLBZXHqzAbSRzERQqRy/iABCRWB9s+rQ
twCFZVq/4LOX+Nlc79VpklFbC00JDzvHHDOjTd84PPoPrubgxK9bWF+Sp28x37faAaJoGCDUOLM6
aNhzFog94XrZuqAg1Lh9s+ojZS7H5HRv0vJbUJSPt1w1yA+GS48xaZyeVu/CyJpmiQUWwnmzZnVv
hIOZwDC70uOrsHYQRZMfNLK0tSkMeNNFnnRfOm6jeuaDQcql4AeBiFnxpmyhv9UeTd2v9L7MNl/i
ErsEimIo0sPCXNqU0o+Xd+5sINwRDLjRV8lvw40q4KwkXSMejQ2Yd0+CU4Bw8/6ReN0eH3GIilOK
KRK880ZKIguWOA6SOaXwb8H7USbMazmHCx2vQWXqDleIMJpUvFGYBPJ3KLZVO0OBkck3z8LNkKum
mYcHus7nosWvMiQtoa0Jxl/mh9ncTRPMb8GldSEtMkbYJy5vKzahmYY/P1HwDZpTAjfdQVK0anUJ
Gz+tmmAqSpO+yW3zj9EoJI1dBrMk1RLyZA3lM6zxMhi5LpopWozsK28AdUVzOny0P7PCnWO4F6Jk
zozM4UnxC8P2XTh/2A470Il+xTEQCq9C5g9fEpT5YYxnd6Fl3Q1ceqSWpF2ElPDH8B/f9ygammsO
rVvMjK7z1rsVxHhitsc4vc1+FRAO6pBGYHnUKSwBmJgJIqbrcVeKr50o9lm8jUSrClyxu2esOMR9
wByYeq5cWtqomzBO9uJJYL6VzJBfVo00JcmiccE+ZGo+6HJhQTU92sFASySqpdA3340Hkd5vuUaV
varbcJfsSqjzpGFMgdQnO/gL6hFU1cDNU7eB7Gg3yHwoYnf6pjXkyTlAMjo/8xr2s+11+wiyiBGb
wN9yU/PnqzJdnK3+qbAGiqCtgta8wtteUU0IaCm3riRueh4TBYR3EqE8C1V2l8dohJtecZI1phaH
0i5eVxE0YaPLI9W3tUaUlYIixUKP6tx++Pi8e11ETEloIIZCkP2aIACufLvc92UAP/GkPo1nY4tI
oUwP/HtOH0A3CRIRdDTwJBnB86U2+kbXSy3QrxjUHWKbxAoLiW0MUKan94ww9iMGKEOTK0K3AVjX
sb1Fe4s4JIc7BqCTFJzWEQ2oqL/N0ScV6wJE1hQqj4JIckmMPKJwhjH69/FxJx/PJJPG1tlBCaCP
BVelLbWbzoIifFIEDYLMFJICVUji5DEE95eyKa8vD/HgzTudFXgpBjSSPLokjzGzJQ4dwi3uw4cr
CMyaX4gjJrdYJLEoKonB8rwEN0AiOq0rNm9zPd7hdCGtVFLLw6l/XqF9tpDkPEB920fF0gtjfVe6
DfToDdh5vkagrBmtCdR7QTHD0rw+xEB6/oizt7pzUOPUjuXUBH7SzNL/r/skWpK8peleEUpX7hja
wwP6Jf4epHVyaedgxrHi5pmLGRgYe0Oeqa5F219rwbmlqrKqYVhD1I4bg8x/tq90QcaK2G9cyPrz
9UD8nvDf3zxQCRa0ixULXEIkncPl9Or8zdce9qDkNLTl+xQdEdnJw0hEDueqcqeoboI4+Or4Wnpd
U1hKJlea3yg/mterxyJdKO8JNHIpiCZ8y2bOzYErBwA2qhI07eF5K3qDI9JFXifqBEGJzqWK/CXm
u7Y6qT1dX7CsTqlaCd1CNctYN9PoD07vrzRlHHRQVFXL9jk6T4FeD4DpGgC1vuQBcU8Ieq3vybby
rGH+HMYtSccvI35W1jm7EceNEMwyun1HBep2A7bs+JlpZHGoRclU4llSHfbNhQY62xE5TesI6dE0
AeRvUGz8DyAgzxqbvDw6zrBiubTSx9YqWeLc1a8jE5TJGoGDDrEpt2nTuLHn0frH1Gm5Te9eMQ/r
EVwb5dHSkbYhEmOSwJZ3hg0B0+ijziNlsTwugAK48FOIcpQvMiwsYvVL/fjG3Vkrqf/ps2w425Nv
GANFH3EIVUOewIQwFJGWqYHsLjGoWkaEX6fv4prrYDy2862FRqr+42Xbk94ZKxLR7uEWvjsey1qe
UkM69EfTEqgcHVVIyjsl5756KRJ5WlLnsn4jyz8C1wA3jGCvXlU4B6RYcwVA2NBLnHcc/kNxhgt1
BX4EvtJ4tB4iVFmoQQBdjxowpCCpkKRZLgfPN9DIAfJE8FAOOdgrhVz1ldPYWOIacJ/FIqlbJtec
XZD2PEeY6Wq1t3rzdFeChT2kZxGLZGlNhEVdclHrH0re055VO9TIzjHA1bHADMLuq5l257T9WpHO
N1+H5fo3MYrptR191Wfui9SaQ8sbFh/SE53ZQpUt/2ebN2GmJzTXi+c0e+3ZHKQCNMRpfytoBGCE
3bsLEVTrb9g/Db+R4Ezq44uAOi8DjIdRSQl7hckk9PRsxhoSUtETDgHScZzCTXEH4j1pWHfHGucc
sgFupq8JCI+D9SMdVAePYoQ/XYKgUtcNean/FabOd6h97bezkrAu1JVzKlvbcEUrtetT3a2DhDpT
SqRORu73WOt4acPyqAoQwRvfl8FsjIhy6M57HyTwSst1QWuRLgNJcwmyjXKeNq1hckr8XaTvMzsp
0aLBWMU6LLjjkS7ZCRYB5fsHM38ymnX0I1fCOoResFEk4eselGyyWtS1zc1nGXquhDxEsQ101cGt
EhlPNUlWGmDap0EdMe581DQV+OM92tV2e91U007se24mud8zOU/anY7eo0rgJRZ+BgUjKYsksjeT
cSdXxCglem8e2Cl15VwBcqd3T4djjNNkgkqKI4V7exFnOdH7fOXlZHAsFFhkG63ydU1ygjjguOq/
TL5H38BuhSJ7SFxwg5561JF/oFoxw0tl3NjFkfq4riRm2WLujklh9lJCC1Vg0TSEnW5/iGrLUFYA
ApeFu6PwiIodBDH4ziJjzgxa38QFRnPO8947debn4FdGuAq/lGxPe1/towRv8zZE6Ffi9QSaVAel
qay5Ode/oihxj4VX5xEr3vW+v3SxH9dHG770Dwtx0R7suRVA1AUKEnPMzyzzxpThKJvSkomnqkDG
b3JZDLGvpbAJQb66ZywCFy6NqDyeyMM0Q/NlZ+Qdu+kS+TWZeYl+PqWQoOAxiEXsN9MpeCENSJqe
sWN1yUfx51nL4vbixeqpbxrkJ0y2HBqHZ8TJxMp6kuZIMrDlSQWEHLEIr+XJt8blT0eC7GKW1/pb
Db8TP/XHld8yjH2LDxwQztwppPSqIJMas69sJAcKJmcl5DFxDG8jIRat3MR0eqHj1j75ZJNGN7oj
JQ6ip3qdHg6/T/+0h61Kjf/bBrSjQ0RXPSG4zRSsRCGq6YYplnk5+e6b76z308FCETkhL1sSSsWf
1cJtRHMYC50r8z31sr+T9dZCPv//Y45z6b+r5fOjE6f74g3fgGJRjmzuy3/1p4UEpTfmZDF/uceX
DjMJPAhnZvA8zmwVP8aD5EUdUVzaRbh0j+p0TQE5v2ttfr9KVAP+d3N56gnONO7n5u/EqBB49a8P
PS9IE6EwIhw2Khx6zor4uvCZkFiJ0qMpK1y/Y3qVK5IT5++wvSXQOGqlqCqrD2DTyW/pNqOZ9B53
9TPRm5OnNTAukQvvp6maGmO/aFhxPDVIOkXIi+RI546JOyNefYJyw6YAhEGBo/+QNZ+DUzkSDcQT
VE6DCNklQIRDbKM/qVofJFQ+cknuu8XaViIhB/6U69Cn64XWMHaXYbnX/yFiNYunjaux08SYhU6h
RGxCD7OKd8/BCbvfdqDq2Z51lKpkvCUIEE9NtkH9Z07GU5zrGY7CYHDZyA7lVFI+uWTAVIuQ/RXj
bMXfe6y/qbrJv8cQIMXjzlM8iu2RUbS0nuYmWe3xBmXGAvYl1mt/pYeZuRQfpwe6VANBPiKrRBn4
eF/DCi9IJ8QlITeugXNaHAXU8v1uZZyl1HVa6rTb2WWFPu4hk1UxiCUvzsX7dILfvbkw5DzTthFL
D78iD+ddbozO0W0QensknBbBjOJ5fGQ5v6s1InvpJPHNoZxV3ph0SkfMEnz01KggtWU4lzlaLZWs
WuR7g/ALpDfv9Y1TpTkRnR5GH/qNWa5i+1jT8trrtWA8g/ds01ipGrK8zl7xvxzPx73Yl+nyVGcN
AbfasB+zc7ZarGwcU8ULh0eS1yhmip0cMJPM+3r5+7Pyo6Zm4ptHtOvb0ZKctgh6+lcAUZ9Z2xMh
w8ybB1vpcTIDsBCcze9gXyKHeDjbco5UUGgHWikZgViHn7lj/verJd++1jF8OEYtM8B4jLE3bqZL
yzPLpHSmza3B7dR5nrK43Yx17PoS3DIDAKZjW6XjZ7dyJKDLq1MIboJUaBLmvUQ9DaW7uatVhuGx
Jtf1uyZLs6EY441r90Vr8Ujkf+8QBEMGqIR8ylkbh7F/+AhKoQCerXxCOxk5dMRwz6YLUpHgiGdI
2iXtz5cR/XMvDpX3c8msHyPtKyuj098Wx4QMD2tnABIlPFDC4N+C708pYlD1Em2oeDrmhtkaKcJ7
3JwsCfwNannXzgPl8AAvrE7ebAfbOYqf/YwB817wghtkiFP22KxQDVU9g5Nx5kqTa7EuXohpXJpO
v/1CY/H1pUIpWh112l8bK0i715qGSYO967BbFftR2JjCuAg5SmADzN2VPVgT5s4kN6WD9U0l5mNf
Gzg2/BTt4c5hqiFZxRiLbuJnGBRk4fJDBX/fsGQhskwKCew2NuUr81FLF5egoNshZoxMYL19T4AM
RQ06hO+iWebn1YfdwAlQ996fZjDWOOczBHiozLNFRelLAcC1ajf+WaTf32FuaZnRsdiie5cVTmKe
IPqY51eF9Yzh/l3bEeEdjD3V71hL6M2khLPMtM86Df3+TicSgcLaW3QC9sAs87zxjhd6wXNc6WML
6dm54ckQpfQhe9YAH7clph9TtTyhHz4eCFCB1yWGNsO1Jbku1VpbqC20of5BeXJS5wsPiVIFR44M
dXUzqJ0WEQ/ozlEvdShg9do9Ka71CRTccIKIt0bLvPgtpWaquROE7WACbWRqFor9wG4e7pSj7T3x
lE5cg7xDlnG1QHpqzXp6Tb7TWtnRZzuo5QNf852Eru09rZEZTRr51Nf4Ar4zyvtNcMuuqS3otWe9
sP3UzkB3yull80pFrFDSFYm8wx0xhKLdKSUqBeMJ1XH3fNwaqQqsXR6TyFgstKUH4Mcw00yUMCR8
kBW9QLwGn/cqmr6pcNazisNu3d8Y2wu5AGpZ0Kbmbytlt9KxhGSZoOC0E+e28kjlj3wRHz7YkZir
9BexOU85DbnFWedBWp6PUo6556PVvYIbvlZaGv5UMIU4QoIT+DqUwExUW8wlp7q7iLUiORuX1+DO
Uppy7ZK1LIpBS9R55Llnmu6/2nRVRqlIqVX/5B2YdKP+runJ/Qa47wmdKGyqQdUM3vP26mvfhdYJ
5XugdL7pHmmxznncoYrWdjDIl9/NQ5/W+VE5fkFNX4F0RrPYCibSosfLierWFNtTKVo7IRWzutWU
808URExSUeoKqQlszkw8eRt76CMt3bdW9FDP3dgmX/2rk4Md4uKtbX35QYEYvEOLESegqqVJanWH
rsBcgsug157RzdWn/QTmk8A6W3yFl1xBBNNnuPFVxhUe/hm6o79g9YHcLu4eiCUwaykCrri2gGaj
ObjUc8rRNlSROJpkjZWTOX5ohCRzbNumTx6AIC5KLfOMB7MRkYkS/UDSMqpF3az/17HZe/XtJ6Le
RIc0GDGMhNu+Z5abg8hkpEiRxlz1MNjm+/StIyU18L0bLOtD+5RIPdq9XRDtOyCc27QNjQ1v6xDJ
oW3qnis3EjUrUfEAEtTixfs03ooscwpnuj1nwXzBE3pV5WfQs/oa3sYKZKO5SyelpJpzARv/DaN5
x19FJUx/hkECItDEmTitwcmJqFCPQ3kPgguJoFw9qQuHrIUPuBnG85eGkqCD/5dkGqQPJt8feucR
LLJW5hp1ARhyxJOhv6It/l9DfYwihvLOQST2b0AyjIDRDFa+Pf9vB4tsggS/hEtRXYejv8/kSGN9
pdd9yVau+NMhOLHWERWyT5jgl6mF9QR84r5uyxiBD3dBbD3iTboh1jwwAn9tCEMrJp211bRe5BiS
4WGmEd6sb2NOL8jo7fH0OZAFJKa78lru9W4LjhEd43rDrC3TqKJvPsXnHAjj5Lrq14AS3VjwpuQi
r9SD49+iwCO3ICZOQKj7cFAHphtZaqtBR6fpZJjfdzo5OsLRiW4GNGCzE1bBY3yqvmNdCRMhgVUB
r/FLpm1oR3hOTywaLr+0L7pbP2pGB4qGjGOLUXZNMZdp//V+yklPfq+atruoSvS9gVWFEX5nYcaE
rKY9iIbgUHGDav6Ke2yoBKYOvHi7FKtWFGghQRtWOnGU742A7asy1ODGgpI7mMPkS225XaMTA6XF
SaPf5KT15ws/T0XMiCT9iVteW031B1RNKtUP8QkrB4Ky8DlQnkTiDBH3LbP8/m8h7AcfXKTaAsXk
sH86A6bzWKOn5GUo7unAUNY9qfhRJeqtLQcD4dGdIJpQO/sr9KcEA3KTIsrN6koA/hXL371fiQEO
+xZKa9w9h+bZeIxquFpS0VtjtKfQJSIqomDAbcsyppaHyH5lZEUFQ0JjuPK/S2W8bDsVMYepyXCQ
ZDuvsEQoPucHYwFBAyPYvFj1JQwpeSwlmyLP/jOERAgDPxWDHRxnt6xL2kessm3sHVFG5BdyK5Ji
0Q06efgcHcYI5jszZnT7b6+I5IjZE1tU4irmv4ALRCTFn+0jSQzseU0YQ3xwakPCdwLsGSRYYMTX
YjUsU7kUSKIGS8Hmfl5p1EZkCECGp+2QjZv2/0b65ixSN8DAhjy7R2Gpiyo57MBaiOfXAlFeVfI3
kSroOXDdUWWyLJFbmDSMMjL1f6PJtlnW5Vq/UzzQCHk7fXXP3rBZLC2JXOO4kOTgsKwjrZwqDhLd
4kKSphRMTi/d8Hibi8AMa8PIBT0n1PcpWc6Y+hRvOYocXlw1wCNfj62dE6ery3Xj0gXOcIWRZ7+e
BX/67XApYldjWtQsWBr8cCDeT35j3H/pXU+Z4KoG82L7AMMQIGHhFclKMw9IAbt30nMSpr5VNpSl
qVTvnrHOsOpkYUeWcIUfJspJBDl+TIlQvl0UTTMfYOG+nfsIMeDBLwiZgAyJ9nCVnxVKKTzkOH0s
gQ7AqSvWJtm1KwwxFq/lfLtW1WbrJo2pDQqtN7VJu40L9xchP5NVAmHnBGVQk0ijBuUKN5CYMX5c
441S/Sfj28/31AKkhWOnDVvXSir+jamJBl1jWA1vWmGAJBsZVieJd1A7HI4PY675kORfY2R3b73L
mF1VWZZksrcjp2ZTae5ezt8npiEwXCJ200yc1Fn8OQPX3p9fyCYoTYBi3aaYWjbwHaNpsRnpnmL+
x7Uz8syk1uJ1zukReNzQ7+n5efWK9UaS49TZeBdOJrpwIRq3VHYccGlGoMRw7xjp4wsmO867aLR3
Rc4wR9pizKgVtburP44NfZ5MFpMsT17KNYJJYEkMGNN4269wEjUoolF6WY0qd+UidLem3benY+Q1
ZwBr4uSVDgRcVQkyebbrunWnbhMFHvwwuahS58aBlR0n/GUGoLcgFjPpnAmuL/jtl7G8OpnEIXkf
sGth5vWdZdZkapkfmMOHoxhPUqKynKZPupB/92nw2peWkBNh6TDa1qj+q725EXqSmJLdeAC1E53R
HHvOvdUmtpUmoXl+otw8j3sjmL4WGD+tKZteZpQY/0YB8pRV6Y+GvtxAr3okhaOkNs1D56FnQVY4
pfRdW+3S1D0QihcdSGlBSj9YxUg1vKoXsR2nz/0a8DWXQeO8UVsWLxcPX+DMF1kemXwuTrWOo/lY
j58o3dElkTYLFa8K77d78tVxngmyKZbkWUKGuqCTVK2xgTa/7UGYkH11M5A4rnEmwBkXE4gkj1Rx
zccgoUNETKL+0Yczbid2EU8ZeBRDQPMYRlvaqADnBeKYAPKvPUBedGcAOvfOVVjU7tev72cOiNQQ
808uHB8GNmPNXsF00ZiRlGoMvcBRvf/wb1H674gEzeprLo8a+Gng26sknTHQnKdXrizbK7dFHpd+
M2gyxGROLgMFSuNS0yAbgn6l7j1BaSQjzW2DxHTB6ay6xpX8nZcQL1hZtRrfK/Pvn7bvJVucZTET
H8ueox6FJsqeqrB9Fk5pwRot7uA/ZZrg07K9iRUjbwO0HdTKxaRACLzmYIxj/VT3Ib/bN9asLS8H
hpFXRqlGSG85pxB9KSlEpeJd/jR0ctaYn9rgGO9MuepkCcCmZJCYrwYAVLn4y6YqSQaeK4dBnzx9
VInqBl7/meBkyhAjsnPniX7i86+No4AOctoOGg+BwYsCsILG+d5de5ZuPFOkLdSmjs+FjqpZJla9
8xO95ZnB2MXhT8Bb+9mIIfP0j216YbgDbUGPmyqMP7G5kxY2eFnwo5kX5Za4FA03ymY/jWdEvkqB
xFpSNxE4Qt5GzbDGZp28lOZpGhoUYwCUS4ZXO2QXTiUGRGlnxOYR+FGkOPa4vM3Xd8oDHcY7as2T
uPkLPSA/yk8Pcb1DmRIs78kHgHdccy1Qcy52jw2X9UF4ViNVQodLKZ9DvHMwo5C8/j6WT3BErwS4
qZcpBz9YNlT07OnYdksN3xtHhE0zYaLa2OAP1FeFKu48oiEPb/CB/e2r0Os4zKtC2LTfEZar3UIW
flmj56b2joNdlkBD1st94JL/5d2Mqax77YkZFZWiTiKK6bYYlDB5/NB6/1RyGnsW0J7oGIXLydY7
72aTDhmSmuxi4BUN+7IV6ONdjPG9Pbh+IAsj2+mCB+pM4890wa92nFTIwuuivoMi5ZYYF2cgBAMP
poLUh6EQ6v81wcaHyAFYvG0Uvo8Xth4fScpJnWu+kP3yR6S8AugTFsfYq2RKVB6JaktSXM7S36ru
26QDLdYIgvZvct/7NqxuJzZad3asxi1UxGTrp2gbZtQqdIibaYnl4edjPiXBfRTW9ZoneII9Iy5u
7Dav0t0HtH4iznrVFyn01UKbFneEZwHJrQa+66PG/oifQqOzMHcMeAdYuJybipVRNolim4PTm7t/
PYZFDaTT8AYWjCLsRolQDJKYqzHLGH7Y3N18wZ3o9Let+oTmApAN99Vd20DpwrbOSpTz9TJqX35R
Re+atIODRUw1PbQB2GG4K5XFK+QYsGKdcAbKR1y/mzcItHfoQrJ2KcHHRATqzfd4PR9Ccv1T0ife
KT9STiJJ7jCcIJ+mCVq3WYGjKB5iZmSKkZw7FO6aoFRCfs3Siz0tYE/DwMaoti9MWCYxmk3yv4hR
Mhxi/88uWc5QEuEspL6qB/KPt4wF5zrhAYXV4W05Smbhk+7G/K34JzqSE6mizpk7eu8qbWnsebfx
m9pKZte729MiEloug8oZK55vO4+FS/yY2K6jtNGELNuxCX/Ax1tlqV5T0syl+093YxPwshHHELMU
saia66nXiSixuWVV0YKmyB4WxUItoPNqj/qqJZqnpjhfC7iJsQbKqEWuB+/fH1U0UxRnM6uBhiPw
4ZvfWZ384zs+SWawmNAd68wUMhwkqWI0yBK+l4iIq0QXWG3NWq5IDbqA31/IqZXIEJxo8GXa1vrQ
1uxTut3G9Fwsn3WZt4wgJXlZzSlavtRMzR32quOStonEGNK7Bsm9MWogLDXKsQ8ycnKEQAIz7Mym
pnjT7TyaZ3oR/RXONTU02SwIjvRtxOK61puymyH/fnHkWKbZ7nq/su4TLyBSD4AzVrY4uSq43KTN
Dp0z3zZGuC5YvABxa/YKT1wuZQAFf4WwAOTt7S93cSyIvoqzRtUNFsjkgaW8CA+DKFiq3SV25bg5
QRiCc+4su3ewJxsjCuSWz+KQVKrYerP0CvMH8xAKrAKZ4LhaKUKfvwtc9AZftdu65dT7GItl+WSJ
AiWIAldL895t8s6SkCM4HYcuwvstvRMc5FsfeMOlpmiRmcZ6XLXvy3L8eOLMV9pTgPRjLrTu374v
2iwSdDnhOdPP0C7ryl7BRMyA7OOdtrK6gIwQHK1sCcSKvWYBOC9njdLD4jLN+5tHMRf5wkqQSPsb
20cI4hAthkBXnRh40cqB1FNFrOkqwmO98cYzQkwiTXk2qQz4G8/lprnyuSwBu6NYcLvECq65esZR
+FjLWlSXQRKYf0N8qhk6o2r8P59XXAZTrJ5F5Nmvm+7e6uWdwMVY7j2H2pKtfN/C6k23PdIf6H44
7Ulwrth7A8LGndzcgErf8drcpa7F7FfmQb5/cHBJkL+GAnqdWm3z2NKAQI6BeIBsqcuhcgQoCLdF
79xSLkTW4R1uMm6Wiq3/9DRZhaufM6gC8zGKKOqLbWxUFbSnhsVa/WjCQEBAlEll+bJG+L4Owp7B
xnVHBRgCrtR9SXveg5E3fIPfpi0czcX+U/45utR43t8my1C2yZ9u57LAzSeOv0IlkL0JGbAv2Fds
rhGoAEh4yVMwSSVcj25UI6KxKb+sAp4sA/+++Q3tDUMg3VOxHgJUwxL9tabZsUJShwK66SaE5aN6
n18l9lH+68WMKLFD+qfdpqXr+x0IrWm4o5H5Yt+vJGy+LB/uKo5o8WH/6eXHbTXNfVKEnNA9uLxl
k8ugHj68dutRTSrs3752aweY1xXwRx5HJ7loEvrAq0CZ3EWbPheNcTWTIRS/hZZsrY/RqzNPMGDU
GWahwu2VmigRJa6D6wgs9RGGvHGR4UH4aGE/SS1KUVSKk44EWjxkSMCXTmfdnDQmii2SAcH7KwES
jIrx9Lq/8vY0YQkkF6IxtCyuq2Gg5tWaLDtVfqCyQmZ36ZbWFJ2y4rvrRHrqjqLhhOONz75B00jt
KRxCvaK2VTGZ70qYtygWkpRfckzXTFbDnYLsfNGVHhMEnPDFuspIbMJLcx8A04BkHIRrtLGi897t
8OlCcrrR2TFuF+J0k1OcKM+4XYmNOc6YdRBWDFOMW3YKdzCwqQ8RYy3mAy/71yn52EhLFHS3SrnE
E+XNlh24FUIDm0n9AapbqgoDgd+tW/RMyIsHyjSun7C1nI9NaHLobASnv7+tSr4PaZjgx+ttYsJ7
Pu5d8Ca7waSGCtKnDYO2ik68kDtYMuAPDogeyM0Kv+cyPvbkONQ0im2BnlbyYQU2MSSavO0m0Y5w
nxXPcyiIeL/coDD7oEDrg886fy8ZoX3q9QZTjQHS691czDWbTtT1W1KI6ayWGNjYK4j9rdJEbLzE
HIkSuMVZVyf2cHoaHHNut7v4AWTZeFNbv80bg+UAKjlj7Mtmu7q4jcOmif3+HRktqcTMUjlpp+G8
ow9hlrF/o7kAlxq0l3dtxnsnlatnq4v4ass6FNJPYXuZnjy4u1B+3PZksSCdP/CVUDIWeKIPpF0T
Lv0GCJaJF473hY2goltkBww0EMLMJnNcGLVLXaRwqAtClWeNeBLgpnin3DgXZDnFUV+OdHaysDt6
+jcfNSWfDufPSKcT76FIhmyau03m3hGjlm6CCbQ5rGELD3CCYWv8E2zXDK5ffVxmiog//74TEGfb
BuR3e5mZqRrcABzxiyPup7AN/sqnU1QQ/OQSU7SiBIygo4uYzKvhsJTPef0LAU6wF2klE36wd80U
Rmh9FzOnkp51OPP7yn96JZ34GHcJ84Oryk7SNTbRVajx97gCAiKIMq4dKvFW8mDogMu2nbeicDeL
ARpS0WjCDpCKLAFjNwKsvgW3cfQc4aL1Dk/CTZC7hcVQAh7rjeBlWTqzomxJma6xeduNBIjGkgGh
QMGt9hrCA7INOg/dn5TAUvK6om6ixwkEaiZnaesgfU+quVgLZzOtqhVCfKEXVz2GSXfpHO5k1BHm
syRMyILaR/K+o02MJyKxZ97waCtAgXcCUCLXaacdKLSz7V4f4FQo1j77+m2AH4x83ODSfJTKjy60
AcsYmvSbbxuVSBBYVipO21biJ1zLwPB9mA0GsSUlcHEPVNXq9Yc6tpyWn9wAftyWq93AcX0RTB3k
YZ4whrCnz8PqOJkaVYxWRbjIRlG9xDspuVLT3nwIYH68lOBd7RffE1k5QC8AMNNsnRlyNhQF0j+i
qjnGkpTAo6Yv0XlEu4wKD1ajJHne8GnyoC8gztsnkEn3UHzmkwIFdWZESrgGxW16mbfO+lLAbDXW
A89FBS386a2MQnQTjUgRkNTaJl1GxzP7T8nVG8gw0uyDOPKoQYrDsA/QMfKjlHs8IBSlrVuHC07x
LNEZAamDZLJXr9LrcLKTmx7HO+EL4VTfgYofnTlqVx9b4s15LI9QyWsHDLJWcUM8F0M6WxcZj5EQ
RxYdL+JzzChUQ/dicsFFFpbIftvWrYfNXDbR1BTdBBOS/6VrMij8fzt4E6CVErbCrQKPwcJNtqmE
9pQoLVCAb12wFUeEVak3VtqyoyKya79qgnDTedOh1pF92gwtGcDbXGjrfMQgZVEbSOi+UzKMZQ3g
Qm/80E8c41zUC2voSZ0cqZ9YXrqMtrog8at3XZ5D7ADzo1J+RpBY/s26eWUDDJMPSt4QW6xL2Vyx
pExaTX5PfxJVRcKyAImhbPumrwahjijRvr4K/AHFmry+gabgaumq7OTJp3lCLh7wnoorP/N6zzMI
ADDXM4xDQXI2knvWvLAZWge7nAqvIjKGAqqQWi1MMdrpIy9C6bSODK3lRAsUNgEBteRr69TN1BFF
98bZhYxzX48nMZFUBRwWU++RFf/cuxBvQxH2ITzAz2Eb8RNSFjiPNew9+e2cYCOHmG2bvCFnmNBf
Dsoee+d9CeoWbDxHAUZnde9Ij+lktR0bFk14ou/x2iv9bR0wqijeaXy3tK/kuq37YG1JdGPXWgwe
8xHqcR/H8lOqW1fUDYRhY3vpmhT2sM7kvaqSWQcAnWHmS1JaI4OcXm92uV4lqDLUSs2tZmPFIOn2
D6Vdg/lMGBDm/HZ5Ky+BSTlOfbFisr0nHyjJFYwhxnvpCuF975RQfTyh7vhaRP64IZuJBAXCNUJ+
L1MYFFtSf3oJvyBp92vkqcmpZYbZo5Us5p/Tx0ZqOSuKKLwJDC5lTeiI14gebNwBvY1ZaBH9mtOn
5uz7CpNyyGkoNpTC4DHD4NbdlYB7tMm5GJquCLwxHoYUO4NJYKwCsk4ihPryd4UlgtB2He3xz8nr
VvQpd9bHc7fIXwz9BNl7ioWxCDZ53OudHwF5yGGw+IkmHCPbhrtY0DiFfO1qJrxmQoBpKs4rbpsx
X+yxe5FGJiQGFDxjzXWRSVc2nxAHsa1AQ2bmuk0zDb7A56UdQfHam+TxusHWaAMkpo4TLqka2ZJg
tPqfhaTNDWCE0X5k/fLwxUn8bfIjiSZrE+gjvZ7wylZph0Y3US3N6yJXhP+0nRX6YnEkvmz3LU2J
rjG/C8NuI8YkTaJKuN/Vf3yAeZW9G9jCzx7Z1RVbSneadPPk7lGsoe6Ef3Ym7GVf4fO8OPUUSD+9
2Op9SjWOZX9nL+oAaJe1+bMrR9jnKr63UKJs6GlF1bDBiHWwijHaIkyAiniWdMHaHQYrRPvQ58wl
Q3RJ0m4ogkfXaCrxAhIYyHWDAillWR+EniiQL4c4RfeLJekolS8CsZPZRnHJnpVwBjlkP9gOPGCG
IKi2k6TCmoIKx9WSFg3lUHaHVRotm+8oa2tpx+NlWYRf2RHId92fUPcGJF6dwjNew1YA5sshDkLg
PUHIiU/jEN/oPhN0vdyfrlNWhPpLdZjI/XeUJbmK4jRMZt2ip7CuKDxw1FqsNs3uCrcdID6XKFX1
Gz++IJPL6rHRNCLSgqxW9X0QntZC1w8CTGrbLSqWGr4mSW1gYfyqrR9Ic2Dar6PWe7WfUxNiiM1Z
BCtzuH0cYhyDjg6gWAYH2RP5m7L62bNeEd8OnCzed24uayEqBknnzmjcE14uP8g9n0om6EKzX1TA
L5hEKS04/c8PltoaZGkcM5kPw4qKzRn75SaOAPHcgqzjHqKkuEILVZbrSWVX7kPoCGpZriFGLmjs
+dpu/+UzXounHJJDD//c3S43vTT/x4apYxw2OwsNCsGT2F8DnSgHn45ypcqgavZw32WROYgKKBw7
CvM7v3Gf7pfzhpEFrpcfg1Kzl3sc7784UpzZl+Ukv7D0QfieS1svGlFReNBgBzLKf+Ob2Zz7N8nw
gz22WXG3Xkkg4KriP7y+v+6CcrOkT/LWaBqJwCGz6azNMwW6fwQVFCGcK21hqg1eFwHDz0tawUx7
FEDgTg+qoEh6cmbRpHk2DV0QKOuTq3bOkGMn3A8fzAKWyEbewhy6ZR0aNOUvY0ueGC9FusGYgPIU
bbisQB7NOncvkGDCVa70vIhNV+kcqDS22TO8MKDBgsbgS6x4uJHrxQEN3pw7985VaIOs9j4Pvj1b
aJFgF3k3yBSD2f/sYAB1SC8pSonNqrBWPu92oCWhknqBpGe4cpBofqqNBNtg0zl93wwMeOZKUNvD
zPOza/2//mXnOnbT2RtqSv0Ev8elMrRc6shion8q9gBDP+AnXBwZulDg/XQitN3B0AD6U2GMAZ2v
xyL0MGrwJx0LgORbr6EMpOxg++Xvneub1izPiVxNxZtI3NtTyhf14+1m6uLkpK6FExO/qd7ISSJ5
VwsDRfdzqyK8jWP7IDUdVSR9mN/ZhSpq5kvLsgBt4YS93QReHnaKLO2YeRWheMi0UcBoPcuC1N4M
yddt1nc+ZNe8s+qNmK0xlBSgyuLzgKZFa1R0IqEweAzsj/R2jbgCx5CENcCUv2FTteLtqWA7Bv2M
zFhVcbceqW8mIhmfqfJUaHMSfA2uhtrryMLUO6S3nZbd/iCV/KbdA+ahUGtMWeE/X3hFWOC1bC0r
roiHeM9xRkKWKeL0qS4YUYCDhnrLx2iQCiYEvzxPkRQ1LB5XzqfjpidhvP3uJ7JWw3XWpWDenuzE
PMvI/v9hg5J7j2CffMJ1Vx4USsj0ez8hqqErD9JAi6bJP63frKjRKMrk8o6meI6fN341pWo9Uha8
WBTFrh4uyhRH0A+xcKM3/0ol5WL/DqBZd66KHoWh3oyNlLeB/9qMb9jSoWkxyUFXptzrD9+EVV8L
CYyJb36120m4kBNaz20LfqnW1jiKTJhUknhx/23IRtyxVK+SswwzrBhxbPMZraSWFHkkCD7iqzsd
cr58uXXk0BT3Ov58twZiwLmJfnWSY9lwzZOFKcygxzQwEaAZxHJLbmTWTznw/8LM0dLzqZDFOkV1
L9Zy6TYa3F+OJOKMnZXUj7C5payI70veYMKOYpw8RATRsbzh+zrgSgZv6sXw6AAfkl/OldPw0Esm
BSGWamg8GuWAadnQ9sqJUVX6nKcvaAIUEQ0/9aT5jiIdgh8YOBCuW5+6F2EYFPgrvVXNpmQNd7vz
I9QJ/CNMPeXqWJpbbEH1aw3ktgjmhvuxppqxNv28d5GR8IfBmcsIoy84zVwJ49jQRIgJN87KTdM/
Dget8fDADGRat09H9T2CRBBfPfCU4+ikhMWmSBIQI6XjuyqUWPkiAOm+i55bLYc4AzjA4A5wkNng
K2+QpmBmIe4We9JIfMP3cJlk9tInPT+QMueLQPuo4n390kmrRj7iOsfHKhq/PUebpjdBlL4TQk2v
TSTXd5yc/AfIZLHfBx8QlZh23xHOlxYpvG1MAdZCwCN7k6/KClsCyyT7ENBAQeyagUtQmG/2ksDX
5Ovkl7wLrqocT9XzTNJLlR3Sp6CvuaxcLnQVMjBcDRzGQtxHkitP4o554is9mcJNFj0TMahK9rD5
+32M8loZ+4iZUcJaAUqv0DmJDaUAj0ft0t0xMoqUEsQ6SktBBCtCs4ge9dkDdun7B4Ikb/nXn0Kx
U9+b+2g/4+XjuKzOc2ojjCnkh27AnfLcc5t65lypGPsVljxs3wgQ7noIXVy8TZu/ghj0J8oiYOro
pvbRwFZPNJzNmwqNoWWZo8VyRCs7MBbdMIDpNhhVs9O2ANHUZxKlmzRcAYY8HcPCcRs3g2JXywTs
xf05CvgDJZ27fIiH+1qqc3r2tOpHJSFi54ecBe3a9Fkg4eGPFTEDpmwTr9jXPCjib8LstG/TDmFw
ajLvhHC/PL29KfnRpMk3JeDfTMoeua3f7NLwkhoe2ciBhGhNAwI5nYAECQbX/RjYWcTVDbk7QYBk
t9ygrE7LFAdkJa6abB6OJ83ZYkTDloh1s/gu8spUjvwcoTzaE/TdMis/4nUg/YXZSXP5N6o4DvpA
M/VmfINw0yU5bH9mzJ+ERVLDLIJPHmVgBVA0pPgZUT56WSgOM0kpBobZR1CYU0S4tbnC42ziDBzE
31HEZuPLohgXcXWE1KBFee9Bab8tdj5pGv4+QAgdwpiOPmKrSBcfRZkF9VGccVv+2LTThqLb8Tvq
7vtsF2aHH1Nz0Ud0hzxwJZHjUlOFGHugnlgeMoImTB+JLyiFnuQIMDJtiuReWPCVwSwIEnIj1Iud
88ulbbqMl9552ady7CPpbxSt7TkecAz6YGIESHWKig06S+sOE+Vw+V5JJHKbsM2cRyVibzOha3DR
BGOSxaFAkuocRc2clGg2r1EqrgJ1bHb8+NLLHn7qj6uCMfad2in3ZVNoNsp2JclD2o2TibEFzrZJ
laKUZr+4GevvGBE2YRamkuc8zyw/T21wH3D+08hhp1oSGBl14idpfcMCfnBjdVOcU11orYeYAyGq
/w3IVtNBmZgdjxwRvH9Wba56tzymk/9o9vgY9mIZF37S/fXuZP2Ynq3+fmhIbigv9ABr6eJVRP7B
c+HQHuLuxu04SDjQ7mpGHaWTPYkO0geZgGc4GBpadMob5rbyZ3HbhvuR9mKl8cy+QtSgB0r99OjY
SK2Tjas9hGdk3X/pgT54wpOWlx1mV1JIFjYDNqpDivFNlEjOBj961GYR/YoKgsazQ2+Qp/NlicSD
W5Z7W3cZ2W3t6+bzWSVe4/RG5bqsAlmTMLncsBo2x0PmBAY5m+Fq1LSWlMa3Rnl8GWlljtUsvZBs
K/+m0v7u8Wy9MuUBdpsLP1S/oCM0CMNZL42D4vDFd9Pj23IWiqye3s7iULIRLjNL3KBTJL6MOTpy
HLJWWuzebMson2msVMxsPQs3z1BKhT34ya3WzeVish9QsHLG5wwCUeToGcRLZ8bYTQiWIecbsKvi
5614631P0q2OCDi9HU9LWTlE6EnBlKN85/sY9GuWSrEawfhvVDRrUH9Z5zdCx0hp6X/xJSOGT7vq
1uFHS5iP4hZiE3DcrJ4TLKVG1nZNga9p8srhWNiytEZAvSe7/ZQkGs7TDiGY5AxTSyfLmP7no8xA
zCOdgFypYuPWaDqPHbbecYGkpM14TtGUasTNaVaNWZDjHdXHQOZWLuSLof37xcwAM+pghGOS9KqZ
6BpMcgeS6GrtqrcmFR09eJFm86hJr7giXVj3O9BjB+hM2xQROzjgOu7uOrp6VQdleVzDvSLwywHg
glc0N2KzA0M9qrUDZBFv6igvtYfks1Fc/bf6ciKWKpsB9Dpbg1EaE0X/WYvxWaCVa+vGEZn4HIAg
0SjzsfxBGEp0ECvOc5EUkmD1BmZZ49mOS7zJnLBjS+nmVSvGtJodl3PcAaHlaEl2vkqvrJmm3+IV
ehgW+UHA4ZT3gRiZiT+1es10m+6CBn9DKksXFQa1CYwvsr9JrKXe5RW8UfOqdOsrD79V+SKQ3zO1
Jk2SggDEaHYM6zo1IXpz0ojxuDG+mbgeKENp+YKbdABSSXsyMq/7n0QUkvzToaPZwmTTBIwVDpsQ
8IlaZ0rmJWiB7kOJQ7NVEXdUAElAtUIcXnTwQs9uA8kQtitNELp7LE+DCBmS5NFEakahaBmIeT+Q
a/xPW94Ggl9739fHPFYDgfKjR0Klxgegc1CIkTbToFiKXUwnVvkkHJd+tmHNZz/J3dPJlBoKuj9e
jDuLfWBIvQjpdOYLxI36jXR9jNyySEMGK/JDYkq/iersJH8EUYQVU5jFB28K9fRfP3gKtANqHIwU
R6p6Pkth6qtosdYDEUQZ0giSlYgu8vAKVUgkoyMat03lbQ3swLMmtjhhZFaZncyYJEDFHWMxL6dQ
ZwmhA7IOSobb2bj0iX8HSKuygVvjOx55WofdMoWkLdKj9qh1p4Ug9pvPgMtcGqPMEt98PoLFSsS0
B5hekO8lDCBiIEE0DZx2upY7SG6/c/ipJi5OKEcLJX4LS7nGerjq1b44O7ra6zgs2m91CUdtzRfp
m0xj73096XNHhJLu8Kyc5sYQDelXm0OOBZBFzBYnsi/SZ27msmKEHyobjDFRZriJ53x4T/nud8ww
1K/zU+7riW+TJsiZU7CwMat2xqVUYn6UMoGaOIB24oL7rcwx62bpX7mteDQkA4NxZi5MlEHrt5WC
UQTcscQOZl7gWiy2FfkkZraQRIkqCoJ8dzns7Yt8x7fvsaGwRw2QL9hqlc7+5QYvD3SDjEqOEJr3
qKfyXsN+EmDYccpP/kGypf5MhyBMYka39EB1fM1JqeKyYYDMzABLlIYyhep877rWVVcKWBv+7wes
Hw+bbv/ROh9MPY5Y6naQKuVE9IneybVoXJJSbZw+9qxvjK6vSEX7cAEU7dXrECvtt8WZFH0gN00H
A5hGPNxsVuX1+DXxNxAccKqf9mBlWl7TLaIysLBTMpvV0VIs8tKW4kx5Hkf2uLUFwAJg2mUvKpRB
g4+xAkNNrvpnpsN9uHGqzu9KPRDjUrsRK1SMbGjoIr2kLipL6j7hIdXXcaxbnkajpQLoriWCCQ5/
CIUjOhbB0q9JTuVgCoUAEInS9YYvxnJb93ii932RHF/2rijdMy1H8yV6eFAtPV1X0saLvwwqVb/Q
2Lh8o86tBn3YDEuUoOp4u5y43vG5M8AV7/UYCdMzuDHIH89inv6XrjGxxWnm5K+8P4ZaCClYv/5z
8+WO5anWFQkLIvxBT/n6fjcW4yymsaZk1oiqMhjN6WZUnkEjYstftxmYaOSd/yt6UBUz+MEi+Z33
cWHELVggA3P5oMC2IqNCoFbGvv7daT6tS2X4AfgaOZGowdE+z5Ios0uJW6ARP1W17q5IJU3TPODC
PzTzoQxtXKv/cwdcozbpXOOixsjgbW4XgW4VNPrH/WiF0ju+7ayQUtFrtDUs6vnMW/q7WG9JpzmI
xLd174bMiHQ0E23x6GhU5GOl1M7nBQ9CeZzib4yopdWWa6ILezYVjS/jhouxMoOx3a5GiJAlp07G
wczlmK1d292MLb2ZMbbrE7JmxfD21K9NyZWm54MtBVX/hHUjtOG7YcW4AQWUvcMqw6JYJt9V6+oE
XOUY4itAoCcfsjs2G6VTBgh3fOIcPjcG4VOZMcLVG18gqvDB0r+AjznsTEBrDZyvQKgokB57uGNL
6Iqr7eQLGb6aOWDCB8ufKcb9+vKV+TOKcG2jN3KVTh8JRU8azIdPIZhi+DYUQM8NAYpS/6qji6Kl
xviSCH8AGxgWP4pitRkGeCGTM530tou0czlz/1lOVpKMWOEHyQlrGWpxHsgiQzB3YmLf1zvuCEaf
pUBF+2+ZBH+nla1teydu7Wc85IhJqwEljbKqgoMWGJfw++PU0dMWoUFa+Yw34sEWHVxGNx2wkqCd
BPbzs93JTgFGlHenNuYB12vywPz2CSIewMGMZ7oNWl+j6lTw8HX/9UKTg6L+16fDCvlpdC53syqT
OcQxWPO16J8aZd67LKsLmHI1nKsnkvHkN+hCzdQeQyhdl4kK2so8aNcFWhs0yKoMCa3i8AVmpLWZ
PGKIUyZLADI/oDTjbyhb4jjzVChhvMnxqlX27+mWdNVJf3FyvS0yXNbngGyBAPZabwiVw3GoRAhr
+Z2GJWUL8uVVkqBFTePuI+e5QzhVdQ5cKUJSXHbh2Roeeh6nl/BfP1BNibr30k7VoNV4qz9ZOIEi
Z1ZL+wqKu5kPsv0z80rLWOEKKKjhgTMdMTxqfVGLldRMcwM98+kwHuSn+lYONfBsMGE8msJVHCr9
2J62geKuhTfGKwHKP6jLEXpspdNvdoH2t6xYQiRxIgFi3DrPMa+iXPVFN41OTmKsaQl+OQhE4kb5
Wk0MBKZ6hf1sfbhRPzmLoTNKiRRtLmbG9q5h6wIzRXQ8SKOIQ3SAqdNwnXh4gkM52Jy1KoFVBh/P
mFdz2ASuxXSqsWE8WX59w5L9cV6FoGc5r8UvI+Atr3T+XeR1v2BXyCoq2qLOFD9N0FluAdaz4LeT
cmme106l1HPRUQHVCEebMEe4ZXXD54p3FnyMgvBLzRxlMpz8yJ7osTS54BBXP9LWWuSKt+U67R7h
IM3U0lWs3kL3uCrJvCpOv48e+yg/qx7EAunXZN9/sN7KlgwQC3GOwYsVMEm5buu7rK5kHHgZAl4R
CkcDmsfPMZUeSpU7kBDgN0TKeq5/b9Cd0h/dYj9t5vmKMnktdAj08RI/I050TT6lVwXN1I50OFAG
9MN9G8WdA7S7uT+pVH3wXmBC0hLh+2sOuJNxejyY6cOtoCT5GnUEZ80HOj0o5hIMyBBq8yDra+08
Jk1/NDkCZGC4cXejFPfb8+YEY4bDo18hAyy3+RqB5hrZkgyigGpk2qdZgkb8fAplrTy3v4ySWbQx
V2LFO50Wx/t2AfR57lNy8OZcaV3STtDeRW3kj8kzAp6NFwh+mcUiLP5krNsLVBVjIEepI9l2JBnw
T3bJcjv3CkuTBiq0zBrPNDqqhCre5PFNgediYh9HhR0itO9qkT48Tv4O9wrmB9Y/U6arbqsVEyQ6
1Gm7ivfvQ3AR63msHXl4crI0jqPCiKWbVvRxDH9lnvH84mJpVneC07CXsJgICX7BgskzcJ/ssUA/
2W8TVquT1Wx/FWf6F2kZPSDKQ0KJfZEkoawZYLD6NJBRW5g8L+u+ZrlVOqEoq0SN4Nu+3RLifHDZ
GO90Vfbw1LQbCfYjIiOGySFZ1I2kyRpviAIeQyTEgb9dcyiGQpqPTao+gmL+/vGhk5Rf3nEiQKxX
V6LbXuBYb84CiaqcuZB1zW1FxEqoVsmEKgy80g3TIwzgABT8Nd13phgBUrObUWOY8v2rwlUGuJg7
RoJLRlCPFF7R2iGwnjlr7j4b6d2sNzsU5rbBelTNRHracxaaeBno9WC6kqpKN7+Ae067uMBcaLHi
aCPokeFJklWOaOGpp/BgmVWIpTyFjRqo7BkwSdRg/SSL1uL9og/0Qa4uLizFvnfVBfdtGun/D275
C60cNR+zvdchHvNp3HErsLJ4hY1kaTPuppyDwCIYHZ6cMnWrWJ1i9qx2NSi0+ttOrUmxU/JkL5L1
JD25/X2XrjVAVhFvy+EfwlfIXbmgsflr55CwAXGVYJFGvwMCI7JLJ1DGPSveUSxOnDtfsfAX4fYv
3G/rRUf6MyFdEqQM3+PCArxaTJgBkWHJtVZf5cZzHHZKpo9mbGtjg+Ou+hy0Ar0jqPpSfOhtSSte
54JCtqv1kY58YA0VIQpzxzJzAaJ/wqpd+AVIuBKKGHWC3YaZu5QT4BQbWgRnLXBxuTAQeYlHliES
bz+6bcTg/p8DKl3/lEFJ/QGVL1YjZVccG67IN6Pih1y4Obup6ASjbuAk6jUz5WmkpBY2YE+EwD3Z
+XpBgbeubbPhC5NVQ/ybs3f/ztv/J5S5hlvPewv8+XWXN/5sltx0Emm/XVdtdtbjgC4qBfayZPL0
9QTQOEh7mdym8Uu5rZyXhznEbAxu7DbJYC7Uw4kZrow2uKDK5vRzrUfd62Quy9S2KhgaeXXhN/CC
7aIqynEdfmt4xJkF/lUVoDpaNxncZD7PMw8EP+aH6lWFg+ub8Ho2IiYo9hG1h9Nj5AACpHvR25Ax
hfrFe8rT8nLl/KccBdpaTizJUyiPVYOPzUcHuS8p8IaDXUmkVMS29kqBotfskpjmAUeYH8u/ubPi
D/2TLH98yiIXcpn02FtuVo+A3/FtuYjcxn2tBR6boXKbt4AY5ZANrgf9tdXuzkuhsLN1PfAW/ebt
1XSC9NMrCZCKV5XhpXYuTGjtp9kRBT7RB5LpCGiQWdcLxUpJQsDGU75OMFNpDh3Kd8LOrM0AA6nj
znPsgoYzxKAEZHS51nQDNfLFR0ol5QDWu19g+YjPKi5NqyvQ28GaCXxFNx8AiWjKqoj+c48v2OF1
uhgbmUXI/+U1gJQqvm6CbiBBjvcvbwSypL2eU6hBd+SvoU7QnDKC++gdTbwmKZz4h8UrJzOeEfdH
dNrJ622x0qupid3GkkUpctwoI/dKozjhXXQdRS2fC5BmB1GzcK6ub0+LKIkDjnl8esGtV/+SLoxL
t+PsIWKh0qw3pzBjTupia5qizqI/pe9vGsPbdEqlhxhnMtnkZSy/z560iz2HEvhDlZfnty4/cgaj
Fs7k7efYC3eerRnyxUPSiIj2pp30/lP7UQ1sHusBGq6XwEo87jZlkC7TXsPQOyIXAf4rSUiDZQN+
vUIZzT8oCPIi3QovWFHjznTRIbWv5aez7Q3i8g1S8PrnKKWMUM23Y1S4nPH1BjqUsJPxP6wXau7m
nbZ6IuYM6e75BViuRKC/tQLoWAgE9j9z15vuLPi4qPUz1uRHG0qt2D+8HAb1vDScWMmWcKpBv8rL
VD1L5oaHRDhd5PIlNBgRON2fyOpAwSWrJ0Z0l/snJtG+LSGkdkPkP60UMJd7zM51zXjimwYXD69Y
k53UMgzMEoUMRPnxRcLFqsAr3NiDncDTMRqu4Y+m6B6p/7Hslep0uo01GT9F8I7X8nxDRtDTl35p
yReupry6UkMWMM7ODiqR3L9G0xH3QWS6lkE7DI4gx1UpwUuGGrcw2scvBod9LjDg6FjF72EgaLP2
yK94Mvy68Sb8PQi6RWYgzQPePULRBbO8R6esGdQAz/JrKfhXZDEVtcAiN7Z7k+h8uTVh+BKHYvA6
p7AoCvzKWHCuxFIPDl+o8YWAu0IONAAs5TXOXuE8OITZn+9BfQUxiDWa3Ixl3XhnmOjboaKxL9Fd
kLyqeJ8wBlvy0ExEdTqHt7He+F0KfhLi3jleZOgcEXI739fFlzUQ8G7JFF9TjqwfxTU4zDw5Gf/n
koLLSJeh1S7qYwmGVIdp2saPZfeOnear/f3TEvnVcK0G97MoD5tuYYMl8hbh1FHlSeRKmgh76c5W
RGGwuQicpNiC1LavpmR5MpvJ7WrpYNuW1bfv0hJUHYySzONGlrfVezggNXfeS8/aF3UmqEbIia2C
cmY4M0Y1WSbB/Qr2lbFdA3wUs1n/rnVG25y7/KuI0MC309KKy71aKnDSwtWAzNAAjFaLDEe/9a7/
/DfJFcM16Tp3kX3od/ifzQkNaJYzJDpb2q3Et9iagCL1LZP/F5TwkWbG9LLEOSIhZcBSdqK7584H
OGFM97kDmaE9xq//erxIyZOIwYX8YOJpeUF2tssYMGo9D0b6xDZsUc0E2VjFbNl4RNtGwuE3zIT4
1rHlKML3yal1A023pSIy6Paxs5k/vlooJzaHcToyKr+/jJZQ1DTHb/RVm3saiJqlrqEEQgby6ohh
aiI2MByMhaWYdqp6JjO7I9/l9mbyguOOUh2v/gYdItsI4oPXwOpX85VZTBhhoaJP2LfcF3hr5Cpo
uRldpzPr13Ksnuwjqrf2DtbHI4lgegTPJAha12RUxGDXLGKto4Gi6J5itWzNghZQksOP1FkdyvoL
ZVECEW/8LciUuvSBbQ+Zdx8PuMdyb4jLUUgnO2KKp5n+T4G5FkES6f68ZEz90XJGk2VlQzdEZdcF
W0FpOencVKpOqzLoiJJ0jo+Opz66rfbyF8OWQQQN6jwa1pUwHy8YxGzbpRlyWxWOd8uBvfaQJFJe
78kbRYHOrjZUkReJXv5lpN0Ues8y4mzmB5GbHTEaiOqSvvPTVxNGnS2AFDta2l85o5xJCfhFR5Nb
df/GzPivyoY4QMi4pFRjPiSolZCxv+nCBx+3LEu0vDFSEygUtj+VfejtXoVlndhySOvhHkOvKACt
UnJKM7iIATrvY5vWSQo09NiJzS4uHHPZusvMlT15OR3W/4cgsy+CAZ7wTjIuWd+Db6GuRRLvL+i+
cbHQXi+cwGclLJ5nzGko5/FDLUfMZAqTxTJZ+wY1aeRxuybjc5ReaoHWr3fLdYCOEobDCon0EMS5
RA1a0Xb+v38Z0raH0gLSsp9Ic1HMVyc+SNzlqxeWUcvH6LT+6RJ0e4//JtVKaR/Aqjmm0H1m/9kE
w6RiOTcYUjX833ASPtxxGoVIYyJFbeAJFfF4Nsbmi44phyOJ0+qCm1RyWssmZ7jCTRCxZnWrc+Kf
whpLM68xuwo0YRuRr9nURvdqwJFTaFKye4PRz6VDkyL3N7XLuI2lHnm6sfZ//Bfv3fwzm+XaGEfM
9xz0xN4+Fiis+ThKOeNICzCGbmEBJKf58B8bX0td7dfaMvIOC51vOc+mzfkxW4gF2gQYVqhJwW+M
jV+G80S/9WzS4HhPqtfpUql4oz/dEs4nVaxtTVn7/RfJpwBiGSqJJcksPmSCFGYsK9HDfd96Zvld
Q3XfG78U/RcKTUusO9tITdmXj56XvZ95tj815i016vH/4A2T5TknTu+pV5+ilY1zv3Q+z+NHYrl/
AFLyItja+j/nVVzKHiXRUa2IHMpSn52OR9/3u/t+D9/dtD1ZUg9Xw5mivVqJrsvTq13WB5o11dHm
XrcLECHryTPFQmp/QEDvDVv7RVqb3e9F+weBNgKRtM+Mjlp8u5VaqRB+mLTcSkUU+mm7/CDIw42m
n3hTxHJILFLqDjCC958Lj1NkcNTry32rrByI8Jw0A8d2dwNJcIBmy7VxpU/SuO2qswjSUmC4ApDD
KZfjrvySj/KEhZDs2HGb1RWE5DRyjO2UZD/zRaloZzMv28wBdTZ+ZleT/Yqm03aJtqSe9l7nNmFP
40SnTSFvztzgEdzIdtrRUrY02/WYJjMYMdmA81cM75CsLab5rWvZ68YMdo5WxpNmZWNgdXGsBr9Z
NVUUCSa3uk71/+/ECgFf1F7+nWGg3YLfykL71nbyeeT7+aKT8nVGxV/e58IEK23ZKIN/Yoj2yjK6
LjoRvNqv1Twx/cIpQn8/C2nvN5ctjfQ53508K1MAsLRA/iphLyN8v3i6F+u+c4JQuALfJ8CHIDUT
ynHEMue8vN+lhQxJXKS8Fru3O0JVAwNDH67Ygzw1W31e8xnDXSg1Crn3kIT1JxgeT0Q4qkJT6yQ6
HamgXuhJacxWSRH25SA373+2e+cv/pO8OC3mVetuNgArYm8RRlZAxGKtSeShUnkRKCed7JprC8MZ
5vJS+JtiRFhQ+UO963CYN0zeBv66EUDpQ8Qd23ArMNDZtQSALnitelDIOtVxRfvALuQPR+8VDJzZ
Furmcck9TLe/sD9p/qdqViIAhe5cDoUcb534GUiMPMknO1KjDMCHTEipXy7QN6j7ADI2tJEaUkN0
mEKSi+ANFicv2k+i99w+94/piyViFiZ6hQooIgRt0O89bYjenjP4+iPzMyhhyUf2ZNgyvFnJ5znV
nVny3VaNjN4bQk+MqT59YIMfqXpIqKc77Gml7WrPqkCrB7icH9gMjWHdNFMI3n/a8T4fHCYDEznz
/QCX65Jv9GM5G2LeQG5/Q3Fi5NH/0wPIicL8Lami45LF5lkOBULPJ0M07R9eNRorrci8xfbu/3It
ZJev6ldaC8jMXxQzQ8XTlbYFP8D4dNxNFy14Er1ZD8b7HBIryE7IbXfDKDDopn5ru4CPZOhpRka+
7pFghxkBp4EEZ9kzLqJ/gW2u8FOERrIwYaP+A7ZD5+nwuzcQb8XvmWm8IgIpWyMPbKLkFnMw05VY
FYKP3ezf1PJvPy7Yk1XtYl33F+/LRm/rXT5Q8+eqkzpulr2mB9vqBzXMqLWLjiDyloPjv/HqhjzX
nvfeN27Xjnhg3Q1820i0rRMONcf5yVr7O+eORggL9GL+jYZ1Q0IttWUCbWc4pqB4RZjpMCRvXa7l
PVw8Gl3PVWgsyhtunqgsuycYCYBkOmcio2d3WpwYG1L/DzEAm4XrJ5WiR1YyKJDPfb5iVGfRlHna
36ThGff2VOsphslHJpStXPIwWSyHmagmCEfJ6avpbscIP6z7daJZng5PAFprzPIqCXjzAiMSEHjI
+B5lpBPeCDRN+tIwuCpXUTm1rROcVTHA8VAREF/1/Ugi0KyyZrn3126C82sGGEARHdo2iNOkQ8e5
zQ7EvxW92/VlG9RXWLVEoPXu9+dG19imqhUwPsvKg6xI9vI60IEAdkzDikYF/Rw+5Fbr/+w8UA0U
8tn8Z++OQvrjYY43ei8eU6IviET9LblHbHspkNxwdBZDM93yfR2JQjm9cDD8mI0/LzJe/iDULP5d
lkELO27Mg0ZhvGecY4x5x1SnYzf6NmueJVG8DwmRBhmGjjG4e8jh6HB/RIajmBfogQF/vrVEfKcB
ALxtUEJjgmAScnGI96M0J/rn4O2lxtYuVKrjyTbusMX/uv34ClO5bOcanyJ+hKBN4tkB/QF0VAn/
/XbrVrNmnYNKnl4GEnFTfQfPQUbOaWP6q0eKIc9eO3CH0zxsc6JESwfKtEf947I5cY2+P3FTB3k8
VE4tsX0pLiCVDgGEjcRYzPZM6fpgA4zGgyWCa/Rh0xL5ECRPqRo1m1NSg7T7PDAh82STaKap/vCr
FuxxvmFJKRaImp7ekGt045rd7aXkg4rqBznpllIPd7r6+uDnB6dTUwUHDGbRil14App1kq/xGz/o
thHN+6zkG4+J9cpO4O/DtZf6t+NoAOw9xdAQbvOjXDR1SdBWDWOPkWCTX3pG6Dw6GA8I+5N/yqVc
n9KYCWtF4cqLeFoo4bJsRwLZS8x5oqlVL8n/wMBYUHFE7FC8puDOe06btRR3CbUDz9Ui5iWoa15V
JYlp1edy5PZeTQRbvK7lly2ssFjQXhbF6+hBzgiLK2GZE7g4KmU7Zdfb0oTnR/gTF9tHS54xVokC
+uf6YR2zn4OqO8sg8iObTWsnMHKBRxK6kR6J2qwVwMmKUACiTHV0CnTUqPNagNANuxHV/adoWMI/
/i069LI5R3rYKtg7PEGa5uHYbiVDL2JmlZYaidtsBOBH9T15gSlcPCYvEHMbs9SieJ+GWmQ9W2yp
SkSIbjkWNQbXnIwaK8QnnbxDnHoIZj+zxSoqnXjnmRlnsBvteva1azBcR+RNEQSwIop0fvfjrWVt
brbtbm6cvUjX6VvnxLQvp0vsaIOAwA6PxkEQV/S0nNI7KXAGZbLNNqTQdG3LrIQ6NVH33dV67L2i
b4LZh5uVB/Q3hJ4rY0n2Hv29y+G4YvANKXovw1aA52wZ7j2TqCYkFMJGJ2c0m0uzE7I4nsY+gbmu
7USufoNUB+KryhqU1MOr+hflAZop0OQCM3ik5Ub+3XcDhAGdlAtEeDLDa3pUbCo+W0JuhOjRVoo4
GQk4EAifuBDVjszMiHmWLSnMmlpcIPPb2PDIO5Gz078Serg0VfC9PXKEf+JKRgOA+ttL9a7M0S73
l23W6s47o590Spe3y66xvJC7z713UyY8pczetrv8BwdkUAKfF5KaZ85FL6xIt1DVeyKDUif5K+Ht
ng0gWdNZITziyAG0WEeQOc52wv8s5aMkZeV0yFvCb0X5Evhg0kLQpZPn91cKu/bgpucFGROY/1B2
5KMb7twbT2JEneG9mIek2kH/iNqSjVgBkiSHVdASRT8ArOSFoWCxRVvewzjyCia11KG3paHWS3xl
jSO4bBOieo32MLWypWlgXie8mSfBHcmYfOxhvgAI8+YngHGJxIPgQTXZ8UOZ0SFxcUgyBTEKK0l/
+ZDenGd3M03/8L7kRvFmxdMuNOwF40zrp2ZEg7NSvWiPa+geNpYQTMJyiMrDExLdFIHjgqoIy1U/
BAcDTPr4/+FU0Y2OsDvAIAwiFJBtze7N1ABa5WWJcL9sHFq4NxvO/xWU2DSUd06+nDWEsK1Ru1D6
Las5gqbzxhkuTrUBYyW2i+0fRknyGK9HqEkpxpPPuGzek9QeQY/7fxVqqqtmtZxh5gwNg4zbU6CS
DCkup0YTRjlDs32qAld0k8iWGZRwSNaTGn4dPMUTdXfnuuAlxdmiDC33PA6jKLF8sQamX/ZUSr6X
GomrAbvumHcsDOPJhumljAB3Pkvw+o8qpg/MdjOFv7M9C3ms7RvEYoR72VqbW+Km41n5o6smQuUC
u4i+E/maBj/Hyel5HmFwWrWX50Lx2nzdRPhddkgVQ/4tTgn7C7HlhYGKIpR+65lVmJ07MfYpiYgq
uMkVufUc19dB8H2VFiusuP5IFoFjTsWzB60myzZARgLHbv+UWXUg26VBj8o98AvzAL/w8iCnMqTu
ghh/mUnfJ0fSX3HB+f69YdWfNqBbiT6VFD+Wnw+nrX3Uc6BTSwt8XSizdvIUNWrPfwdHDyDvih5I
eNikLpqWr1fv/qyStJidE1acX+I07tgb0my4WL9e031bcRrmtyuVt2y5SvkQ2rhpyGAj7ayPnmAY
48yA7PT4DrQ3NAtxt9oY/nIzFgzwq0YxSavnqtu11bGEwCpe6+e3HiAIyfDHEyMQt6iZ6DKiOIjy
TmB5gY9QS5UhmIZq1V1mga3xnLUKMWDbVRoTk3kJ674YirQg0U166UmpYCGLDQrhO2ZNl97SS9kv
+4R+RNrUw4yxW1SP5qeMadaKXzKcUTBAZJikjNIlt5+2Ot1SGCukpk6MiJYWdvvNo5I/XgM21P72
EV4DhlV+WA9tIf4hzkcU7pEvWXBddyyHxZ7+j1T4dQdK/xG/XzybT+nYC1CuPefbHVkc6Rvc5HPl
uM/ck3G4IJOcgeUua1/ULafbflvOhvwL2ExJsWh8rXkuwo+b56hLdivtSv/hM9A5vXkgwxQEvTst
FqF8retLvk2qXkUTOpQmg/94/SouJmGXjTiKttl7OdaNOeVZWd1rp4KvQmA+zVMGij7T6i3lIZe/
6qlfEqsrmoGQXhWK0+KpbwLDHHkAfn0zeiTy5S3/c+rhanCKql0k25nRNJV+tiACmGkChlBpmey9
VcVL9oh4fSRY05uWeDmUnZos+usxFVQgs3i3g/cSdbGbC6F9d13EFhGESSEuJ5kx8P9Qiyn5V49d
o6iO/qpPHZNAa3xxI7Vu92iq+jPFoAqP42DJveweCjuvUxDPIMkLJu+3ySlg1FwtENzM7xNX5T02
Nz8llAp8DZ4RRpCEevqgas0YXetQxSlxibQgrG7A/U0tsAg94Tr1t+lTR9WPMMbQtVI211+ayg5N
mLNECbWoKT+rU8h111XEMLF//kPrVlA42poh8ebwsUc2HaSsGEZhCng29H0cTvFj6KYmBhND8C0O
31AS381fMp/Trtjwp3vFZ6X6AUO+b3VgYNqtphffq4sho9Vvh4HPRXkE3SeKvwMrIe42OwVGiFzu
WiFkaFCGxZDDJmRxMDOX+UODP4X1LuDBw2qCT/JuVWOQ+3xbY3YODGpuLsMQsz203tP0foMlEOET
cTPWQQZ0mplTm+Xr79p30m8pdrp6Qx7xZGkEF4H8c8aBeYgY+yMa3cxBc/TjEoRBrbPMUJq/tj6c
mF4GB0ONlxXrrmrSB1jBAeSg/zwulcYHRsio56JMLsix2FvFcmji+Mu+iwSP39vJlIW4fk+LxYwn
bju+kAtEl29X4GddyjkpLcCAT9HtbcElBH159+0Vf7JGyUlq8nfF9NgvKh53i9NP/GhfbXruShIq
yCNujHeFRfK1vsyA65T9Y2am3/jCaiIjfFyTUoYe8nHu8kvAJwRaI0vc6XmUAPrBgLZqdaMJpIfz
v5iL3/BTcfdohUXufvgzac3Sp/GnzFx4tiEntWF3z1eyqvKLOzF78Ok0S3/VwHXN/Pr9m39cF3NQ
sIRZ4BQsZQIUx4XDUh1psaIyKwEV9wcS8ajxVtCCm8cQaJl+91o5aWld501Wpfv3U2+5/3anQOqK
6vU+nbDThRwu0aK3WX9YLmhLek9d2qnTT3wn1eQfUVRfsLTYDmc+/6igHSep5xj6VZBw9mEoEiZ7
OZ4cjfMnLUSIib7gDPttBhIYlF2TLL0g2eYP0/mC9HJVVT1BNQvPew/KqGmfs/oaM6HLMhds//AL
sfSMkdCTihszBuTaPJ5X3T+yuOcY/5glyxzcRD4SaJccf62g36D94dG/rnVbZWpF9cYmvETmDlxJ
MT/MhpqnHYnp3t62mY5R9Cyf28BVhDiHixtNkXfAJiYbRN1W/7PBMUNYLY1H+HaoWFGk9Z8Oa2EZ
xAwMw72K+eusakGz6EVGLJgVmjeE7vVpaJgOtW+Tr5bDMp+om63TEnl98tkPfnjFImKEBsnqAIYx
MU23klGm96yUqGtKp8rrwmmMMno0PhLUDaTT8KZ/lQYD7DMxyql2jBBoGHi8uFqhyaGWPkAk5O70
nvMxGX/srIctvTX2TV1e9nYf06H8LwMw3zrJsWzpgncJaWjn+O4nbDe0ADT9/kfQ2wxoXJoD9W9a
KbrFtbzs1acmG5CYGbokFIFr7WPmQYiBEnC7FoTtj08fypjW+N+8He65MJL83Nvlhg8De+7J0Lhv
SKmdje92rpeO7TkBac4PDrIXvJraRkyBJB+CeasUj4Zu5dgWPpMmcUJF163ol+czFLmqEZUeTAoC
pEh6CAPEGLbBuoHzKJotXjhSvMH6XMhUf9IFnyL27oKJtFdrccSqmzapss24CaYKVgeeetg+BMR0
pwy7b0MCJygD95Jia1g1RRAvcCGFo8Laj+oleMal22xHLsVeaGsqWdTAOKhAwDW64XDR8fN7nnT7
9APgjrKjGFDEhnJQbFfnWLLBoa5lcWgls0XJKVnxZcJ3EnrMRMCG0MMvwFKmJ8UZBRhJCJ2cElH0
qFY72n3wrVUn3VMP8hWZsmq4THQ7i+OCJgorma5yclHR21SSc7TcaGkX4RkrDU/cOt/MRDGhKrwu
YbdJM9bQ4L6p4I8PbilpknGfqZV3bc7v2YAWq6hBgan4q+yj2gUv2B5bn+kwdEco1MMEaz6s6Cn/
5Iea7dEnSeeI7VNXvDCDOGhZK4fdvPGbHVo+Z+X4i98gVAZk74fBb70zu0DInzJ+8kQpoH08VliN
ikYzO199bC+Q5CUm1Xhhyc8zfNKYl9FM5PhSuwgHQeU3dNlogZQQ5umRdHa/tcEk9yQVZlOtJ4q1
Q3k0t1CIWD2J1sxCrKO7SSGws/bk/oYwMoET9TU5sP1PTJHIKyq99DZX2Zmuwk3zIZEV9EBVZgIX
VfnzqDlRCUoUdRe06nW176gKm30/AV3+x7N/3ODoQv1IqBrbGCQOrliGGHCBMnnP28S7kNi8sU9F
TMcaZEvrpbB5325gliQ4sef3X+rjAl7pHkXdguOxyvyX6zA+HMSiOZWMT6TNMUQ+zB13MM36wrKd
jSzyZ57KWSTxmGCWPfDkTVKs8KPnNVvO3jatLNg6eo9GxHwPWn5yA9Doy7sbuL1TtG98agjSdqPQ
24G5v+avKI/JI0IpAjQDy4U5SSCaH0hOQurul0xjkxmPyzd3SQZ3IP/AWcFx+yF+bSA60oZxLCfd
weroEi3pba92x5RQosSrNivxVVj6PjciHywSyZibUhTy998KTLqOpEsOcp4D1t39uLWzAWnLSOq5
M2dpdvhhBR78UfpwwMW+GJNRfCKOiaAGkX85Bg08WJEMJeMvuae3yYhaMjBDyDt+0zJZLI+BfM3t
DwhZVKQcJbFHOxa1vVjICIFGbEXzvEZ1dWg2ZsOLbZe86DosLyCEXAJqh7t5CIe4MiCuO79AtFmz
fn33GRjnD0/eGEi4E0YqT0Wf/RTnpFXX9VrPMIxr+Bj8kC7ps7Cr7QVUjzJkY5CPLimdZoZYlrGu
lC93qduptXAj05UvIljqbc3QRWhlKEBxF7I7i8ur7+OqQzwrWPnh5R2sCEZYXIb+wfNidtdSZfen
LI41fWZ84nw/MAFf7IQ5I44NBslRn6bSqMe9bbHphBT+Ob4QCMwsjBStsE3Us6b6OZWjk9tfnUBt
7RleloPc93MXxPYh5DSZLCyGb+OXFPclb7ekFStYln2rggqrUCAMEfpfrsJr5GJd3ydoyocZKdaM
3p9VMogqALlFhJpLYrOjxP1SNfTgttKfeHlc8Y3STV8KPCga1LIETkGmDQgm7F9Lh3g/DpkT3hbj
mq6eMZgVScJArslbOa8WqQnARLkUCUnb/OlnoLIWgacvacNR00bsDI756OQJtD/u8RjOm8cV9ex+
qzfvHIQUgKnQh2UMZQPt6cGn0jqyA3t7Ro71BBLDLWKf4FKGQT7BJoaPSekGWs9wvrKpY9q+jl9k
LIdJ8RzWJQK8hjuyITpofSDqQaBT3tZsnfAUY3hDv30n0+n35FFjzlJ1sSwKWlpyQsW80mFRSM0s
CorPrVKQDBjqxw8pWFXZsixZAiOWw/JkdrguEStpI81BnyEKAjSPiBDbFzc6L01uqetbGmR1fjFr
ly56FXRLwy3ZPjjCbC7QyHqk8v9bkU5BubNIkw1OflULrNsK1o6tDs62nymHwOQLG47x6RQJYAmo
2t2eGyRx0fskDPgWPgv2H7j4yiDVPyCPCCqcOLeYVfHXbR3Es54ITvKPCnZ2HCYxqQ+pL8cuXeCN
s3gE38lQchpT68yFeKhO+03+Tm+5FgVGFNLSod1hOV16J/BM+ggVqZuS5NvKghkrmJs7tOOrIOAr
RCzGPcgQYRJt1oR20XlFWYeIqnsfpnwmhu41YLBCzf1U0I0iUnnTutCySBDYzVXXvj/pFqSYaKFh
4yoyc58K2EpRbot+wwviysJ3rWzdarQ3t0NAL60MxvTZ8kW8SvmmJt1QUPUwugZzED561ARdpaGg
RWzGt6uZ0HUYth+xYLEs7J0Ofkcpy/2vv71PU3o6XEhAVcUJ0cHv27tMgQ4SJCZx2WVOvtJKI8ht
f88kJIlzS082QUZf6ltnrEvhMrEfX3fc7oKQOpYBezqtuTxvRTy9pT5fcPu2F7DU1+OmctzRdfun
JuK0dU2EYs5yYidxnQdPCTd+B+/zUWXq5SNtXaSkfBSZS1DbcuwSv2OOm2MtdsVDMJ9ub0xwzeHP
ub9NHTnczSZXMyRowN+kPKtZorcRNNyQZSk2v3nWCa4FLrq9q39E3pi7GVIRpfGzwq/pHc6W5nTW
GZlWdxVHnfWT/tpsnWWSXjUKRwF57qfljoFX3V9yClqkK43iG2ZkvuENQKswmTnl4gvEGgRd8UOr
nnu1k+iGE2SXu37h29S9aNvTaZV1hZ1zsvMIpZKjUBfxI26ERdYnuDn+G53OksXj5XNIJcKB62wR
v3HrXP8FvwJgOIX8aMx7ngWYOju7Nn8yRDtIRR+hy5jvmEgUBWRc7MbhQmukzfzgCTcHt7srg9eT
FqLGFqThnOYZfC69DOVbm6hOfzLItdtrTItmkYbCvKVvv4P2Wwc29gMEyjMI6HI4mMjsyFQLF+dP
us5ExgQ8o252MvW3QA60NkuK122G8o/l7KY4ZCd0kLXxOuIFuDBD+9y/n8lzVfov6usN9szM+E3v
Hglx3AjdHtC8BW/TGb1RkbxiPJ864gxfqbyl9zjWDidLL4aPG2eQWKp4ttEtHddKEYLFazz12gDq
H+4QB+0I//EW9moc1uLZPUyxpyiGYkMwA6rUx1iyihyhzuZn0JA9f8fsGK0+B9TKva0tb/KkUd96
4lizd1ksqaKlnj4C7QJnX0GqciUUilns8bqYNqNFfZ5hF1Jx1jVuVq/FLf7jcIWeDLOYFZbLEBQG
Aj1BIGkfJ3U57AGrDPik6QT0GmaQmAyVHDvVqFJ+5ErvOiWR+Ky2tjSeiPaefOS1fXQNU2C50Th7
e5b4mczsV9oBEkJ/1bajV4bhZn2xahnYJSR/zXYZFZ07j94wVfByfbppEEZY0Ut1dYb/vUaSIJfu
9GwAdj++eWo/Oc9JEJuojgotjwRXcwxuW8r8RoLplfQYoG40Iuh6q65xWf/DRwVaz8eFn0Gyng0p
GijHaferrMIn6+REi8gRJT/wDFhnRklZITOOeD1KjPxjwB77m9Mo0HaZhVlIM6xsW3utyKQfSTJD
P++diBRcoQmALgbSsozZJqudAYz+AsGoFChnLaEJnSTrH68Gl97vrLn5Nkp2DrEakAfatTi9TO8K
iOv8vPyUW1IwP9/xmBLpZkn+Fapsl5sAf4stiUw/Nvxg24KGrDIyHMUP3c4B/g11hFrWFMYrVH31
Hv+kU/nW4qzDcv9gWHIBPgg0EI03GTOMZaa9Rdvlj/Kp2y7VGwAB9p0qJTUXz0mZx+yPmDIDfI5E
/HMc5SKIhQ5SDRDK3SA1dznIhu6XitSSRmYIAZ8X2hp70nDqAyU4vCv6S7E64H76rdy2pLGje/I8
cq8QBc1lmh4kHScFkMrfaiW5ruBbQAxtXwzD3ZjLWzgbWFypoDhboBesIObK5cJ81tdKiwDOVC/6
Sd75/8iZgcXKYCWaNXq7uMG7Yqslgoz2roAA2F0gGiuAROSTBKsKm9HG8fk39BYu5a5rp6dT82lD
HFmNBDKepfC4o4X5M7/TAZn4y0cr86y7s0gWu5020KdtrmRVv41aM75oFuw9bxl4CBXE0trcpw/F
b5pNf0qoQJSQK/0YpZgSQDEqTRJcuF9iFZVvze2y9IPT/0WEPKXPYwxneMwoJRqASI9t27pu2T7P
7HCotasI44ducJUkG3oa28DmOYJDdk0O/YPpalrYytALSWvstHApRfvn2S/imBDixKVPm9nawenO
F6mFLeMWCqRsRtZmZJtg/GZOxWtfJNsgX1c65XXwmhJluCyQqt8E4sI6XXEwZqCmMpZJ1bUVk3Qs
EHpnDjMqDaD14YczkhJWo5TC88loIgn76LBn+dzeWCxxBNsjqA4rl7G3HA6hSRUPCvkzrAjHS7zn
Y5Lncn/Mu1z6Wz5KDv3eM6WhqhNbn2U7NEsveSrIG0NS85Z9nW51L7uxhZUG+SCpIz1vhlQandVl
otOUFWggn/XMK4NGceOcow6G3r4a8P4tu2Tz0aM8oQIBrCSHLXcwXVfYZ4sDV78l+pmlYxV+4DqF
OHmN5st06ZBFE56vowZXfMbctX7Tmk1OTF2MO5zlbUcILtx5xCDTVvwGNxcmUtVkE+IECOm8eSwg
a2cA0GyVg18oY2aViqVqQV2NcRx5ATJJxXTFBqDe0YskUtI5mHRWqZcNx+yg7RhG7mmsqMThilkZ
5bRHBKFUK7anCFKG30SbhejglZIrwbHclc1XcGiyEGFv+4pyaokRQjgcQIkwcyUGDux/UsQ/BNXr
0Q2s/BlK8urBg/mUyu3amYEojYtpATXM+/TuJVEcyNxi1//q4LEAZDWUdmGFm5dTxfKoUlzyVDdY
+mUD7PV4G1qS3M5l2ya14MJod0QoXyxW89cGAiUDUyy+jlirV0Gve3Yfy/eko8UF24tEHYRVVuqb
SWJkzPgg9+s2PAvxv+fKz8t5h7iaJuAw9KSFPfxqRMX+jJp7WH7LP5+wTxuQBoClTiMymJw1WUL3
Xd/yjTR8A5dQ8JHPVoIcaW01QVXtXfhxLcDdIYUp3ZguEoXx5zgQcyPHeyZnnbNJiv58a4Zd1yF0
Ct5q7F0Z+px/womrRmsbTuMF2irpIVSyauWc8U+ov9sNHCYxLaamnCb3Wvy7CrWvIabENlcENHkr
4z0XvlqH+prM3KMjSc851P/UPa03bMBxmlK5N8bT0BN17q1wMpDsSYunHeKh0iseqU/5CWb00epl
HWM8b1KDDEQbHLzIMW7B18Hv/8uT7sLYAb1gYc32SZX2fjnDNuzEr6mkiX8xT4mraaENXcN3OEgw
Ja3wEmGqXjPICoruTKlAcZDX19xxKqKo0pFkuN5IePt7JaXc7hiSkSPcQGMS/XuPMfFsMn+dgdTl
3Aku5WiVQEJnFfhCOkvWUBho3df62r8emb/SZ1GLJse7wkbBhX9fy1CINiwk21U7YN+i+CbPeyMT
OKXtbp7f70tt20GhhSMzGhpTUKX49Rar6zBhnU5QlEFwV6BfOCcXMh2/fuh0nTn0I9SWb0AQ4/mg
GK5jLrZsZxMLPXkgqNUHercF8tj+tM9O1SSefxNAJByovIwEXgaZwaHfm6U1Qzzb5176yNRakWPj
g9gnJQ4LAiUVnjL61+ZH4lxcfMUvTuSJq/wnZcWI9pXP20Q8yhfHhLxT5y2gJqzFkeW+s5WlxC3y
qg2J7GuZGWDXYHGTQ/9Ucr8vH6g9fRt/+0ObbCZpwRysLY3KvJQGMnlNEKBhnfXNyVfpcPYOrCcb
F5jYrLxcDbd78b7AHak4LttfQUBcA1Re3sVZoTZrjWF80Kd3Jhd9N0n8sV+3ogf7XEXm9dP1Y5bv
K14PNBR8alOaEi0xeThHFg6tPaZprdgNnDQUpIG7QcfmDyz2cdVAcK0r8VhYhXzm26ZZCIr5VHub
iQYfS1nzubXdqoKyEPBAjt04NV0g7CzcfYUKw/hPzhr5CGdlkK65eM5R8EVJd0KkNbJq9SDQYfeA
5ebQcaE/UaHjVu+ujOIcetIlXVn+M/ZDmEFY4RqCzPl+KjYP5FTnAAtRVP+Lx2SPQrBMimcJfa8/
7coR58s8Ufv/GpH4KTCCQfPO2KhT/n55zMGMbr8S5a7YmWb6SQSqLD+cYAhztYtMnHGKRCPP96tx
uSAygpO4RZfkh3gwdfuEhZgGk+hxpyrdUNfFjPvkykjliMor4SlnmUqNtN4ovuDrTULLOqL5CY9P
s9L3PndkAyld/NkX+H59ARuOBeslhgnLoImn2T4tpN0l2gv6oQOYXV8N0n7GY/mtxvSNspyS4xLR
Km2JXJGB64QNgSMqvUHSVn5p97zNITI07atF/qODn4Kc6ViInBHYwKwkjiyeKTpNoOMRov7nNHm6
GEa7M1PqJwKNaKDwB8VGJpVJzJK2LNzFAUgeoUlG1vCF9rRxRq7x+XEHcUi0dzAEF52f1iJOxzaR
d5CzZTD9YZlU9RGu8Bxdzc6XuO/AOwzZrHmuZsQx7r9wnLZ/vwp4WHHKsBsVE3+DCeeRtqXYLDAI
hacmKT5dWqJC28qwibhsCQA9+5fihyxvNQSGCQbKlI8w6s/Z3CxvAPg2wciTpqpXLvfyxMWIdkhh
Ad+i5kqFQZTRZG6F+oYgNynrfcZ88PDre+rEw6J4/HDQukklk/Gi2Qn0gkGSX+VzWfCnxRIm82i6
BWRdNWLUavNQB+poFoAI0bwk9kvvGhi1gInNq1fWMn5O8EI6OHC+RRWa/rzyjuAQXto3YIE+e25w
p2ZhgQQaN9R6NZWWQx/f4J0sLMc6FxH6AL8cMpQzEZnbvfvwfGrGvcmwsD4+zqKaJGzYqGHD+b99
scFfUwBq3+cnqcKhI7TyjLSYKSwzbdDp0CwgOg7srPvBpCjTYkt3RUDA3upSVIdm+SK8aJMVEdtP
FhUjxiPGIXO5+T10zLi4F4/OQ0x6HPYpw7U6A6fJkxGwavF9jCTxg1isAW+nzPzSNuBRBdt8bCwc
8HkBArKwsFKYeMJFFQrjWjP+0j7Zonf7AEydvPD0CQkvfO6pUousMHk0lNli9Mle6XsQJk8v+JOO
vSf7tWmsg7oo/DL1X2yGdaQJLBDUSZ2kjLVd9EBpiD8ZdUIIZ5tQnPq2frBCWtgkg2YPKMOytGaC
4agGuaIfrF7R7/svKT9KG+ZzxmUBLoPkfAQbbkinC2ytJwKktBm5Ybi/GgBL+Y7U39TdIi1abgnQ
5gJEfP/P71RHh7TFNoNpGNAsvhNQJwcF+3A7AbW2qWz2mlfC6vU6LXVAtNflE3HEwnFnDPHh8KPH
zZeg0vlJc5Lu8hQcfJI0KCV4wFy/ZeOvfs+zu8ZcYweJLWZ9wKu91d/ROljkLexCegVSzRHLXonS
miRVmX/RW4QQDssxO23FrlP2hI3wv2VMWU/xrfCY6ZWq+JjWO8+GyGMz4ZFfySNYRYoweqQvOEYR
Z6bYuQYCkOCG9p+E8CjAOxGtlfYczJTITDJLFpfWvaUaTch5JhdpjEFl6wkKRhmri1rfPx8Z/x4U
SKDB8JRwH5k29mElj4tbjDq7D9ggi/o3R/TYJZSv2s/WSpkSuCNjGpTH1Okd2xo3OCqsmJBT3ppC
6u6Bi5tO+B2BPtUhTGWnXCj9OTntWEC8zVRraSisiQwvBoguAFKBiNGQItVO+IGt8aSKOIhmpsJ8
VMjeEaPmzJyMgHzB+bev5mdtVmZSRgEFxreQnpqH2+DqfvBeFQOsLxqgb+1Pu3CIwwvnsGo2LONd
Fp9SaJo/cB+AlMVKruskMxXVTKEzPG1GGyQ1bFHv7A2LzCtDv1SKNQYqivFlxFUSE49hPAUO4W7H
dD2eYrpK5I6Av6Ljo51IfZxIPBJ0Ytpe96LE4Bry67/DYemJsYBKOlksyYjVzQ6+8r7q+/e/HpGP
PkRBbQ9DLMix/TLs7XRLU2emSO/GxncDdaLfvvXlwBYDg/io24xrfQisyYnpryGZTNPK3bdiWjyS
mIIbcbHVbVKzfyFCfOYsxzkFzsesrglNzEgk5xGzV0rf7tagJeo6RDQrIQloStFbv2aCgByEmGiH
f3UB+m5cb9GBTtzaHtO7ZYgs4iySwFfuIMOS6F4hts4+zaZlwhSBQjhpwsSrDSH/eTixsVL49Wrg
dUBh1147ZACWwFLs7DCazpKrf0AVvCh/IJko62GG8gKOfdYDFCPmdF+D00JmhMX+n8rPYyc3LBlT
HHNJOxs0YlCNi6DsMOZ/6X+soMYFSm8tyUcn8Zj49UY8wF1pVbvg127WmWnS9luNxUtt8WdandPq
KdwrrdcUvZW12tM77iUJ7fKkx0XcDS5UG+glRb1RIhPuUEiZYEYekdipxWtKg92/Udh9RsE7QzKl
Jkil+FPyldVwWACr9b9mxBPddbQPeDM4eUbV52XQSH9rGbZJoVrzVN+01gVm2qA8m6xJfphbJx6r
zpXT+70NsdMPtmbp7ctpFymATPw58A+lfWJteKs1yUMMrmOf9HLFMDs3imqoX05HqEDPo6yIoDVM
iW1Fs1nvU9/eCK6qgR408qEg6vHsjdDCyzl6x1EzwXuboWbEwqUB14TiKD4zxC28eOveSAxPS52u
M+37xfV7n+jOoWEkWI20rUxYGljdfQr9qh3K7i66I/0u4rlLf+/D8AWjykuCqrpBAxD320cormlJ
QKjk6OiKj04Mcn3Khlg9OZAa/LMmZ/NVNWuMx00Ny3JqAy5+58ha3wDmKl5XkizIWgm5MqyeNnhc
1+oL8L8VI9wzzAntCaai1wX0HPws9jcHC22ixAkrCIHjKwRS32nPVpl3dAxZfvZpLgMD36EXRR/Q
QaJ7vNT8AwTIyxk/pI4+ZD5j5Tqo40fBEqaxRVtFCnvt8BE9e+WQuxcnpU8MwMItCkBUFCYyJXsR
lmB1eeowRQWCvoxrDjmHTyK8C/A7RIlnxaA8Z2UogrQa8nNOdhjbPhf2gfsONWb5Hzg0OXKVjTCC
wftNyQN1/Z4HhL1AuX4BXp89Y6d5mLYdcmjrqhKi3znqdT4DAtdWE1zDOgpLdy/cx0Lwz+sUayVH
Zj4r4jCVU8YTlLmGHbLTTpGn1xDDmqDLXtxJ3tp0q+mMBCROsmBmGciQRFbkmYGFNYLdNkUCaqRm
Q3n38bsIlQtiieQaO00Qlqsu7sbMTFKdGMChtwKMYvi97G3APb8nTLsvk97jRvJmKb2Zukb8moKP
8r34+WIIfOO+VAEkykhM19ZW+bEJJAHap8lp6SOXQAWdofRTRTrlDdls11jQxI3oqlWHFyYO61+q
NDoqHzxDwhs2+dPYLlv4woXCpEEw8v46Oep2TEkSw/HhGravh8f3iBbh85onDJRuJFOZfkLC3q5Q
PVSnDayB2Xdr+ocIk4d8VpWsNj5iVZe3KpxXMuEHcEF5MBi+k14YGRCrQiqj0/4hZq9EqcfVEZYp
odKAZMXkLwCYH5hR5VzleZ4VNMn/fb4cg7Kr+JuP/CYc4rC5piHaXF0+OTkh64sLWE4jH+imR9AU
tupJqhLnY25+/ghVvFOFaS9LmjIemognyYYKHvNCPxw7UwQnK3t30rpZe7LM9uqjJYAuVGMRqXuf
5+gb/32Azz0BNXLG9iKs/wVhgtdwK1xOV0IcJXxGSfrlJK2u+1AAsfNh1C7Ka/nNFOeCP0Fax6tg
u7co95sKYkOhDeTOXoWx0XaEHEBC6M5EaBI3eFliS4tHHicD1x54uRX8V7GMh4zuWuELH+JCRUFQ
NLh+5DYbR4t/YVQzLVEmhcd+5hH/gAF9wwR1dSLMnZ+bZmZQeLZ6Rokhx/2KyIUXBALEpwdPreIC
Q8nC9Om793bUA7Ty/Jp5AdUWioukxgJpRe2lK6Gx+ufF2zsaL7zKP6oKp5x0dm8Gz11sIWrZTSV/
j6+KMdfvrUKoaQ8huGnHpSxBVgroiZZVqkHWsJArZX9nQkWZtqA2FR/IT89LuKZQjA821Kab1P+m
i8cmlhWwqfeUq3aRgwdezJhThUf7yNudORvcsXCOCfwiWNEI2I17TKwBun9hQrefA7GqVo9LrqP4
U8CncbFrnK23gvDY5xnm5ILXAIURZOs0CF7RcWwazGNGkFzOPTiVl+eOaqr3gfeV8+iGq20vWeVW
fGwHc/72MNiXXA9ovS93IkNievfJ/ENfp7dEKlidbP99q/GzranR+iCCxhPeLjDONPUMwRUmep09
EqhSYGGidQEs3S9EXmTATMy482jUrU5gg2xRyOMRFR+clwMgsI3I4ex1jyRUFj6ro4T8I/i4rsPj
9sY7VU2G0XvqrBEjZKHa6TvzbqKyIJTAxtRb9JCgyoxZ9qGRoJW5KiZe4KEHsV1bmQ7gAMfBB+r4
APsPQCA54I+CUqQW0eUhC+M8ZMpuehmsrFrXQNR4ibpu2j3VjGvK6aR0hEETMvoKIJOaXv32TAx6
CXrxHe0XJ5NzJiAg9NrIRi+aEP3FR7jwU6aMMyS9IsvVGRrUY0Ka76YOXRprSNojGIENBMnnok0i
skTpl4sh0rE6kmWjpGOu5puyhjcN+KVdGAu8wahpbCaz7CJplC2TTNOXxWLr5IgZXqLJe4CvnyGe
OiAKcO95ZwBqzdbayRthco5tauXuqazHaD1Ok2UJ6+7bZ+6vHRaCQJRQmCJB0Ay3yR0DcQe3WpjD
BUXTg0sXLLz6VDDg1IunYAgcuze9RX797avw4suL8Q8nPB9d/wiRTUUztLuQE2iyoh+eqgri3i7o
I4DoZoL8mvORtDO6GLplJvW8+66oFtE+1rUWBjAqq6ObKLkL5Xs1Fpz53rwbvYRD+2gOtws+pnUc
ujXKfq3fIzXbdIinZ0IGvhAyqnVBji/ifMn7IMkjyx0oU2vvw97KXC9aGuuwyn05KfNP+1yFSi39
OzUwYbZj1y2w1gfZ36YTDSK2b6J+eopaFgm+HPh8Uuv+dlw8WXzRIzYOQ61RA6hRM1T3M4ln+bgc
3XVumLUqukG8J3bfvVgMtyrrU3GL2hhK7GOajm8+jv7aUCFmjmI7KP9KDJxUtZzjW7RyWqpCBnaS
hSGaIboReX4OlhBiS1WdfWHwLdWzPyqMO9IneTa6ZrhT04NzKuUMW3q6IBEONjoPdK7fJ/TtiuhX
YsL96XdiK8krU0u1dD/nh4oXn8yLGpigP3yrkFd3tA720WuH8HaDyCrcpmZvaFpYxsga2WFgF50L
ElAMvX808Mmo7ai2+fKpIlO/+wO/AZD0puh1jO/u0fmtmZerey97BVu37rLh0/uHhyZQRIIQh089
B/4uPb30tLmTY9OzQautjATuXHCvBjbyMybt6KIU1/oGxGP4V9O+4stkJ/wAp28yNt+qH6WEQJYR
uG7asIQE0Tw7pJWUpA62H/fRvhUD1mYSaXiuT/NXsYupV7UyvOwRXNHacV/ihrgvIb1yfT6dgm6f
E+Db+IZM251XddPWhk1Z41R0/OmOmIldk4aUvtc60gCRW0h1gT0J8/QpRPNihYcOyOfdDFhrvSLi
gbNN60CTZi1aIYJ7feTIJNN3f+kB0m/bc6W6Eo+9+wzeoyPfa1c3dvl0pFlFmfbLT3CSEOGwpsH7
wqVuOBRHc8fVeSje6s0juXEFRBDKK5uhwwIsnBoEzq0gakqUUQyciwAoP9IKkV2ou6zvbXqmA2Wq
qTZxR/7QgM4j9kyDsBPzFK7hlgD5UfjmmNS7F25ahO5LLqeBKMUlfEx1ea1qYurfrxeCeg1TEAO4
v72P7LV5ChSWHrWB56mkUxWBjlJ1bsRHF52zZJAq7tWRxio2Ef3WUxAF1vs5PBdGkhTX3zHWCokO
ebv2mRnNnfu4eZpjIDX6f2unHKkmERgSSOKFUKuZyzdduijts8x42czmqMeN4lFc9YK8SSZzZkzc
+dnurbcFjdxPh0zS3Rvig5UXg+jJZjuv9LMGniAgRzgRCplOgP9Yyqjla2jaNBZMMYRPPrQyMMVp
ESe2e76pO73KNVlAW2TkIYYqNeHFslTxuT8uLUO6ijSPwWt3JkBaOuzTDuR8K/gapEJ2Vuhcow/z
2F2hu8JDnoSvmVTw1zEAJ+b5NBgdJ+gFa3kG/XLdRpM1x4+UM4Vocfd7kv9m1xLc27Mum9p2s9H+
PAJMR8AiZwMKmDUoqxkJ7M1sl5xgRRGF0Gdwi/S5V1d/RJ7Tv0NJ3IwSrRjPmyMncZZ88zQukVp/
gWlvGvkzmtfSRaNmjnBkR1gQTxhZGniJeQgfHtBn6p/eLymdFf6tea3aaOhhQSt7/8/IoCXgcU5h
Wh8sLNOsDVbxCqTAt3yAG4+JdRQdcJuUmP8v8AREmMnlS+meGtm/q0P2JRSQSNZ9r54TqaSBCxPq
g5jeLN/7AZ9/lL+fSKFrnR4vLPRn4bs/PJvFCrG+eE6f6BH9n2KHq/ATIQhQOWkL4WRJQXqjTJrq
m3GKEdbYB7NkSW65rrTGsk+3e45ZIMGfuuWuogxYWt3Ggq4WDHd9NKTEgxQTz8TDDhl7qgebZNgM
Hifvsnu99kvunvLPxVAUidPWm8AvI1s063A+qQ7JCDT/rEJkAVKwWijWZ4LBKgsQtKduP50flsrx
rWO/N+VRtjL4xtadMlYejtuaoZgtT5V0e5QZWjmirsz1FOTyZ8XfBeOMoZqlGhspiuG8zx1mK0hD
zDDDFY/ejbwBQv/+ltBLdc6wRoMU6cSPdxcZmHQt/J3BC3WTc1oMVLZT6xkogmyhbmh/ocFmoik4
JYe4+YgV6197YQ+ri33/zbmCadacCJ6Kg1Gye4Alh7r3JON2GGDFkHKPi4SosPEyBsRYk25hA2Ds
cHH0rBY4qy05TihLi3jtsXZjZvsQSiCWEJ1oFUROahCNryHXoQQ+2cYYqei/6RM884MW23Ubp5qs
txMXpRaMM/3QmqffWoC9oBEajsY6S2b6pXtWEVcBj+Kz/0QZyYPPMynWaxEZLEqaa3orYw9BR5j1
lUYfv+LtSiYezqpYYgjTbWLn/OlS11nnYBFMZ3VIHppkPwQBoT/WEgsZfqy2aHgnazKQ5pnI/zXR
yz46dGInl+OZDRfx2oVoHg8uK4cKozxnk1jichLqY/gTot8/WGhkqylXJsHJUQkiMX7+MudGSkwa
yluT0ArAO4KlysGq6nTnODTGre+1lhzDju0GRdTujfLeSWRkVyVKj0aH0FDEALPxTFQM1/k25UzT
9rhxufIdr+gfm8558OWFPSu1Fkrxu71+Cjy8GT2FJNO4uXiinlXugCf67yeNpdaUw/HcB7VPxnYA
G+VIz483ReSGxHQW4nMwY96wfbS6Or1FqaydLjPgtzgDwsmelMGzsHgE2SYIiLLirtodCDPIxAEQ
cynICdpKjBNtNbnHF0beHwbiI0PCF1w4M8NSdRdKs0oPLjwcb/dFW8KSX9QdiLFwAYYAEtljm5CL
7ibfcJni92M0qPKv+kKpO4woh0HQSb/GPiSLeqe1p4TIi0JgfACPOCpNgot1hxTtDC0ukHGkdO1d
+wklb7LRalu/EHniooqMSt1iHspz2A33Q7rMWdqzGh0fbmovG6D+hvyxZaCzpCnR9Za2XCvtcVYU
i3DGED/LohDUFpPCSQzcKxRKLu3BrtvPIlTPMCb7mw4mp/yJr1hijJKqAMM1hK7N6JBnqDM14nVr
wcB5NP7m4rSWek2b7Mi64eoyTf32glkTn870impW3dDuAdIyai5Fn1tIXhnV9o+Orl+aau/VtHe2
7AnN+Zg0j7zgOarpgG/tnOB2gUSX5Vo+bMX0X8MuNJ57tB54aB9tzEjSwG4orJ52PTQFk8TudaL+
odBicgYQOUl6iqk+rcPxepUlhAor3YY7CaOObW4SaGI51998KTzcRdXl+HzJlbEUcmeNDqSfOL0r
gx9S8iv83PIvqz8BbgCapDSvXIdZyYX2QPk+t49i5xfCRZKCQ4Flop9lmU+RUtrGM4q/p1BynX6D
Z77nc4VOFNNyr3EZOsKDFn7b5vQKBL/o5g2q516KHHnz6k3fyTsr+WcaTz28u3ktixD04N7/KlKw
uwmP3sSC8gjpMhriscjOTyzQkY/JrmoXJcE6B4ZDTPuBm77aAfi1Sg2B/iXYuq33PaQP8bdgD8z0
LkUag82tXzybgWPWEB7hG7GTWxHZ+eDyzX0qLj2MUOxE31q7txZbQIsYSeZEi7QEfIr3ZLIwrcH5
DCynwJtmbQzrWqrdTkDvjxSDva9ZJd6B87J9q7puYLuAtjdxyQ9C5E9+Y5waDA4H0+avNre9hYjn
Q0NXnuvjbdAsB61hfkO0yc82WyTBMBcPN32Af/GdU4vo9/M9wtVs+/XqyzxbzDddnSEh1PTpAXNL
f0wSggZccdH3TMezXNW/JM3LYA5jfTeKfdbIM3Yirbz2AZnCSnaFEv8omAPIXS/vCLbIMVvhZ8JT
Fbvrj7hhW3bHiH2DMLrh1WjXYW1JgwugMxscYWj4FlhfIamow84RMkc7Te7U73Iw7xRQbT8QmbJK
3WAVEFglzmvWT8+XeSgDJMWJnEttoMTA+hg5osHEzmbVD+8DvJaujXUqkRCYWUa8yXxM4jSko24E
iv8yB1jx7CyZCWktOLKj3YiNASQQ0TrE8qLfUssFQSpWhy+YGGxb5bClJ6Bh7CJYgZgYtCTgrNQ4
j0l6hGZc5Y/TfJ9iKibgVKtHhF1aFqEREnk6/BsBODmtV2W76lvJlWBlPGjj/lkYiuQc7KTIVbDj
oc8FV3BMGlJSqFkTQ3FBVMPdgImYOBe2MsyyrgYOaMEO/yDVcNfim2kC+1jQzyNnvHF57pMlG7Tu
3R02WlemZ6zKyVtL/9CZJ0DhHyYsofgaQ7MUQJg52COEE8Q0XJbPM38WIqzrYK6DCrsdJOEw2KkU
rD2MD8MbKQ/i9frGznNMGEWVBHbaPdbNmh4WqmaMvySUbnbg9Ym3IKUc6zEXXP8Q9PMFe2aYhvYH
mH169eoHd9VrEa8J7prLKUcN5xtsU9h2Tn1nYluH/gsj6dGNjJQEE6CFN8qxEPLWFY4ea5AbyX6c
JlozqtGNxStFNp4yakIiC4cQUWd87DdJIL1cyMnRuiwAesu9DRvQA1BhPxVSGpn8W6loCB/y0/Pf
J6nCby4lz+np65ITKHC8CbHlhRRt5cPm0hC9O09nPRTky8z02+kVAX39VWU1cq/7jCqZVltXscXj
hXtyaF1PelrUUQyNq4+S82F+AKjK/2sd9AzunWWwbnyv8pqaZDuRz93bDQHN7y+tltLqErPon+jY
7+w3rApeJvecvKfNWqDYabbLdhOuEergweN/x5NvMgTuSr3xNWSFQIdV4AaMPsEhsrIw9x1Bl+ae
r7pgd3pldXnhcmIxuFGsXHdDG8c08sH/47Mm+SxpJfu1TwKEm1CvRDuD1h/sSuZ04hG5GMHuXn3h
fIqZzls+cMz/d6y2Y9VB+N07w6HSp/yRS8WrO+l+jm3FP7GTHmircc5qvip0UBq5MtdZsAhOrUoy
sLQ5+Vw3FBbT2WkeZLXCer/fPi6gz7Wz+bv5E8bnUPJYITTNMFbFwrntRvvWpAz6az2THYHzJFPy
wKkrGeCkPmgSzkN6ezM06OFFUDIg48G5STqPQMY8z8j4ZfY8+4AdGvZ5M0RlpoG+ngbbx0MI1z2z
7972WRQMMy5VneGcB9do0iG+wXO9HUI//dzwL84gYojyME9tf1gggDv+hdo0wSyYvG+wDv9gZMrG
UpuFZuNlIGGKwP6iuCeniNmXvscjOLMuBhDFv7Wz5yETaa28v+0DTlG5bHt377o7hLJZvuKEG//O
/vV2UaKaiW0C5LZuo+P8f4oKZit+jo0HglGTFqGQrBqS2Mw/zDS2+Fv9kARKWWaKL7LpVRV4IbDZ
AZIOCcYVZkjwDt4hE1EiJKS2EKyCrU1DnmcBtCjW6A0Vb89pAmCl712vS0is2jRTikv54KI5BRX2
ZGQVclO5YTPiev0mJdfa2BK0dI+p1wpWU1JzfTwTM7TAtt92LYrELZAiXEaPHkgYOlspZIHuvv29
2ddk7M4r74wTWeQ/6SWRpWafsoUlf+wXlgQWLy5UfUwQSVjf+ag5N92ypQ9zGd+ENmYyDFFgUL40
CQCY6LL6HQS/nQmgDSq4sqRerSPHjQIfnMGgYqAZXNTB8R8Wjf21Dp1V2z57hSdOim69fPClBAFI
htZV6vMiAxtEfNrWdOSM6+oLNpc8LO9a5UTirGn53Q7y+Ttr4542gAg+2y5ZwEfxJuNbZxiGk/XV
KbD3I7NwRRxvHaGQjfwdTYDqH0vgoKf7rGse3OBfQdEUNFaQwlSv4Sja/j6PhN5dvIfH9fhC6wgf
+rQQPR/1gEXLtcdA4j6IR4V6RbO0eWvwYn4BVB3eh9DvAdp2o58WaQKmLZ6F0W6NhADuAaIYa2ua
QJxJYednlPiaIxQ/+1XdehE/mc5uLRW9y6Zk0jWCuuf9hzxSqasYBSewZF6AoWxJ/Z5E+LazDPX0
4HXmZFXeKWlnE/0Ew6u3R3V6fALWq+fzHstlUpn82xy+Lm0DE4u9q2ZCTJ+om8sQ6cQK3NotyqKX
Cl2K2YleFEkVqVY+12W6UWTdgOOKWEa5BxWH57RnEqZ7/ZBEVXvBgmOZaUbFZpc5j5ijvrW+yTH1
MPaBH5vphYr6dx+Y+KJdLTcaJ2tReCr29CTEzNW3WrnB8J6REjcMmqGr7J7NjzRhwLkrStfnL0dL
Bhwf+znanmI6Qc1/PQX0oNwTPaTNfaWVMGGuVtLpEsZoN+YNX/hQgo+lAWRd0y6fmrYdtQTX5UTt
izqRwvDDOWj+fPjsclY+yact2YeDPS81S3pBMnBmoiJV+Do57/VOmUQl3JB252OqIFQd2CHUGkqx
6Jc0y+NtjddkCS0SKBMLcm8dY3ti4/YJo55JNnc+b9sc1UA/4GIywmdjp1etTtTGFXSM6V3m47cl
YKCl3qrA4f8sIED5+WCYR+tPX5ERwjjhrYYS1xRWPk/OgkfIE9MTVkOCLhm0rS95OwOqVf7oGl7M
kgKrxS3ZvePeqU7d9Fk+6vuYvoqfz1uQL540XykDovMaHKLJJeRqI1s9RWpjMqxyi3gaQGi7yD1A
9JFZBbYP3cVgwWrVkjUdcrsLcssVgIPIcI+3AJqbQF1kfdVXg14Q1VysWifMaeAP/EyQpkLryBjL
Vm06jqJRf9Yl9RfkWqbLpIRrAJLvVajjf5kwHLaL/KszwZot3fR1CvmkLmE9et0R2Qc1PzZz7cL3
93tvFek3y8qaOt3YOHraqCikQURgqeGuced40oxO00CF6XRooSlY898KAE66aCUb0m++HHyUeFPH
iGb5xn4tnbhN3q3lbq91JgVeBC1Zt5vVasK2UHqu4Nv06HWiauSbmRmUezJ5b3d6yKfqcasZBHvn
rGRUaVp5zavjjNWBFsaVcsHeLzWbanf4kqyjf2hLQD2rcN+eoZwoB2Q6pM41Kw3jslz13DyxFLA5
msJVycEs5SBt+odfmmYBFwBXhZRbfX95Oy4wpZ74VZT2YgRIgWTGLQy7ArQ05rR+/3sUQQF77Ovm
Bl+/0EGISvNLYU0GwsU4h+1T/A8ZTZFeHdhGfy61vh6jSpNVZFa3MTmx0tTN07NTCs18m/gBpFTH
l0wrjE8EoSV8o60VAbf4tWd1SijuZrqBek4t/6U+1rhg5YilFF5l2YK2whAfBm+42hA+829X3Ual
1I3jU+HWErZMUQTFj6PZc84xhtW2MMRsbKTBYozffweW4J6heEJ0oEh5n3FgyvvliKet7IUO/z0y
nmmb6A2VsYR2/VGlDpj3bTVilZDXjlsro4I6hfn+PDjQ4mmyXmF4jN1+6TuTZ+76O87EOx7Ccibe
u1bAtVx4SwM4d7YpzR20Pf1WaAteciW1SievE/Vl6gMPMSbibK1rWVbXMDtlZFf1HWo1keid3iO7
4jjDs9KReBBOZFjmzOQUTqUo3ElOT85Nm5PGgDromljp2V6vNber1vUWJo263K9lxOW4F4QckL9J
h0Mc5tUe1iOM8Ge2pPA4MZH7GFBL/CpLpjP9k5z5+1Nq8DLJzEOIK0Z2iH8bsXcIGWUrDscqHZ0h
m1p6UrRHNQRinM0xHKL5sS8mlVmsvE8rHTfFXgs4xZGp6e2PxnbkzBskQiiv5GW2UacoFGZFM9W0
vPladf2eZ3KfKUj/dPs/0ncCbAtfDGOgyRkc4McCAZDBbfDsGP3FZ/SRcQvx1VYs8mc+V5lZsDnl
WbMt0/49xYn4PGPLzBRs62OYwEpzkvof5XGDcULQWOnyFC9cpezsheTPWZnD7Qt0fCtKcmvQ5VcX
lWzJlcNlT2FPgowffGfKQGSUjdrK90JfQA2APskI9p1DbbfmJcMEza+SZTDx0+Aph1JObVvtLipT
YmPGOsbQmeTKbS9yq1Zp+acK7ucFivQI9agjm038bOZFmvtnMYHKOQW87ZkeCoiOi2YfaMZVNTIf
GSrLjfedgBVI0XdBbYW7qSuCfs8NNIQ3CF/+6s5qrS23H8FInCUV8XWrn59NJWYizq8cqpP7GM4o
IXlGqMqvCQ2s8pLDww7c26ZZaDJNGjTujiQaqGNuZmT2e7ZRHZSX8GaRWe5XN8+V+qhpj6EnbR6B
T0J4s1FrgJw+NSuQTBUg7VJGhTCT/MV0wQL74ZAJwqyZam8Pcg/TgPoLWwqWBJT0fC6jAffqmlCQ
J2JmBUvDeaPRoypf5rsW3iXAZJj6u/E1fFWvCk4uyIIw1h5eAHFZYPuEEU8PxrZwnTayr7DwM8r+
CIvlwnBjtUfU5CPRxJPap3HB+JS1KxyxxElCH28AmUmdEFw54OwZZ7bGpe9YBnW2zBqPpRN5wF66
ucUCncGFBK+feIwdXnJ7FqloXwiknslXhgd88P7kkiWzjdyTUrGtyWsyhDLRNRepoY7uR6abTmwv
YDPWn8zppMGdO/UhiTkcQsUe7UZ7YKT6VeRg9R9QbiA5e8hfB+a/e05/o3zsImW7Riwxo28R+qbP
JKccSVLkKwPserFXNha3aWqv6ozdK7ScfRsBenLdCb+XRzVWYyirSaup5Po9ck9YcDFMAjVzatjj
Z/OWuvGn03R6nruA3tyyk6h3JDR5zb9sqMA574xmE38FqMAmKnnU7Y4VSZhXu69upjnFKrWsYTUE
7PMxVp3URrr5O+s1aMfa5wCPQrjRbcmS5u8nWUM3LX1GAm7m4AUbSZ/d9EG9nSYnuaNdbzkD2CW6
YB26+RPBgYU+G2odeOsk5fjHgpnS1CvF/Pa1Jy2q972ZZrWuDQcCfKqWvimdAZYIsrL5DwHVpl1R
yUgYH/T8EtS1h1oso2Dy/eU5/pbjW2baIZtK1TG8FLd4+p0wbGbhmM13xw9lcyfyj+PcZXsyxcSn
CQLntLxD3te+nhGYmDFG+ANtAkaB08Q2THqyPg7qlXMUOxkMPn9aP2ooSksKse37yyi9yRTl/3G0
1wYa3bBS/UThs776gjVsYFsZSvPOppLVXS7+okUIhUjdrvB7rS88iKPx8cFzklpJZD3e8bbjB/NV
O/eInPNPXcnRMuVHoUdNm8gDugdkpitEGr5Dn1csSnnfDpfAyH2lSfbkC1vDQ4pSct6hmyjSq0JS
rknWqEU3TgGBZoq22D5kcM92IuOt12xgiMBzeD+jOE9rBjMGovVdzGadMdiyPZQZZZk4SO3ONabF
KQ9xHqo4FOLpyRpFOatG8fMUTLwoi5GF5hyrIW/4GyD07W/ReZkzC/i54B3gALjSUZo2mxxtzcfr
AoQ7nRiqwZ5DEOrqPDd2eLYqTQ/iy7pkugDWj0QBmy25AbH5xMDicQaCjMOJgs+dJSpNpCk1k6eV
+3wjQ77hwdoRh1c3HHxF+qPhBHlTGnVNBgHoLsn0afx3kBwNS+ac30h0VVqHxJupUDibjDrqnR2v
JpAbiJ7rMihuEpQMBTSuIv7Fv+a/6XUPbAMcoB79Aey52TarsFNel8i8+ED4Neute9wDQP+2BA/6
5VqBuPiZkLWp8vZ2kaOfckWN5SZneQOzob1Av5eip7PhPuOc5+Mi/w1xHV1T3JCsMXXZkmYyV6wf
DJxkpz7RxtNbUMkmMWqRbdCOaG7mMV5j/RXM279mFyGwd1ZSoGn1c6YLIY4DCH/QlbxFQTeshcyt
OwqZwh/J7eUmFbUKbOENW2TxdW5Yfyb46IoZ8fe+pDSak+0attlNjspfb30III62FekLZg81b0BI
ja5VuEt8P30K+gvHhZp2GlJZaV9GZWzhRQnE9sIZRmP5Z+yaTZVF5WKbsLwsBmMeEKOLSOO356u8
40eX7ZGENNJSeCmOcW/kqDn+ULAcL6KUzZyxq4KLbZnGqLeqaQUcSre4BWvnOiT0ECCmA+CHQwGE
MLu/ZnDZHOnPuFS/DcLoazwt/yyqMu6Sb8xTmSzN90SvgPJkU1ZJlFv1tS01TYIp0j4+vH8PIPqv
1Uk7tPKWB9/EDAS1GQ+IAoCq7EOHJEy94PKMCxVjX8WtSVWjJDyvgotZ97f5HglyGNrXhZj5vNsi
UpWrBpl6HPfn0ZEJ6vUi756MHwdX2qFW4p/XwzL/byIHhb7hD3K9N6jchOq6dTfGJCRLJ6a16cis
pjpDYd90SnVmk3oqQNbi1cv7GZDRvKsxs1LS+yhjHtDOMNMxpPaPNFwZev/HJNhas7CHxoLJn484
BLc3w2NK5ii/hfAJH9xIj1+RyBfEy/dUVoC7sX+nAno3OO0VhwgIy3S8YSoAzxT/rUcHxOScZtkG
pIARmR50Q4+isk+9KUFszfmJFoDGibMzqkf0oZUmMzFkIhEfbKWi3rrPNywPXqNr4eKNH/O5mvrQ
RpnExcuAulq9t57KRCWHYvpwoiRsZxI+yoShIML7EkZu2qQbIsTEyXWV/n6+1z4UPY3nGMgka+9P
N+kUTJhTR9cvsczsuRcKN9cT32+GOhJPkrhonJUW3eU7fH/ZW0u5r4HGPOorU8DQfDw7iYwXuRpd
7usJ2fY32n4zhtPcGS6Si9IWa1vYiL4gN0oS2bFtvkyUqaUInU87LJAMIUXrsThKa1otultcZ5eu
U000G4tpPhmlgWC8g72dPTGmGUSsiT14LhemEa6jv8tzhuFtoOFqmjboMPMIMYW+EWJxtieHeIpe
UFAdepm9PUc1U/y8vQi5RFIP3VDctEY5G5UDWnOtzvmyvGrCygako6Yp1t8vEzIdEeR8GyQyQsD+
vcRMj3ATSxc9OQSOlodCKXM0sDQ/tqmyeMSxjtDPEBlpL9i6+9idC11TFs6g4dDR536z4knbFXi4
URnqaOSOP5Gmjx2h9lhvSYTvFqHA++7sqSOJsILMNyNqpidj4F6YJhwsjngdG7BZxOxcDtQk1SbS
PJWouUdak+hDUYNQucCAkOhRKErEHmEjrtgXKeBXMZCq+T9D+NEfHKtddOY3FEkXaCmG5gXQ8t8l
GPlWiZDvqspGGnSZlQ3RDKjsj/Av7/g/jvquDo/A6LV3HWYpQRdcjnHCSH/fhkB640NhEApGCguS
XW80otLLvJtE0IAdChCp8XiFKzMDrEBfGtb0Z9ajJEs1aLXTtlok9Cf94RNUPQfqGWlkkExcsmgw
WTKN2g9DFilznB/g21sutQaTb3Go5UulANnX1Bd3Cd2tWBMIvrmlRvPXxy932c0vzZnJ0CBbqUIq
yYpGktaobdv8vfkS7KBAelbfGM3jIPfIfY6nzxioEHkJm5IcqHNlGuCKfCeO6JbmyPJsMEcra6Wi
nhpOHlr5mB3/fcli0UKT1q0ExGbbo6Ud9X5FsCrVEkkvYtid2LmGv6+w2CKCsWiYEzXk2w2drlcw
05l9l121fdW2nhuZpCsL8b0OyGAAMxXrc3Kkmq7RHixJ6lc9iecCJvvzIFbvSTiV7oZgDIwm8YwJ
QAat0rP1vGb8vU/Zy3xGpGyszk8NOb+7cfAv7G1iyxUvYvjObfxPvYAStPRcBukPMEgJzh9QvVda
kmtS1D8NJlZdhvPK7Mc/IZWbUpvmQpHeJclF+F5tGPGPTawGD8RQmTTu71PJyn1pRBb+IaRlwhLu
5AftEEg8LlDHAklca6+Zu7o88wmOkaNIMqA0y8sc3zXcQSBqkrN0KgazXKny2fQDFLhOkXAlEufk
pcnoHK7di5/N7yyH2B1RosCW/aqOfwUVQxIcydAY2563YQqFXZhCzDQK+FSjKtN+HUEuUdP8IjCj
r8HRSyLb86zJMGlTdFHwhsB8p5vSuEtTa4qS2da+4NhomTWAQ15A608sEJ3QkzTDmYFf5yo7vZ6e
q4VGupX/qtoBeaVghAsCMXP5mFn029P1CvVaAoV2T/bYocck+Ra0oeY8R+Vd9WOZtREZ0AmtwiAM
uPyM13IgxdEAUwzl/LftOj8An7yF0QhmsHB8vtmSTu4J2SlHw/+fwIOdi20FJkgjAcFj20tdFqX/
IuYVDnU8hK1OuLqBQSIwvWd8jjsnOk/SydiVZ+kUfY5W+9hKHpMIy7feTM3kHZRIlzeKWI/suaEy
S++KJ+62thrXQvVZGo1LOLudeFjT6uiwdRPJZT5K9p/zBSIv8W4nURuOn+oo2hXWeA6pUM4tLlhj
Dp2v6VHbCN7WUjrvjp3+XbIhhxxvSWrj3D+f/4nrgLJrOZWAWhP6S3mvjRnJ8a6DC0SyWOsMvBGY
bbS382UH4H2BEvAi9WBDRDPrWXtJx4bDyqMBF3gv8ziZZD9hSsuHGGkppWpCoLqp/WFaH6U00Bd+
E00KQqhK0qShvr1zYJa3Sz7djBnqiNX92qN1uDo+GdoGXxfFbXBlF5qtBv2uZ24KAeBRsdLgFqzC
enOtdNW6ypfMXk0gR+gmWIYZR0rbRA8ib8rd5ZeT0QqvifHmLGS9jXhsqXXk9SFAIPVgh0EAfRs5
BQ9t/BJRxyQrzhFEh5r4p23vaZ7uD1UqLOzaAJEF6NK99a4VRg8w8dS8W/TPbhTVdT6o+N+uNGOV
GfnKqDnqKffPfqMqQL/U5euIpjnTDUi70EqMJCrm6M33W4MBXV+2Mtsc5py8wTszEzorgJnKyUhb
NAuhVvNKx2+WBqWHAGgURySsfRCe1W51HMo5HPyeNc/FrvpKTq97GBNbLIzN8dTx4b9fRq+VxPhl
UeyBytLdAYNeKiOrCsFG5NyphB/ugQ/Ky+hScNCZ9tki5zFXipC/YDIjVLWLigRs/fb4R2zxH+d0
1Vwv9QEN8/jnHPNGEejVKmDrezPbRhc0X+x2dV2FjXWzVagL+7IV1pAGNFa4w6Q/Trfwh0HbD/xR
kxwITzAKUuYwTdmyreLnk7mz7EckAXHwIv8C8hEnUmIremy9rGyiDjh9+s/gqOiJi72ztnVZiXCk
DAHGHVNcfT3JKbtiAsEwU2WZ9AGoICg/bXLTt58aec5hDk8QVhM+FqZcdngb7TEN5DN4eiEmnWHd
TW7boylGByO8kQVVnb1+HGGcqMQ3+15DXNvkL1P2FPG9ncMcfUEDb4IX1/9KfIwborE3/RKbpKfQ
1+wVpV8fVBnkhNYx1Yc4+NpwMnbpHufjwkOi3fBR7qeahhpl3OOFZLVtgri1hW6c+Zk/pL6Lu4DV
2AT/4e1mkvuYaJGigm17mJqZhT7kGNtdyhBsiUY7T6sTad4n7VPdS6OVZU4UAspiL3oIVGstDDJR
hmUgQFj1PqsvoEzE5vPY50j5TVDUuFyNbKMJN/pIsZHz3tTrcN/VU8p/Ei9yA96WmL+haXPMsrFS
6FtGnVjqS+WroY8/7ylGR2XdqL4ajkUFiUd9KjFCUG4ibIky9OGwc3mpx4BmF8gUw8dIy+3a+Su/
Lu7XLU45jqr872SNLRwG9lVk+fqGZGW5TykBBFrGf1AvvOoQPnnaDNoMjEZ+D3oQEEOiW0Egv5mu
iYWYl6XtCwzLFZpJowhvuPKPFeGYPlVuUXksZ4mYs4dq0N4ED6hngxxpI+knW9EyF49LOPRmbq5M
jGrVD3U/i0KJWUl8ek27C+5Nwv+HDE1iHv/YouAIKHi/ohL8YKxqdhANTYQuydvxG7Lgxu1yLMt2
iGTgqiftm2Q80cbGUbukPflkf2Gxmgxb9ji6O5cbnhKOqWJ0LLBR3F+Espy1s/Umou8UiZF4wQ2g
XGHVZ/8mAHRPmIeYQkj8m/c76YhO+6spjcswFsvV7FggCVM8GW25QoqyoeAaRRpyXFv35qQIyZf9
0Hpx1uAqZLEEehhNGtdjmOQ3jjdvK0AX6onqK3XTLKYxxNse1kmC6KTxT9JxON2KFdGjcE15J8Nh
uqXLwxktJttfcKthY0rqp08Ey9VxTlqi+zwyCFDPZR+MDHak1kUXmtEqFkN86lQh/kzWlVIYNkCv
krVf42InM+KkA9oGlUBe+ImWM30NPrbrJu73xK48a+e8oIMD9vghD5Yi5YOTiB42ePiEd0O9A7Hl
ioYzr4nGXVzX+3ubG+EBC5GkUv+/hq7o3akbkbZJe7Vpw58we40D58hZYqlw2H+4ehMkpcuQmT82
n5M3pRrrSmW8Cj7UoSJhSUFqI55IBcRmRcwJFORVPacD+rn8dZuBU3SLjTnMog8BMEVMrb0UCWDi
nKK4xYQxi+8w8IzrbjFSCF/JaWn0HIvxZLlKB8lRliwkwiey64GuSX9fHIL4hHtJlWjq6rphXb9G
VI5B1zH0S/YxBIL6VIyAf2Kdwr9Q2CUGyRSkI/F6/77bBUSn+NnZVDVQrvaP5WC50PisAGN2r/q7
0UmCrkYe3Jorgj7+WNrzXDQihL15XZAi2A/afcnGRcw9tcguQ9x/cpAcUPHfVLyXgct/VDLIDVKc
vc6dFCIQmkH5kQ6BGVcy59m52sU5SeOGVHnC/Tb9iICLbyQ0NEscEyS1nFDjOPHp4g3aBlYliSML
H9i8OtoEGcpE3FqZiVuocUr2PMgo2+Bzd+h/2dFpsc6IUDKFdDIgp4nGrFkZHnNwo6KUt8XIZpQq
gpjRAi8uP745LMs+pF6gjgo4Wz52pO99B0RA/uilI7Vfw17G5wyFkHstY+yEOTyijjhWRUqqv9qP
xkAjjihbHF9nj+PXm+W5WJIxj9VVf/0l6ZlsEBoXZp/HKzy4Ny87RKYEfEAIJFYv85xcRXGWvoIk
VQ5bkMZgN5Ji5nCC1DGgXWH8IlBTphdy/11G1JEW04ufJqq/n0Hs5TQYEXZoFrTVb9OPy4d+fNjj
iB/Fh0c4/O4sqxJCFjRP+hmJibXpNJ2/Pib0+S/JSQb3NZHHXTaCzDRK/eR7P7iz0n8cCXj2WeHl
EDj/rQTMguTpHpelvOr8h1/psybmqY4KVQVOXHDjBiiyrw7ijIo/PN+R5DwpDlxBdb/ewS+1caPq
kX1PCr2bdZGebSTwDPaAFLRqgZFcstIuAp42yY2x/49O7uAG2l67YehTTB1qPoKyaj7dAj8Nd817
r1piuUZUSbVLdPxgcI80aXsbYmkW5hAbMWBatAMV0lEmxk5gBAbH/zpF7kPZYlrLXqt0zfZUaVvk
0TSm28NZeAlxrFmmb+QHEC/YNS/hi75ttI6jVZW+Uw3tkPI0SrSLy4x6KjKXtk7DrXa/oyfPG2n1
vdUqjhbxqVFl3Sbcxk56uIGNpA1JPzpegL6iPCix5y9AfYMarFTWEQ8WWKwkUAondDTbI0A56OMs
5zTch8lr7ZrOwdYQ9BItM4ZRJ7hPj/jI+pJGiyby9nqmh27weyndv9w7zOODLegt2g3GUL+ChvCt
Ufh2aq/ieRREwbvkOhEXLZ2UsbIeoYIc8aoPK3L+yCuaTPyGTmD+1D2hh7l78tfBL0ZHQzAwIlKf
inE6NV+YUO3AS8nVtHsZuWYZhqHJa+gM0pz3vhrz3PztlwZSwm5XKFWemKc6PWdybXs55tzwM/Ap
wug4zxPxU5hsBzQn+OpeSgFUHIx8JbVSEuVWoCTuwWJx3Ji0ULTl2KzLK+3YnQcX09pnSWFzt43x
fClk7ueXI3PhoEsFmCY+5CUG6UnjmkOuWl5CEuflzsv34eDmBPhu5w1v9LssAXuvninCzLWIdOaB
R9IMcYhTv7fY41sEgwqHrzzKF98txng9e2GO7DHO3RkrLFUd3/cvGGNa6Eohk+3/dAz9zM1OPcEE
OolHOv0uwvkoTxYzs1UlPPQNNImhiTGTk9Gnjs5a1W6r6uLkbLMmE7x7ebHb3xzlzp4S2k8rBNzx
vXhUwnvrO9JTIlYwPQyrskBPTMKby1KK6u1WGFv1IzW555OdC9rdIcRoFYWn9TDOPY1HfY1nzZar
6VsB0xcHpi9hOmL+5jaAm7L9ZmQ2uzZeN32BNqyCqSdPHGWJ8CupWTFjd0uFsnZn88Ksgcj3HjfY
jIMDgTkAre+EzPBFmvEzPbHaXYpU2h33ntcTfdEihVS5ZFd37t8EtAesPCcPbcP2fatv5jrc2SF1
Cq472RJHWj9VpgOL7hSLQtXcBar+q9MZJbmX+SOAojw/PitKNim6JFF5rFkaIHajA0Xm9UfNwbGj
bfU0NawWHSePfP9LbyrrrAPZNCp7P5mHH7FN596hU+bFF9LFzvmIB/IjEP+otgVQGHRJ5axx5EMt
tMyKY7VilkKW+5gW904XuI2VaC1UqQRpN5alPOvkqOSyjEpravdiWfY6XrIt8q3WtPAthg2tqdGt
OM6QsnB4ogfOEiZLLfw4aXaGRGqOhwqaktI434yNmyk66RZq2sDRCHwbPAYJ3CV6OozmgYtoUaMl
gxPPakOK1tfHakmZvxHq5DnfttO/kUw2P3QARcq40LcWPdt9vzkZ3FHa7RrIxJiMi1nRdN3WfHcw
kpf0IhxDSrGeiRnA5kpDdbkOBYOfIcEqYYrx/ZMj4bmq0QSAbEh8OA4voSKukwQqGF5DLiW/fj08
Ybdelw4zNJoNHUHFLRMjltn+avLyMnidDStP2sr/+uFim1T4j0shq+XzwoPaSWRhLdyw5LaRsSPG
ZvRUAc99SXoZC8LFzEV6tkkmNTQTw8hN3DHTUw+a1HaZAAqFT+6juYzfCdyFF3dLfwvhCA7AyaJo
OJkjyQ+tCVksNKOLd1ZmhuThd3AxkafcwB2EE/vdLFbj1+HwvNC+D4S46nGGzJixhr5U2AuGxmeK
ZMq4bIP+6IQPbguVWeKOYsiqjvahJHDo0z01R0XutN1mxV3uIOljBY0kD/t+BJE0BQEVeQ+CNJrA
cU04Pl+zCvKRNa4vGdrjlOF59+zg3euj3955KWZwvixrmsMRXnnZ9GiU1xsscmAo9ap+tBdWNqyG
th3qYbd5U1eRjn+xqueIMtSx3TipCZx2KSmwUjLKKfvIJnUNC6aICwC558OdCXx9XBhvaYDB0bMX
KJWPyE0KAXlEzlCTtlntp+vY283j1dFkJZ6uFlmOQzmGQzsonzrGdNXAUP72a/Mdds84HXuiA0do
uIU1mjyCvd55CjlGW7wmBoqG/RdsayrlZCWw1g8R3YlIo26aN7GbaGNUM8ipEEBI9zh5W2qRepZW
GYf0eZ8trXSTofKeAQ4ECtZq6/WvKESW0GUJkB8K1G2tPz6PlKeRg1l2HrX4d9pXDTG1dPlfU2iP
foAUKw1soDOdlPIgYxyBM2wY0M+uogp07zqLFccx+HccoVvowKXpS5wfb5IGFTjf9yq8tMw/1iAe
DPCVrEp0rBhdDDrmygziaOKUBl62nLB/XcuuR4ucdw+UsUUviHMzgiDoSNryGZlg7529loIjL3Jp
w/SbD7+e1EFWqj76fQ+5yPWGgYvUPB1gt4EMBd+tIcycNuClQutd+OEEbHIF/lvoNjBpkq7AJC33
uBCvkoARlSTrst/MD8U2/3gcNdv6zbXZcjbSo6SuM3mo9aPxd2hk2z9C/cgyOC4UhE52zTz/denG
V7QSeNcuhHtRnaHEZ8vEmbRtgLu/ECsKYd0b3c36FZYY1nGi96JXDqqe8p+xkl4z8ISi49GLNK9I
jbz2b+WDNv0iI0LKG2mdzoWwZve3HdnXg2BZG8WGiO0tWwsOrPgvcYMCEj+F+259Ju/dSwBGhwLR
fGELcTVx3LqpE0pMH6SnCqde5zQ2hfSSO3TUzndhmwpR/5nCyDR4B41e0skadhga5bfQckGzVWAl
MYHKruZ2U8x11dVbgfLb/AztbN+ojJV3lA8IYf7QqqRc2l9SA4D4eW/LiW0DVbDRuAx14Jnkq/f2
HSHEF9c63+G1tG+45owL68gnjNv8qlBEe2v6toJ1P/790P8FTd3yB87ALJTbDlzDAUT0GXGmScce
h2P/slBCZQjNrSLekUo86FhwLuSsHX3WgxVrpVwCB+vPFWJ8oknwmHrx3Uq6Pwke0nJdz31GP1h7
mw48gZePc5zPoBem6GktqsHhUxq57mTcOhkZHHfo64IMoaEaupRez3/RF1ymwqnpbcNVJj9eneov
SaVQyU7SWlkKu+en47UVIgG1Y08TWqNu7ckJ9ccU3aXJi/P/0xv4asiHokHha/P/8pyNjq6RqzH2
gxnJg/jGDzcCo2qCpC3r30m0acQQL/xpLl6PQf405SbJg/J//+73+K+COHquyY5z7iB324tLeFKP
jDBsFo8HP/QxNfaqK2Rd+r7tHa+FL6VLCFK7zsGzEeGOXMRWm3/OAp98npuZlRizEpH205h7ZkbQ
61RMuhRQJOjAPneuxVyvAtabFG6ypI20OyDZ7C4Ivljbd77f5WPGOfWQVytsUrJf12EcLziY3kg2
rUjIrN3Lpc9c2QA/snUilIx4H9505wxmYiyTYU/TNN+xjThzBeIhJXI0DQbcP9sWi1SvRJtWbvxH
hm1bd8huRrIOYllAXwVlTEfYR9DVySp+aqkwRRYHFMywG0c6titcpaeeYeLVkmhFjzYvKS/XDBOz
vbPviTQtV4lT2J617aDauZ1GkcsN320vkdCeyPnySyfupL3Zm0lYmqKnA7adYEX/mQz5VtuV0Ryh
hJDsKJHWqst3lvz5QQrogxyL29Iy7p8y4HRRwpqokifEUxrjeIC/xpJE5DqqOxRodXBgllxts1wL
qU2qzB6Q//n7BxGCzKSjYiqTUkwybFe5eMzlIxX7ECMBFyd9fIR6f03f+X7QxLKv+Cf8DDq0ng45
VpazCKncxieJ37Bxrh7inJFm4CSQtG7Yta/L/Yai/rLo34b8scyDKEaahAHbm/kagmkWy2S8JFMd
n3U0PfIT5t2UzOW5hPN6bXG7ZWtWGhug50F7pR+DmenADrVldHeDi8+YcYSCq2ixSMzcm9ICg0kS
zvqipQL5HgIA4TqXdyjUo+fCh1S5sKnL0X/4fv+KVjK342J79Lc9QTFV0BhTKB7x4aoivmHSHg7J
GtNjRx5ORGL/5VYjoIkgeErRn5fGD0ydC47/mvgL1zeu9WH86raM0DkTiGloEythYySL0YuDgRQ8
/dqxJWZWPe822BtZh4ynDGE+0gNso6xRyqMJZSZmSF40yfORdl6uEt76sIgrSAREU1/ku1OZw6TH
G9MvJ/hfvf6Hfrxrjho8bJh6bdbCPHnMhv6sSumnsYY1JboqWX/N6PjE0vYbWXMdjWKVlt1qk6iE
doqYLTnMR9FTch68qLcoTq1cYXUcJ82hEwkZP0T5BuColIgi9bmvdRjiiKDkywxIBXBLS5wMJlxI
5GmK+7LozyBulfiwkitDd8ke/tQP7FNgWq40bTsoUca8bFuuMhdPmWTacgxlih2c0GqxD5/zFS6u
Qf3Utik2m7QaRR/U7gU0BWMcXcQJuEvkOraii4KfJLWWrOJ+Vi6jpkAgaFp/Avwmjn8Db6ycjGBO
ywDi2X3WgOWDtH2CnE85SScgYwXdhYgtbFFoZEh8OeE5sX/ne5n2BJoyNp/Bqge+KUJcsxAbnhPE
FNoqq4kXFs+OsgH3lP8Ut9Hvu/K1ltgtgdNxTeh7F8QR0jHG2UanVSMbebDHGFrEtLWpePPL5UWT
zv5ck5bZCHYev0V0E7HMrY7TSqH/Rmt67qq0e7E42Kl9uLDF4hH9tWBIleUAlVmzfGI5g+hY5T1f
BmdeJAm8TQQLVsV/FxXyUcHcs3oAly4P2fcvfREqAJSZDTEjl1hS3wjUDUWmB8JCqFESqww3haa3
yqmKU0tO4FqFKOlAVUi3dVXn7DKpq/p6LE6KNJlUy+SF8FEbyjZs47N1zylJmOIbOAYD6wxK1tzU
LoLA2fpFsz6kmuQyWulPSMGa03WO0pAHzBVN9eFHBNBYJUgrLvPep+M/hqMbEJ75HO3AkNgbyJLh
n9u9cr4NHPfjy/csR3EmI1fm4/0ziXFUeZKVgsbPTk1PgJNiL4QUVb/nFUQZEXI6EPq6jCa1u7R7
C6Sydli+PDd4mjXmBLryDXQHYYEwLDMKXGAP5qMFKGKrh10JBRouztrDdBMFtn5O+TlH48kWcqk+
hx/jocpy3LEMPkMyI2iFQMvsBAkl5sju8kaoOHh4H00qyOSY+8uuIlqWBCLwrSgwVaRZH/4hG56o
CA6bpi9aCRucNqdBPgBCYwxJXm+/ctT3g/Lc1Vj4+cXlEk/RAogFDRllPyan+cPLRIKGKdGf641Z
U6JfaCM+p1Iyd0QdpwfZpcdZqBwkFilk3RPqlVN+/SpWkHQmUGS8RLdBQhlFTZ6ODfpWUGcWfvHk
qJ6FkMJMkhCvWSslN4B1Zdc0kEBxqjqwM65GmEAjCuhGBsJk1sDfXLA78nyfBvA+Yx5xiL7/+sTA
OD72J8h+GTZzwCfbDwT58/5b9fzWSNvY6ouIrn9RkemohkAFm2Pjltaky8kBc0qhXaVsGYxtfXoJ
LUIhIa4ozz5c03YoUH/bNgiDcqO0Ztj3t6zSLz9L8RQlPKcUL11+gTYqqU/R6v/IySNSEZjK23Oy
mfbwBwXGKZ+wheAPwCg3r9gzM7HltwnoiJaNwMG7Zcy2NXhsbNxosVsLmIBvz2JJXAnULr9H0n3x
jIR4EWrpsGG2S8ljwpew+L881KDqKHpO4MSyzrmN8/0npcGsBaNjFtDTOsj8NmtpEReFOiYFSXWj
W2OeS3cQO/aYor7wxyQ0grBbV+hyIGRG/vT1KlgEQMBtWz0diPWdBhZ7P0IOfA8o3N6lQ+w0ob+c
OCXShaXwoiM7v3OPo+m7HCQn3voEWff/lDfG6kHH02C7FrD3Gqq2GDO6TXSzI3AwG99YuixCGFDu
okY8y1uZblk04GaDTTOScWKJuEw9Iuln/OE2leTJ1iuDeS2pvQe7MtJK3JRmkADHeONbgxVNXgwz
tmVU2a6wEd1OzkZ8M/nHTLolgiAzMVPdQxBU0nBAuLCXPkBbhWz1WBDH0OCc7lTjV4ZRmgCF5CVS
2s7/Zjg9dJu6WxAAJzsogU6xnmzUPtt6uOXBxp6wmC/vmS/88sAqZ+8uofYSWp8Lw5aMS4JlPkCy
Jfn6T7rTAXmAunylwfzoC8UnAprcLwtXbhH4F2QCfZI0ENGDsZXeXJkSFUEnXzVPfFEnClrI7pZH
BrA18+wPHbx4mB6Ss1yXIn5EBFv6H+dSQ0iqwW1BLu2Qa7FbUwp79EOOOT2oP4Jq7T7TsEFYhPFB
xbAzTgOIrt3+XWvBa4VKoGjynQAmfcKdpi7WtIFDNflDXotYJnXSlSSpUyjipF8svl+7PpJycJSo
CpO2tqCTeD0QLn1PLYFIljjdSR3SkPEpdvVSqUVqBTPx57hRzCJUuYptEW/+S8His2FNZyo/MTEu
eJO6evFrRyQ13anJEAhhgCIcNxiVUBJXem3qZMyKP000dZx1qE98rWyzUrJyPOpoVzK0uHTLNEKZ
4mrMuntb6bjqdNY8pRAudZEcP7dAUUWFMM7R8lsg+Ie6Q+EBJiFwBmXRbJso2wmsqj67MVriPHRf
oj3rD8FY6eOPrbHym+XjM0magxWmFT6t2nQ30/Vngpp9PuhpKjJvjU03XdkNUA51Frjd6DPXKo6B
qKs/nEgqeQ/mfVEd0S1f87GHv9kLv9/IH3DmKNFuL1aTzz+MyRobEq1VOSYHEVbN/OClwrBCIs5O
FlJ2mT2NexhRYc/0oVyyBboXy2/eZSEOfL+Yk1lB5tpK4JZHasE1VxSUY89Li2jjseY9UMY5GLiU
SMEjSY3KT+oio4Nvw+gr5ZOLY8FJ1gKfqkr+shosBoojIIpFcynD2Xey6gA1Azs2U1NS8JPEzmdr
Jg88BVxm0ioXrjHWdFYYKb/dCnQ664PejeDynBglQQbF1TmtCIYw4CxFysfoQNlo8afE2953XNXK
inIVCgSTtML0ugPabCEZAta+xCDaRDbycS2jrNVRqgL7T1j07T11zBHkDRE6aWhCNjujo8jPhmvJ
TWU0HDOUQc/AN69P3veOdbC7SsWXM/BOShhiXYACohVKWdz0iUWLXoynCZ9E9tssicpZBYCX5Xdn
QvT2o7stl4sKwxWQahhYODhiUF2y7qfr9qz+BDsmrWeGGkTvlNfcDfzcRS8OkvMsXAz/k8dOxPYR
KToaJBTW0Q+LZYgtlDC8IfSZVCwxzX3uat68kSFjeDDvVxMwafqTrtyIimezLLU4P8Q2u6DS7WBD
3DnTlH2YKD3nUfRiN4o/Mg8e009nbDy1x0cBQ9MycdFaTlU5QJINGXSOHyUIKZ+nl353Pogd2Ugx
c73ZjUkh1G3nH9HXKuX3GR2NcrlfQNj/OUGv62+F8k/ku5XEN8H3OoHYRiO4i1gMTASweP2vQ1fu
tSS3JDO5fHgM6uz80bh52xqZmdArruS0ZsNzzL8aUehYb1RCTjKv+vI5Us27WRRLV2C5v0eU6Rj+
n3j2o4tY/SE04H8AEk5ARbohPIYCpw+uMQSG1z487CDrGmJDOr4RnEFNhObRt5E7kNa2TF1vKqyB
KzJd3cYy2yqxdX3tpj95BVhgO/Vrro6+DC0DveOiFuBGMgrefeHNdNh/TtIeOgZyJAuW6QzECjbl
whulJs/RZHtA1lfs9gbG/tgwAkzYPKFBHVMYhBJfAAM6VPf/krwoynZmdFOcc69+lNLl54dZJGC9
U0J+BSajHb8W3vxXhZ4aeUEn1fGppqvDMUKlpL1+kF7y8sYsMFHeSWhOQzjNZbgtNEr0hgfF2D0P
ePnfQcI1ATyt3qbduJURn7V3Q6SwKpOdsOzwsZLm9w9Tx0Bph93EFSUeQ2Z3DVCSD3v8Qbs5cdFL
MzNQkJr5wX5Rmx38K2oUsf5tz49iCC76noSbgEeZgy+6Od6+f06pUS2d92W2obqndMlG98EA6X79
FqazXgETqWtTY+8TlwX0CJDe9NqCqryoTbmjJaB+C9mBrXiaHIwlhhnAL9ryAZucT0B4vxI1eKLZ
NPPSQGW2Wy3KruWIPDGBkEjA60HN67K9MDvi7crQnCIXadj+FXmbo+jxCTNGJlrtMv3dVLd3H6s2
7w9OnXHZK9mfoNZCrRpCAY4Emwbg63dzBXqq2auSQbboXdXpbvhH/dOHNWhMhFLdzJBgHeIqYxZp
jTcmBU93d5g80pThWcBEHeWs8jrThIuD3vQ0QRoRjsIK+EmpKAIwwm+HqrHDt/fr8R+7+HzjS7ts
fB4l/o5bgMU4hqvZ5XJXCvP6Fyi3ps5gLlE9t+RUYc4GOjukc0L1Qm9VD8od22b27lqKvjs2AA9k
ruMqkEE+px9HZAn5oi9FWJfJ/UdURVKc7Q1z1pSDKbd0qOd9xEtCUvXfFtUpCrJbYin4Uaml6xXJ
HjVbV95LfXsRDDbo4Xum9OiMzSuw3ozTqzNoyQsPvv08W/xNAFSJGDLTonF3x1LvbsBKGiMyTcwT
hOkE5BNzDyDppqqzcbFPqBauTXM2/FHYiYrMVMmHD5Jkhhtxg7y042fXYTVzxUBJOkolSX3VtX4d
uzVMSvx5zF0+3nwRrJb4fZ4DwdqvYIoi9NdWoBwON09qq7T1uZIpeXDRnuqVpYAceez5Ohaxe+o/
SRH43PgHWC5igKQ283z9/oN4ScRO4Vhioxuhaa0w+pQQdILE/p9dKLMXvCNbmj6QFlvU7WJZGVs1
Zhm62jA1j5dT+D+oMoiroTEptU62L0akE5lSCPj/vKy3MbURwb4mJV2JHbwP2x1T64CxFZhSBVlh
woiCc5Pl3LVYwKVgLTZXjYaP6jK9bExZT0Yemj2qK1sQybA+P3T+6QcQNq4l7qjBOaWF7hap2WJ4
BQnQ2oHBu0g5dmaAg02iSJ6+80c0h3lxHdgMZ0zJHRtLvMe8tXiO96t6mfo3SJrNKgQTSxxxzaFm
QYMoCRoZMHD/tqe2Cs+qlRH8bRJEwa4sBFdVNoCndU1t3CEdsSUP+5/ZX7VqfO50XraCwSQ2nrq4
v3ijLO7cT4FgYtt8bbro0hzhcXPHArHoWLFPQEqRzbbMioMA4a6c5VTwevt1/RusE1Td6V7be3DL
LU00Ha60zsHtPedzipdqmNPvXirgmeOqTze9HzHMpWslV1xLlwmymM/pvmA12IrjXSB1VYtUBJyF
3f4qpZlFRYT6K04fFasOsmVIIR7eGLIfAxVapdEMDV7m5e6WrOeYQaYER6wVLphnmfrTEOnk6P/9
WCZKvW9dvFW7boh70ZsD8YzuWtwkxfEiy9clwd4xMxQqGrU8go7Tx+KdgIcaxxe97Wb1Q1WWwHfq
JpDIiNajn7ddZ2uO+qQxzpO4iAHIYO614w32XrDapgkatvldjdLEJ7I67TGd+AB1FDaW2ykwxJOo
K9stqnruVzOsvmY/taf0ZUJq+wRzkzKQPuL4nmuFFZX9hAkEfDz2YtlxYkUJFS8jd1KD9456sl+H
/QqMYNTvADbPxVXwZ+NWxjAgi3HI5jhUeEv6RDOEN2kPianpw5Qs5yzRFTHeGy2fvhCj5MD31KFT
q1Q8a/C35Jeo9UCNstO/vLOzmM0RbGQC3+wUOdzb1fHWsbN2nMLBlHMyuZ5PIShLF73HFRbCGDN/
A2zegZOlTw1KKivxMds9rfvdgyxnOKLWkwjdKi67rExPNpeq2WS4UFaAUUqIn2CgQ0lju2JFjWLK
UIM0mhe8tq25149aHN8ZIDb0bG4GTiKN1Ztu7fRspaMO+mcAfdq2UwJChFIJmsNsxPFVpVClnjQc
tfGdnJmvVUM4p2uEyDK8LXFV4I5L6vdLAOxvVdliUb1DzJHOZD1TQsc1nebTQlz29DmL+Jb93uYx
7iOsHmdNmDRm4jtt9V0t3Ro/6XODVNiHhX/UzVP0WNoS0bV5TvFKaPAyQXm2NUfQSa7dZm8si9go
iNvNvFtfVmdVO8xBxt9/hw/vb6OoVRchofe19B2vB49cWjMvHeJTRCppEXOaPt/xky7mUY+fbxNu
L1o6f2okF7PEwZgeogBNCbA28rYEem3/rwrSWxcxDo/xFq31XFqw4794J58MUO6PON0thzqE5k1R
bj4fQuvcqlnVm0PQ/Yv5MqJm+wLQuKQIHL6rI+h8VmgQyrNkZqGDF7vUIO1PS4Xx0nl0i4yjxsQ5
w+dEVusl7gtpURntXNZnAyTrgIIEPaviq8wkb06LvoRF4S73WQrXb1vU93tPNTAbgaB8jKV2JgMs
04d2IXdCkeqNGtrWQq7gqdUGJ1vIbQyasxjJiAYqcnU4rpdWA12dnfOcVtnZhgCW+Yxnh+ktKynJ
9ghnCEjCdSk+sVTCbM3aN16IqxK3t9JDawVm37cN079F7lIyfmjOlC2GJVzl45AGFf23ohlKgWzL
mZEVNyNiSVoKmsMXLjpACsY/wdYKyWci9QorkQZ7Z2iTm8zjbsC5VDqAbdIXhqHQrGbA75mp3NCq
2lAgzVdFlJwV3O5uAUV9R8S+Ns5vuRIad7jjBkCngzuqRp4TEawJGIUlMNSyqV4IlJM7OemZCdiq
77OgjnYYOnPHd80YsPuSpiyogRoAtNkNe9RcPPBpC/3kYb9KUlSH8rz4vbp3dDp2DC5s8RFg4zgx
0jcxsfMgLG4/XlDiLXj99/wQMLntDG8pvsjwNm/5UgrWLEBxnoYCOZXjGgThOyYsBvcT5ynJZ6/W
KiyqCjp8Y6PRnT8ECFzQzxv1oSV2V/JLv+gIZiZFHQa0oXDGdDOrnvHE2DimJ2EWel5+X7Z3zBFF
D240KAXvgFO0g9Kv+qrW8nbB1Nrh0XJZw2euU4fNDLAyOybsw2adTGzChsp7sxhcq/7aEU7lrIAj
7EpSVL/i5OlDuAedQnbscNZGLdknfYT33YZ3Zp4KoHETtqn+vyVchDxL4tMwtVLiV7mJ6TISjk/E
oRjNEqFS/K3pe2KocNzn9eJ04kSyzWRGGCWpYqmKf2WPEhQRTiAY6ts8g1Wuqu3Bfo8lGFyCnx/l
Gqi9YnLpIOqajpIYx64VQAGCu0rq/Ax6XpG4S5wONKoWdSr1e6RiDCodgBNXcnOzpOzDyHJ0dvog
LowxlBuxWq46S6mnrD9YKKfj/2Bc3NdWEtWeQvUNQC/xJ7W40+PIOyIugzycoL7tk9hk91u6FToJ
3fHQLwpTSzoROcch5SDf7fNUldAcrjbnV3PIh3Z8bWFKcwFkVXAFiPkEIi9G6QxYEBR+HkU2ZVZg
JSzS3CjF2ty2BIPCa9ejXIN+HBOrolYMjJjCbR3T6mbrR0+i/4bPUA3X/1HAlpcf36KuPJL9Zv5V
UEH9P6u7NC+LRfBt0CxqfZc+dqP+S8t5oOqVmQtH5fBS4B0KsOGQ41pUxS1fpwZSwU4uNzfra3rq
tJ0/cbZFAymScVhmMryEhtMyZC1QzXhdRDjQFTN2rrs3/t7b76bRYI2ghhfnIM2PUWVEowu9lI75
Ms5823tKfRLYfdh+2gfyt2ZqR7mg6C6mmR1qIZ77erxSSvpdPP3v1sZaStz1CANKEoBVzD+2c8X9
2jjqk2wb9ZX9BM9zFnWMHeT5GsYfzalpFTcekl48XJG/IrUmQeqwRvJRLouNt9LgPUnqg+DT8Nlh
TRFCxg5H+p0f2O82jwS9tAc+f7/O72fOHbs+8qrA+vprsZw8Z5vr1GZHLGYAar9IaDCdIoR7nzao
YyP/TCzlA4GAxO5ccK8gPldfmzQZF3QGyf3A40l/wr1l4qmAOL1x4OBWvnA2UeQwxrKR5CNgbpW8
4MfafvplYNJ2Is/DBNN2V3tTiXd8g1TeTk7gIBDUrGqXpr+jowPuRvoZvvbzLAxbGjj4tIwYqLJg
6O8ptu6j6Ite0wprn4R6WlSRP7fGjA7vM/V5YSQGRw3RMOsUMXsBHIyysj8AXFDacOjk1q6UW7ST
4qWZr7On/7fkanpFdE+a7/jwetgpMKngWMupfqKROlb247Qlw3jxu0/b0Rm7f3P7lQusvaguobp2
XObGjlXygXGIMKtlZqkXlenSnxQn5VNFf/6cLvfwYnFTKUNWHtJrC9HXPMNiG6TLh8jSsW7m1fXX
qJjQJ3hZkethhmmpU1NoXf7d1z7hB8QNaeQt/X5t9hMinuX6FiggEOLpF8Dlw6j8QjSWcXZ6+h/m
L53Nu9azNhMBErBJR3EbIRIz5ZkUgmSpRR7y1GFDIeSDR2DDv5QUAGi/Mdy9qpZ4lnqNZBJLEYqh
nG096QF7Cx8C2YpW6UqesqXOL+E13WAyBDfbJxwYv2FlQXT+l2dyoovBBUwTLo/bi7RImlnI/1NT
A4sNP1wy1I+hRKpqkTMLiagkTtzhvx5Rv8+J4TM7rCNjSV7B4qzFO1xyiKTUniuKMsbghVmax+E5
iIa7JG6nt37LQ43xWuusfUOwB6tP+gtZZ0U3C+IhQFqdpxxwnfTbIhcFeEJNTRZladoyzn7JzwSn
HxWWEhhklbypAgoXZQc0cmZfvod+Vr1KjMLvgpGijxam8oz3c/gPyz9oe0a5+Ae4q0EJuQJxSQ5R
yrh8ZmnIPvhtPll9Hg+7NHPWxv9p4XLGKN9vZbd3uijPTgqX4hPMnX3dcLs60smIK/+mpTqE3k5J
Muh/toEIX/CBMfkOoft4mSwLUkZVKsokP0EbVYYS37Kc77K2qW2Li6K7P1p91TzYj51hYcF8XTPQ
903nLZGa9kVqIi3UnvZlmb4oyDQUQXRPAEA+W4xwsWy+aE1DJTKylWBkCuRAnZ2noy/AFiuiH+ws
YkLluyjHc32oevn7Jng7uREkrSpy+1W0kr3aI9PSlhNyEf/vAGo7fq5X39QK6AM3JhSx05OZqgTh
mdhghO9oO4Iqilm3ABAYCy03i9aPOvjMf/3vm60CNK+K+03q9SJF3XWIatwCWSXV5cMe0TQwLPms
BH2avbmb2CUet83hnA6Stmzd0z6owoIyNi7AGXHOSiA2DAWlrimMb2K6rkCK5kNOwqhWZ+nkqHXK
o0PrTBUE3Qc/vFI0n2NB34mTzfXjPba1104skC1lpkF6Orq7gF7S4dw+dbLIndiR9DhjW0mS1L1E
CkRjY3WFXHmlDi+5C6xHiVUwwmgrKHhbSYtRY9TnN4oDdLOR0pDxVyJC0ZCHi3j/D0VbMF8HSRjo
NTWe3I8vcQ8ZoPNWIe5/ZNycWw0qZayTK/7tbXtiypdsYW1hPbdyE0L1CuB1ux1vjnEFbhS/geaQ
uSU48iDYvRPk2VoC7J33ps231PZGd3KG8oG8Rhla4/0eVnuiBHouSDGpzdz8vgJXshTUzhQiXjls
egh4tL4mR86ew5cPIaYYtRDi9qyvjUZdleQ36C5IpYRMnZinEpJL3499H+d13au3XHxZZNBPwRth
ygiVS7IFpa19oJs+xneo8Q+B1WhedInQ5qyIHRQsdJUqlKfAbjxe+zQ+OWBSRTU44cU0LIHlOasY
26KOEEHhjm+NDhsGeUV4p/Wk7L8ksBZGdLpZlG7ChdcbkQxAdzE8kNHpzMAO1hBy3tL1BFqQaNba
WW0JubuddyzQjdknWcESm5EMvzOAfzZtjC97Zy98TQAmhgMyT40vdWrioL//KUvqD342mz0CYzE2
7L/qYGkSBEzD9op0K/Fd/01/T2FLMa4K21y7FMXWT1uidW8aBQVkzl7b+MCVa4wA93TB1cL0rIuO
X4qwvhokZz+YqnuegWb+v0fWvnKLtMl8mH3nQVSQhWdlTQXENN+TYeVBsJuZ+cnknFNWZ95yL+KQ
1BXwmd2RHys/qwrTSHPLvTKP9fYPrYS+4qrXNtTDOiRHilkBONCQzGMs5z8WGKZbatvIZrEZ0FLy
oWg8ukuJ33dCRb/Xfp/SQy93hn0aG7E4Q3kg93VBjpCvBOqjnbMcuquwnampgk/UV5yqncrq4drV
lKlGs4VBBKs7hZbkXRg7lxvi9eS672JvI+eycSd2FNUEBccSt/zCdwzlbkK+bVGAr8KJURHwxCGP
yunP6NoN0ZL5/kNgzGevKYhcqd/RjPWIcAzMf2DDGgvRofqS9FmZOv/LZmFljxo4HJoqHhTh2aPO
pLw/s0TZ/NIVXqoAtyrRtIcgs4Sg7OnQ+FxVB91Gj60QVt6686cD7973uEVSbWSdvKykC/gcx/5C
5bamptsSvt/PclWcHvtyIgGtIy4LPeRo1JviscPlRXAyCaWctTOSKNXi+xjY/SXImjudJ3iGkzHM
V/D+ufN5DxnP8c68Ygz4YAaltuH+OUPLCq3UtGYpVdXLsx+VTLfU2WkUTkcN3InYMmJU/ABB1POI
ybmpfopyvCjZLdTfKPEcuek4Lz398AQytJuAF516JbxNk7k7mgYG6hMzkARRR26iegjzjNCGQzwp
zKjko0Sy+njLLmv5VUspKsReBw9zKx3EwHZIJBfykziZ+feWXL6SDY0YztBponklaQriQoWmdih7
RaC4Fn5+1yGW2mc+7QhT4B9+ewdiaSkG9On4gvCOvMEPUPAE8RUQnNnTCdYM+HLVhN5Mz55uIsPH
JVuu0+ZSmCsSyd9mwz/pqSlUYbEk5QTUZLLl1zdYpbODGg8KsXrquoAR42iQRQd9JQ1x8uY071/Q
bLXJ8cPToUzIEafQNFXpsP2tpj8v3guGqtvWsjcG2XUWEMGVKhb1YdTl0uLygp21BEoaAHWa48FT
XsZHwzsXua7RZxzn0Mxce/yH5kpeujBiDtdTOjtgxxgTLsGVWsQSRRdDxH8uAJ8kwLDO8kb/iLsr
Wwg3HWgmWwgKY+opnL2/W9Nptk690E2x4ij5wnqqE4xXvVN6ic0HWMKMcn9+YyhG8P97C8zvqXz3
mR8zZDVX48vMzrStWnmd0iBNwD08H4gFZWWtsHZGZfNlj1WLUCCvgNYrTT70zNPlyzdsJ6BBeZbg
iUXQRg1w8ZWMawWxAoTrw8Ic4QPu16X+xM24CIoAj3UWTrx1Xmjt3tHr93zkf8H7MpC8+bLKhjrU
GMvTJX8EqY5FecI407U9R6SrFbzn8SxJgaTuLwp0Myg/lUBjPxETswyvF9W9dN6ODw52aNUzYvfc
MhSRc8tZmoYzBNVgprYhhjbQZNXigArvcG3Og5e5XGWWUSRNUI11sb15+RdlTuPKOWCiPvRhW5e6
BFTner0uVr81zxuNqTOI0lRod612FgCWlV5/AzW2KUjsBsBe0SDGrwNf6CzL3GUsfucBR1yysmp0
sKwZ2F/xgei3LvbVHV8mIqud3sGBsfhBGc30SCjOLCaAD4rsrMMzwEcI0KxoJ4O7PrfRvv52qa5Z
zSkfaphDN3Uds/JTddczC7m1R/iNwhmC5r4OZYqXcDissRIgeWjm5JVoXGH61uCi74RZ16mxG73J
qBKbHRME0h/yFSQiv9MuYfq5mQRJ4wbu8n9rF6WuIlTu4jvOS+tOuTe4SKO5v5drugoQ31QiS4bB
dtHGhkgvvg7N2qxB4Xu61NyAqT9fV9Fs+yHyk076JztBAoavhKvDEYX5eM6SQqVwJguEI2PqsE6x
Qf/VVjfSp00x74pvLBdhIC1xcsVMShKpfeS1g8zQkUSZVd+IBY3K7eYIe71BCFx7YlXcGzuCjHUp
cOxFbdzueuL5pZAxmguTJGiAiDfTFCG3fBZNv8wbjbh945y4wItI/L3TRdbVCG5cY2bSbbXpUDqD
V9JEj2dnuIGTSge9sDmTM3TX2Mv4Gvh6QFe/uhnc9vtf3CsPbqUZpwSMVL3XyI6watHqY6KbhWZM
SN5XBlLQjj6dH8pqw61EM4gCQg2vRaLyEPg2XAm41GMQEFwKCTsiYPHpTWWFCNVwN1TiwtBLS24c
w08mYO5VeO6uANsYxtbUZjmYiYRsC0aHuZqozF0MtocA9acGO+UmhZuerd00GviMB3w1BEifXL0h
Vy5Y0v++yFbD+oYWAKDvi969IReIoZk3tEmMpUwC/3cJoPfmqDnb0ujdTfGoP6R78p8EkVt+/aeg
6HUvybjwyeUjgLE19W9bjX/kPklXec34gSzqWaqhHS/e84IHOPpjQmRiqsj/d0WrzqqNtLuAuFam
ZKA9nVyN2Bf2Ahk7Ym7AsUSlLzGwjePKxCdUwlWqzkbZuA9qS8urQ4fhq74tbHee2WULA20aOOIy
cou1nFnaTiDnmXxljeTu09DMv+ha4+3xW6xD1GgN0h5/fW2KdamTwp9otEXBE9bI3uYtmwn0q0Bi
R9vcWSs81frPDaR2tMv62GoARLLy3htZ4vAqvqgS+RxhmPOt62fFWk/GvM1tEHgVlM5qQ7rUF36p
8YiE+9+5PPSPRkhL01iygNUSh2JFq6RhZGILn2o9OPiiOexxjlb5v/OPc3Dykap9aBjUAsxP/1Dy
6sBnnGxIAHzVYsVZf37a+qvFh4IcIh6jrqKjw6Z3sGqZN3jaMe2mdW9FJMyJaGgOuW2xgvKvFUY9
9Kc5wDiiMMqYsH+CEgfsNsH1WXGn53YY65Hzm19wueWHRlTd/S/gV7S2yY4uvFhOKitcxpxL/UPO
Az+pdMTu6YVYbpjElb4IosZUuC9mOKvVEwF9yFJuBSalUBV8BtXyf1+YeDL2Twx90lU0WYnytiQY
jF/vSftLiJ9dRvMtm7mVfcEukcSHMXJUqkoIy2TztV5SO3lGrmQ6+ApWbTSkPYI/hXyZHV7bnbTA
mhgfnBNCwWLTtCM3KFrMAYwjRrQ+eUHrS6Sy8XT9vuNZQWhQZ8Aq3UP+JPBf0r13hSqN4czJ8lSd
LEqqmbHyKGRFvdJNQDaZPLRpuKrDlU6HIq0rE9qBmnBu4i6Oo/IdB8G2nDuwrX8J3U6nkYbe6POL
MLnHClWga1fVIivQ3IwyygBX2ghqgWKwgdbRAgg4Zng+kacEirAfnA8v6Hsf2aStHkEYqRL4r+eq
hzkTg7OtlSmbnfTDxIlHqiE7zurWqPTdAkcg/whCr9TK9DtCgEhQ89Hcq3ESSY3TfT/0EMNOvJDm
51U9NW+R30T1U+cGXnH+VfIcrovYkNrcEIYjvxRQEJVMfvmwTmOAUiUrwq1+z85amn44JzpAfW4e
/GjLE9blqvwTAr2Z0AVguSIzRkd5tql0nSADpHtSYyj4Te7KdchfOz39l/qktcQHx4SCeGwNOCDE
TjqwrJ0a4cAU1EvdCZaRxjuZUHdCZ9Sm8bFGcGvJ2+4U0XDsHy3uSqcAOIGRdQce0hnweKf3/j1S
h4h62zavkXtOKL83fUobjN3H3lH/6+tjNnxdpOQm8oPAuSHMU5VUor/F5yGjuMF5tEm08C+w/tQE
84olUqSdgD/PPqtlkq828UIypZdwIeRekGCojWeik1Gvi9a2v9poSmLWG0v1+KfV0Tine2KzNyFo
30TYsE0WNpcTjFhpcG2qZKJE2q4JJUwuA+upcfXqEfIVYZROYtVsZHgq+9Zjd90VjMCkqeHbq5Ze
DzDaZ2dHHPE5fKesxTOdSmEWumZY7uoZi1gq5LuVx8NjKUF6AHJr9OoSaA8Z5y0Zz7KLh/gzQnTP
dd+6R0UnfxYR1t6rrR1zfsjFrO4nJxdxVIk2+F+Rw/TEsJ2CgBsK+THolwS0PKMXFYT5PfV9mnY2
yBqP+Jds2vC72ikdpYJsPuTYaEZEmMD7T80dqktchi5JuHcO3Sx5TFhy4zLdpZZoNPFm6YqI5acS
McuI1rlfGlBh8RZKcGnbhNP7ii5EvtBjBCcBvN6uQ9fqMbuYGUPFqsOKtH+jOU550zEfGzWXXL87
uCHEL1Ii3lVjhEOe+ZS4FoFwTX2DDZz4WbXcuLKmGQEE53efxu8/5BWYDYYi/95CGvqIqohFAaet
u1u+2jXdRoBhtVgn/Bs2HsZDmeuyU5DXQm5bGxvTkpa3ZaegWJn7wkV54UBQiqGSW+K0xTTlOru/
qcSwTxWRqjUFepl8mgaDdf0KlrW8sKiSDcdXKu/DTpAJKC6X/MfH2w/KNqMrPIEhyA2Okeww2ef4
warOKcGjNZFJSfyuEtQEf3LlDZIT8UnFmLB6NdGxoO0fQwNL4JIubqW9PXXkxhaWCZ/ZSNVbTAyq
XibKdHt+XF1h4s8+sK7Obb4U0Tl/NwCdBDnZGqF83XMob0IzXsC3i//V7Ujb3auaZjh8QrfwuQbH
IU1LfyjzXT6Og4j7gYZGpz9j2VzYxt0czvw4Caj+ZYjA7nWnKvCtqrEJ6MxQmRXfW3GkPO3LX9I/
fzOhGU0RJp2iE83cZq7yK2EuRSlsTmNWQKOLob01I5uzTD+7rie/0IdFjxHeGQbDlqSOu+NNa8YF
mWDbkDTR9+iZE8EzmTr/UQTh5940oLWUeDHoYh8lRNuyNSroK3RD2jYQ9nOJqDRfYT24+iDtf9GM
LzSQZ9s6aK+YoxqPIZytf5TyO3mYQoOfBVLVF8SO7/VajAAI7tswiCkYlCmiBctjW9J87LIGGdbq
SWQg2lYlcZIK+bzXbJdv+SdfAJZcELGicuV4Rx8QObx2bo0Em6CUrqhm62QpSBINgJUAYyWoIRI7
Ahj7ZZky7UIwZ8uFbMnutcKw6mMOfxx348OK6qYFn9ldVi7+hilRqDUXKRgl0Z3TRkm3Jz/JDIvg
kE/tpQHWUjmcbhU6Nefy2vgavmmupYa/O5eH99RXGPXjmAY4UzWgFd26ZFR7HaDlZPYjC1qKPdcO
glSUOwMdolL1Akg90Kz2Bc0/s5MNjOX7AMjRERFY/d8gNNdsaweIZyxT9dC0CHJ9ssY0Pj+hxHMw
S2vpiEgMfU8/fFJHttaaL0cHN1V0BmmotQj2TEUc79r6HsOdx0K9ypRfKLtSrX46bB8LtQDsfW5s
3S+fh4daEcqCWbLy6b0enDr9EZz+hYWXygh729ZC4zAhjvGZGJVEll0PMw9NDEy+7KMaxmxlqKYc
5FLic2McM60W+p71txxwRndQ01EJQ8mWO/tSLTnLZL7hj4S4gvwPpZXe0Sy1TE4D/1jmLGPJLqLI
SQd9t3mgWS5dRBZ2xq+RaL+By3iaBvlG1+bcMejkE7r82sA3nSqMMKVcvmihPzMPB0SGUU/JnYWM
1Lu74TT4dlHpJOMSAcN0OF4v9CcdT6gFf1l9C0iA5NgTxQLYILWuRySdHNkpSoYbHt8UbVw9ZvsW
nZFUX3oDBYblkbIXV8qOoQMkgkTassWlLPU72Jwwx1ziu26DTYoreK5cCtD35HEiSGzy/Y6sE/JL
1ZItmLjTt6jFle3kW2n6RV9KE7Emx3zWdkDUpY8q2lvKo2YUD7B4Ln48SmtfHv3AxEer+Y2OBJqk
36P0xsEOJgzbbd0KPyEtIqN+iw93bzpbqcW7kysoU/XWclVG0ETwj5Xc7xNZGETZVIRfQzrWdhBq
Z5mpMOPSzvz77WmeZvvUTqT2nHWQsq9yBiAAd8w6oQ8XQ1MIag2TFpWMygMeaQYvu3ssefLTaeNe
PSUtEV1Wlt3/JyYENX9DMtbYkc/OZbRm2ItpluYJPyxrXlc83P99xV76iN2iRjV+ECV7+A19Yu79
IFE8FIOHKzeOobn00+Y0Ig/ZAIr7o6OHsE+WhYLGWY70WjGxIv+yiej0Wc8IJxjVp+BfVmRtNtJX
mkELS7S4tjKZ1JlxzoI3hSiZpvYK/txRomHW5dXVE6IQHy9kY+GeoTeDPhlMkGqdHVEHoRKHNzgX
KeehAbgvR1cbJEUMrgfQEYY4d3/xRq3AZw3ZPtw2BwbyBWmB/VM9fA3VsmPiVojUXJTHJABZCcIi
ySazvz1aH2Qa3C1AC1nOXVD3ZrbLrddyb8zmPKOqfY3FqOy0lO6pDM3S+zY+JhtEwBa5bWvGxTS7
4h8h4cWaQ5M7Mu5L6TNDv/BoSE0isn9GqijhhivehydYsfFCyVXRVY5XxgoZ3XU6uZWtM6NmC1v6
OULo7dTWMLABqQ2EHlulEcrjdUIyHKlPIX4QnRS+HzpXy7DmTBfOZrJwDHphCtx2/2z6NvtvHP8K
4/ZT57ylOZREC45SWPjrNo60GjRXuHKkFbLpY1sF3rqvvw7U16GyIALIXFB5410ducYBdwy8XyjF
UOYBepSKZnK1YUnr19Kj3VtUKLQHSEHIoTdT+SCuF8+w2nZun3cduawnQz16zOHD6G5yLqJhozil
3rkGfMHHILB55ZRth7RN4DCqQ7b5wuAHocxlzLPFLIj9yNdn5uSI5pwAOiuER8v8TLXHl08c8ywI
/H2Ib99XTdg6Uc1YG8hGLajfVQFBuIZt+gvf2f+cCL6VH9LhrkhbRcU2Nl/RQUW6MY/koTQekAlk
e+GmS7CtzmbbOJtCF9SVJS1U4kn8Yu7YRsPZfR4qws7b7xXnPvza8S3K6JeExjittXEP+ZMq7bTe
wDEYoegFpnNll5hf0E0y1Dpeha743ScIAjwGCrnDIIWkNkNsrBncI6NmFsszzTCh2p/fS4RoxE74
KECQhxCI9Mc6sL8s19nEhvGx54rkSlRPbVfWodmX3ZGABeBaSAhaKa3BP7V+5VOxbzkKbxFBTzjf
EOf9++lgR3pa/UfrIxncL8IqoNg24tdT6YHJW74Fs8qbKnMq3eBWv9+FQzQdm99Y+bVVozO3K8Q3
2ZpbGQ/QGe5oAbucnPGpJbBnRn+U8lXLddOkUX4LaatEvop1nxQGwD9k7xUVEKkc+xswbNJmy8KB
LXBvXfSBOMEbxs5Vg14BvYuNtpASNGg9jZuHFPDQ8/o7KLbYHvOyDjRlKwlWKQNGOwyyZoNtw0JV
qQsZsB/Y08kzjjvHcqfKOLgd2CN3c5D4Na2FKRhw8XBFKOdtly6wi7xlnwRmQFEDcG2x2yqc0Lqb
WIH8VKUwGy11WDWcZaulzN/9HD108kKNCRMlEGXjVi9RVu6yOFIcTUwXRPfjh8DhO3aRU4O0fLrp
6Kfy7N6R8IxmiohiG6qoaG5JxNQoCw80EziNm0slXA5Uk5xGGznGhQC9wBGH8Z0A8ezvgc+ttulH
vRPoCnOVFrKviH2GJNxPLWFE+3ctVjR5Otp8YEhzCn9iA2ItSmO3DAu5+P0FpKPwsSwV62GuClKh
ZVFEIReZXNULpFxSfio005XY0/pOT3bVkq5uztwH8Rqxm3/4u6rmTJFKctM/XDmIDhvCDSWFYgLr
LtZBEHEGE9+WG0MGghaSnZW67uhPAmtyGhWYl2XQj6zODn5jKjYPRxQP7tgd7ToFYW2V6mwvqFS2
J//xAuMqQMG1axH9mvHYE6ptZ+80BM9s7ncb67hcuQLApSO5G4ccQflEkHscNRdTRKYz7/XdtMFD
mMN2OD8W0f0EDmtNGyYRB+kJX+Fh5XP1m41UhVLJGCj+8nG2r54HJdRd7wMgxe1JnDXZs6QgMShd
T7dWP6/I9gHmLmwzftjy0cVsPHRQNUxgj7FtIZDksggh3XDj6tTRR4oOwes5TajNdHY+19N+yBdF
evRs46z9IybREldTBnf8nOhevGGhSVIpKuWz7LMtcg/xHnIrFEdsG0SxoObaSqu8HWAhBeLBW9kX
IohZ3KsgiTJ1S7+OdUVUxWk3x+yQkUdEv3lSBKIOJTAXRsCEdGOKIUjsusLFNSBcZ+aFfJVNMygb
o1FQjAAGvTL0OuAIZ+4Q5eGHsGs3AV7FbV5fDIKkCRwdXyioqtsSNicXKVymslIprX86rOrjULkc
OVH/isUrQ3awu6d8d8Ihb02UZs3lw6YecHhHLTukF8qOs+qvp/zJbGa8jH8Q/ysGnk+fhDAwX797
1p/+C1VBhPuVePbkKaJ5yuoCFjfSiiy/NZx3QFndxwza3ezEV5u4abzAFPKYxDqbAug8h5VryKyc
BOwGPYh11bocNv/BlXp+dK/8D5pr0KTsg2++pHScdHFXSJE4QfMl8Ymx3ung5nSfILNF8nmiGWiJ
TvpFtvYGBsZ/SZOEWjtWsquzT1RCEwajAuXgoVRCAixxDBnWjis1VSrHQP5KcBua9sFH1HK7ZpC/
nhorXiNQy/dZSmNbFhruD82iPbgIkp5AMwAXsBG9OYYU3x2Em1sEKRnqJy3ZhnP55aD2XpTAsQrx
HWz14UwTeYgtio9qn6UWLq2RlMaVSmJ5RrGcFigQNKBANAToDZv1TlXKnr557A6yyRnZ+NtPjw96
yPuALbHbTvjk+YvGwGhzsosbcn0H4F6FqMTs9nASXRyKjwbx8nBKn5z3aWjWlRP7mOxWso7T1wsC
5V1A1brGoj3PeWcMHsYT3Hl/ap0+AHKfsJmX5kbuRi0GPk8/tUCzcHNRsu8mhlLQ5MCXucgrfBva
KD6Z1ZAzACBnLyp+rW0TrpVPy/DQf4C4cToA+iqIMp9WSjKumkxjAZvn5SjCT08mg7NtqHL9II8V
80YCeYVNk+fWSXwO5ej+Hw6sk83G79sJkSkaJN9EGQ2JLpCb4twlJ5VmzBJXpE4jUHjkfTmuXk3w
qEhqaKym4N9xe9xi94HWR/PKz4fK7lzCN7udisEQ8fuD94Cpk9uvu0tmhJscCi0YM5jqydy/rbnS
5Wq8c6VVpY8J11F1cFH3HjeIVCGsIHFk07ZcTPVgzNaYmjM6daZT39xfreYrEjD4ERKDJp/ry5jO
D+2qWglR96PHbWkNgeAYCme2YNLROQLn1ytVfJu3CbRFgcETy+g0ML5prezcjalKvSTOxtuzvmUY
F901YYMwn5GuRmeLgvMf+gEJ7GVwFffPMkcGC96tveW+M8ah5Qv8wd1Qm3ZIG8ChK2c+EeknF3RB
y7E6Pq3rwY0mETJ3vceEYKgQ+EPMLZIdp8lcBGaafTqUOOhai8eHnefRIdgoHXqZJVW4ZQ8Qtldz
tC263E2Zt6ESAJFLYdD4g4iKDz0GbYSOkocxfsw5Ur3hfzUQ68HjKCyo5c7QY0ki1VHTz3VcevzF
19ybkBoxFHtteFJa2JMTue6/HXFs2lfVxghe8MXrDbKvdQ5HMeG1LVNY9PgGQiuy7KgtzvQiHR4P
f3n0WhSDlK/2ArCdIbtriJ4bx5mkN5JqwWJ6Jd/Cm8WzNgVENNVUY7lUNl7QOFh2cEGDdu/LlB1b
7ljU9t6SBSNkKb8CCtvSE895X1JftoZ0C3zCUtTKRZRfSRuPcD6l5AGn7mtbCpExrcuw/2Ihq3vi
BvtggwAk0ddCzNKp6GLs2rk6xd3ilI0s8+DNjNT8F2aww5T13+SxirYFcq1BSx0Yn4uk1ZEADdJo
Ni99PFGj7TRBvxM9fzHh0UEurUg0ruaS9QFI04Jd+S4IAndCzRgiBvOs55xhPf9USwXyvRrmYmZr
XEofgaRmpBk1ieF5cX+pmS/de5wxhlmwLCbmgQo0V2NaY+hqA6Ms2L6W/wxhh18OQNDcJ05W6rTc
a2J0KmY9kQUUCXApnNpACFspYbh+uhhamEs3ijBsU1x/5Pa/9M95KHhyG/NtFviDCzcxoMjsss61
BnxyGZC5WVylPmn4/tMNVPiLBFGLc7+nst8gCrQ9Skt5dtsl85X3OvM+Fm2xbo0l9QHdvDDmZOKr
TNayMAdB48sgfd/b+WjOYqyl5it4aXxPL9E8ygbNLMKGfBb473A+xOBtVg+C3J05fC0I91cZXppl
RZSU5UB6jj4erEVrraFC94jcDl2dHBoppdWbrozsApK4Om9RolEk3f2TGj0idCYY4XjdTBjq7B6K
oag0C4zH/dGzgeXB2K9iNUL2T1TwAUNxqWil4gmDEE23Qd/koeOSlkKTjAfqU5/CigPAl4q6zgB4
FEnhEsw4Xi8j6SQcWTlTtO4ONSiQ7bpi8UDIOv2ieMHnKwXRxFoZbNDoHUmK2grD40Kzh0CmEekc
PU6ynSmPwXXUbeIMBU7ZZJQdopwTZ/nAMiw046nVgJQVm31QhflqnpBnFBaMkEQl++DjBhFueyNw
NmxC6yLRqs521w2tq62M0bJN0+1h5w04pgndm8tj3z11G6jEX+Apk6XJ6qPhWBeH0vmRAlcAKWvp
l7wghoWEWb3jcb1mVBJS8Q9wr9/HBAFqDaTzkA/oorxwB71n+i2m1mTqaCLSu5HxAnZRxMqcCXNc
XyaEogltspqFrdPgiYOyj8T0ErfP9Ye+HbFEjSZQSWEPdpzOowOcF37ggzJUrVC39SF8y4up9c2W
x0DSpx6q3MQHJOptanC0/9GK3/ZmDZd2I2oSQzJUsFExQrzuGwggIXwhu8H/L39C9dBYTIhogKTS
oC+hY7lV0Se6H+n8TcKUnyi/GDDyyJE42/xfJfiCwcEttbkfwMW8/Kw+LFveIMYXALCsIYjvt5yb
oI/lUIPDpjO8+ccl6i23sGh5NyjpxWn3GKOJ94EvABKkjevsjhtfqRGhJVtTvEPEnmDU2Km9vu7Z
SC2z4CSqOWPTM+W/TSM2iqSqhJbTAaQOA+BIPZqr4A/t1iDoL3jWAd6tFMRfkl7MocW8prWO6HvX
TWgGUp5FWwCHsmnuAaTSCGcMH1T92kArRJrci6CrHNCKG2vs43BCGeSs1DmStxVabfNUrxiVB7As
rj3OpmUhSmhLPk9JoMlqXBWno4EWXKLhd7MiOHZ83k+aGOLYUzTZnDvP35PsbF1ltlmQFfcK1Bp9
e98mknKRrHxOPS+jcq0DYWfOW6IefeU/LjXwfPvEZjnZK2usZn696BdglUD1m+zlvrUMJwp0v9D5
HfGScPFBdukPmgkLDQFEPQjC6CxHz692AImJTX9iNCZxKUYlk8ATm11CV4ZhFye0UHAHVG8U33EQ
IGu9UMnVouNQe/pkkUwapSb006TW+/tCn6z04blsMFOdQwFL56tuVAVAXK17qW16Pv2ELP+7cCFQ
pbA99C0bN81IpjIcLEffRUtlUsJHiIsVy5uw5iSxWc8sk/j+T6NYcOI2VeWmRU9i8VHEQ+4pBaBY
u1BCMu/1GlEgwwki56gj7X9YXLTkRVFkhUXCPb3jqMuCGMWg9jwdREg96pYHTxtbVbcp4Jaf4feB
/tWAdHeRgbOxejiwkBK5kGNi52siiuUdLkzAfblSuXdjDaqzORmFIk59+FAA/TWgLlgC4WLtGpeP
gvaZWmDf3OW/JnInx47AP28iHKHbI5cnA0x4mM+RpgodfNkkQMNcwrDFM6WwUN9MMaNEXT25yCQP
1pKQQ1LkWHkad7UI4g9Pjo906XVUyHwvNCMkZG+1y4CrN9/M7UPPj5XjFWPMVBJzeddmvKkKClN5
To5eiKmVSW+O93hIeFJpzjctl60e7GE67pZsbctx0SSrA0VNTaD2hdqirEPVEapj3QhVv1lLYggD
aOFGrlGTsf+5L6vUZrP0YxWwbVpNq9nSRNzdZsjD1bmd2xuLX3e4LutIpBzDIpl3h6XHJgqB2+gG
0kl0u+g1hx3ApFHkf4m6PH7tl0DFwv1FnGMvoG5Wd19/bsyw9acqFmKlEcu05RRPOiGMwKFKE0+t
7tLaU7GJkyMxLGIpgXhtieCo/TincF8K6VZE3ltQMewlPAOUOPXZyL2O2w5Jgqoetl47urGpQjJT
DamVWJbLQ7SZfiBRo22RabRsXglldWQZdGP7lx1rlAUimwbUym7YJb2NM5Go7IwI7ZxsQwP5tXrf
H0VTk9/l+QKZbFMPP4JdyKU7570YIxehVui3kqQfwb2im7GZU6fg0YUzS26NOmj11kYDZNZirD97
LATueNxcE7e2E0xZqOpju1x4fjuFauRb+1FvlymuhO3o3MBhTGfDcBZXWTiWSvM60LEEQPHauPop
PxecMmMHzawZVjZFtGkoW+YxBEQ6bYu6XSMc3ogFSISBgmUur20nuM2yh5p2118paVu8D9Rq83KU
AcZNazDhzEDWLM6NRZxq66QzQfPZ0JXweSVlAjNr0KXNsG5Mp+2gpnN5Fey/qykQoABgUUsuj/JC
X7H042GF5SMlQzgefmLRMJUDXo2vEPFVgokp1IaYIt+hULEA6XFmEuIOtwVXRGp3FfPP6ZFkoYro
UiV5rURNM7Bg9sI/3TuN2ykuCKILZRII1Qjh1CJI4VDXZAFVqBVvLHuvWvqDtjGIKmMMGbbsFmZW
Ya2oWfWozQTWMT+6z8zgUI01h8W8uNMCzjpi7jQzt8v09ScQvL0Sssihcpu/GsKFoKVux8vjQkp2
ZvqppBRdUU2c8+diD86Q0ygtdM69ba0yVfRG+zwAeUw/XwenSrlYMC66sRnqkOLMUVi6xju5LfhQ
EFMBi3ACyPcyDEg4iyI2zTx7Sf2SQF6k5e1k5441rAUXmZmhgw/1MbpvqkHVwvMtZ34HrLmyPeK4
b5ZnVGayBbCruEfJuOMygpeYm1HPQi3CC4g20ud6e2t/W47VYguVFd107KIwPPzsAXIr7ZIel2Kv
tiE5amJXh3MlUPMnC+bIG+26gnlL4b4UbakDOYjD7sUHYH/fKxmNPr9t7Yrf0FHK2LKZJ/M1WPIJ
B2CGl+wQwq08+rkfZHlnj6A2UcHkqJ+9SwIWP9BiBi7hPerXaQhb+y4cGBs5YjvzsjKm7+Hkn6AD
TPlS0brrcDGJxwkykUlI2BXE62sNR8Fwq9wE5ubbQUoOQVCL5wMs9nScTYRPig9YZv4HR0d7qTb4
axOIev3IpkkDYFkVYaNxythOlJB9L706/i0j3sK8JX2nSs1SP2cevtRXEc7wrUTtmwo1O9DqOzSv
cfvSMHue5zhU+akrSdmup4mnS8wVKC+gjGJFNEGsc8FtZDMSnp9Xp3V5735ZzyCLnQa7RBRiVzAe
HJbA6fFED938IdH2JRKsnKE7Wu5gFwFvdOrYaC9+ax4RZR8kv5IOaOlGKV6HeR5ltzIeC4kfkLpc
sXHMucZ1KSEubd6Fxs2a4YIa1qaFkNhtRtXDiGpt/VOVTCfNDcg81q6Qt6T/czL/nPSMOU0Zy/LX
sprAV+j9KScH20Vyet8GaZgcADi4ejAF/XE612OyLliAgNICOxv2hezQbECoK42BKof+YQrznCmh
JWYBR9EScRfHJ3XGSNWOeUN87nNXPlpDo4nymdLM4AygcsQjnUiTIALQOY5mcW/G9hQiR1jU6RNd
OTSR/tsXPgQrfocucO4B+CM7tT8TTnsvSvSraTZQGrmeIB6Inpe/jiHtoBOvl22RHJWKg/C/a7FR
4B9unLSdckNhpjqHJMpRGVXXIRBHBxqWDwGIYD8BG1WdpKfukPCgESb6fbXakmVHPai6Y4VBbUL5
w3pKaK56ylaUQKudjOWjTz8hzN7h9Y0EZB9Bhjtqw1rI4lUiVJnvY4hURaGRsB3bezivoD3ivxM4
nsjjF675YThCcyArNoBe0ilk2CN/oK2KQdMvgniBs0pvhXsYaYFwL218jxF/CEMWWr0ojVEnPBx1
hoSFgutjCHAvGZhREGsXLih9hYggW/JIBC7vnFmNlmtA5Qown2r7R+XCwl8vCbEN06S8f7DD6NYN
Zvbbgoh3oXcBCoLbMVGo+ZsreepgYp07lB8sgHjgmGLQPvGFkQ3fnCB9EjEljM6J1vleV7QZkAcD
mUUj+WwP0/TOKoh9rk856OXvhs06afVtSDOLAeptPDcPd44FfLEv/46YE1OjAvNtEp9Hzk7lW90O
2pqXoM0rqc8d+b1ll8B2iRAuxKNXl23sluJ+N+ZmN0Ul3OTivxGs2o363cIQIXNSs5wCkVxW6/60
+zY60sAxP80cCvPTJmrmvs6a0K+DUQ8lEkBVr4LK/j/iFKnUa/elEm+BMHHcnx4vdeoBrt6f1iY4
BGwcHkh05Kmw5GODxbRJbyw6FweiU9cl+4wrsPiho8ICCK3FBOHmD6Z+3+cLPf5B1WCdhzQ/T99S
Qsbd5S51oN7p7eEWIT8I2rxEj2JnRrQ77bWeBswsIdeFLiW8CBwlpNZeD3f4gO/RIJF7Mqb8rzkf
NFtlGWr4PumVcrZHWUNVpbx3uj6Qk9nRcMa/i1sfUHQBRZc4bRoaqnHQsvB5f2Bfavjoyor/WZ9a
LVtDuk++d2cyIIHc2A3Bmhk9+Qj0FTtHT7XTX28+2xOyAeWnYf4yzSIRTUD1WvRg1Kp2To7hkNT4
mFaa8/MDFuX2dVVmArVMVD2AJqzSn64ZCybUTKAv9cN13CHJLC4Qt9wQ/ZAQMSrwvG88MS2mo2DM
DXRSVRW+ffzkcS51zVoAfbdDacm0FKprXwUxoM4OMvBn4ga3QnH0wB7o1QoLA2n+dZIh2BRdRed4
sktDTyLzl97UWvxWvRhqydZB/4ELv2JRLpjfiqB6Ky6Q+mKIRey9koE64D3NmLt5X1emHhVLtyct
Ld18z9uS4PQypM4/+i5E0UIB9uu2WHIYIRE8E0dyrPrud31hjaNuQj0S1TW0eZMjmUrZzRYhBvV7
uFS0t8C39lIFPkMD07SMjUbpiMSH+VqBXYMqPO9s5MCBpaLl26m/q8A1aNYJbAogP1mb37dMqAWz
LZKoV1a5dBPMitPYQvbpNqn8uCuA4NfSGUjvWkCkb+smn3o6BTvPj6EHDaVExxnbebEZzEzR/xa0
oHf1GsEIwLC7dp6drH1/SskFI/RtlrFwS2RUAuuaxbuHss6KSZ7cP4COzs42rmiXjnxiyWSnOigs
mDgGyHByKZAtUTTCK55e1AOdHA6mv7eBtJSwxO1DHd0ARzATYnnc/6GEi83lAFllqgrOrkzYeOki
sSMF92B/DTPs6S5w+hLTsX2TVa5bUCdT+zEvHX9XwF2lhxp3WTJwVqhKaqz5qqK4Qr5odcdqISjD
mMoqy1q6S4tiizQt9LjGhmWZuJFyvngOog9pI5qRpKsH3xS1HllTldzSg0uzK559QMfzzllkOHzo
1NL7ds30o0newDBBFBj77JJcOm9nlbdE74BUSRKlqTK6V2W4bj2d6OnGAbGDzrJeQb5tG3TXimnM
fxEUBqb5Mijdms47Ytstl6t3bK3Kzn/7rcmx/WtgWHQrupQelBTP3Dr+ImSoqUFDplbBa7xr2Y0w
+NHUPVhGLsyQg+IDQxvxlsTQ7zhBaiHerC/6XSubQOIeKEv2SglQIeCduFY+PFIiWFo5oaeY8Y7G
/gfAsu5lRDMM5H57pOqp1lIEU/YdKKVOXYcu4Rq5/TjiPRTgWmfnvgZ0VoXE29pwAS6JhuFHGn8H
52alxYPFMcZA278PtwA+lw5xN1TJQJS10X24KJGzLWj3smHagfFbB1WN26hDf09i381Xp6oBnqDq
60Qbl+wO11wB1FaZ4weL3ZNqfilRJ77UeEsOhofaKmQ+WewpuQZWMB11IZ1yyyThOIicwK/66+1D
I+hrMebzgipK+uxbm42TtC2a5MaIcJDr/Q3e4UD0nYHdGjioVXCC/TdK7JjZ20mil5EC3KRse2CG
7r5jcbQLDkX7mT/Hw1+KXRZMO1fO1OGzT+hM0bFRbpvFpPZ0ebZKEvs6T7oHycD4RSsxVmt54q/x
4d6/1I5dyf/4oUfaGHM64EUUcajUjYNoBR+R3WDbjudefBasZhcwqEM1JxWwRSl6LE6tMEOKFTJW
QyWhYBhJ3PqzeLRkZKqTloadNPcI+aWCiIhHt7ip8o8hSShMQkSNSn5In01hrJ6BhntyR2sP9KEb
ln9PIx5xspad72TT/xYa89FtCEo/k3OJ14AoqNRXSk0fyEbvfGB6cxRwAo81qWMVla3gX01Xz+Vd
yqvOjeE26t2eJTYKXezo4NezWRu9TSzofnE18RmS+E7SbJIGfKhEneIyQ+pv6TrfKiGJIJe/XNbL
HFd/R+zOLbNgKQPbPEoZ8qLMhYYtupJbqXIg2ZsA+i/lGdVqR4L5vCyS57Jcw8TkshKNKProYq0c
f32IMs7GZ+MtZ5mwzUNziD1FlA25N1ghtE+bIjomqeUqk7NRv/t5aO8+JOYxAdgDRjfjJUzeZNup
347HtPcKzOZHofzAp5UJokiyvKWAdbKxrMxY4Mwl7WHCPqbCo2OTEXXA5rB6VhxsPIHzMqjAoLb8
ZrF4PfhVy2bJcFNmU3zJ9mdI6q0tw44mf3CUxTH6oAoPPAZr4dAjMqLq7ifeRPPbsHBnApMF+02L
Z+sVSclSd7ilY3k8HRMm9miG8zj2RKKzEIRPv/wsmyi/L70Xfk8uo7/oj+RTI8rRGvNxzAP067iV
r/3T47INbGImPtCbBL0EAqzBvJeoMLNffKlyDdOJP3rvOgigXz3hfHHgS7kUCUFFEHrFRDQ0ctZw
tC0E886vTctClAOtXg2QQrLoFrL4bVhqI/chnDyvCtA/ab1ib3YfskJ6mAL1L9Bi6IYGjaBrANbp
RCL2Q/t9f/zhscAUdzou4Fc6uTK98MmeQTWIU6IGjRFZ2lg9ZBhfHavsf0Oruavni7Ueq49Ftj20
0MbKFEcT9UIUmsmw1GRvjfLUO3fzjpA4DW5w2UiOzL7d/nfMd1FomiWPOm4K7gWsb1iIIVUozj7r
l55x6YNeNEk0po6pmJjZehRe/dmnC7++mg0soo7Wkjtm6XIOXottKrxdKEjDFYl3QB+2Z5GHS1AS
OOis1AQ+MRbgFlszbBRgIVX9g2g/98704AkP3Y7/Z8HwEdsPgW0BdaerG6m02Kn43WCDtS5wDzMo
bzeu4LdgC3YzBRsHCMb7diUKSk7Tb65X4pF6BuD9ZMc4m25zbf7PbueQ+ECcrgNRUsyN/SH7rct6
i1HrT+IEX19zDHdyjx6QbssyB5YkX1RtQQKudnB+09OdMXOEzTwn1fKA394oX7xWKvXVkrgoL9JT
bbK43d6vwK3hLlL8aq7YJMhh3NTOmrV/F+6B7VsfrMpvMH4dNwDEtAF8cNT9VK0OJ8vGlxSBCfP3
kMx6WTIrYZGZei4vXZxM0WR0+DotwKywMGS95CrFIK2a7/TphROBYEe+kcC1wLDlo2moHxP/1JnP
VjyjD8MaFFpfDzfdtkppcxCjpZ/TLCCHqlBnrfnMk5HshCupjmUCfcCGIxsC1v0PnuYl6sQOQTIL
YlhLos/p8Fn+xQTWAM4FqP+QvWAZAbHwdzN619wxYgDMl+vpJUGIM49NAGHi6pdeIiiS3Hu/xQkI
kA9ANDhVlelQfvfekFDUvX+HXpwrBZuV0SSn7lzh+q4G0F8nXpkF7n3p+LD43ghZwjnwhAIUhD66
D0eYEnx8LxxeAlKv2wb4su/hvk0PmQnEeuxkppBuuotQ0who62w1Kimk2Ul8ETVybYJKM8y7Bny2
/fcRwt1m96nvycbx0APY7lgS5bTucDD3j82yfE+aJu1HdmEsvuainGUkJdeu4JVESOZnKUb5Ws+N
yism8v43C15mrlqwAXijwc0EAVytXwjTc51lO9QgPGRfLE926zjrJadoqi6//k2o8j8Y+IQgj5sp
ka3zqpTS4M5557+ji40jWikreXjbp69chOVIdYTfPLaJjwAaIDHDn7fy1xOvSMvQ0Eqxz3wcLZ2S
fEi4JDIVbHirBNvEaGJlThy7PfIXnnwOnXQb9bhJbqPdyJg2Xg/OT2H3CLq6aeuev/p2HYoP2ofz
PmM8X5Yzf3n24Y3isWQ9nJFj7dy3fPfc8fZV728b2aNAHDBowHPzMjfR5ZDm4J5FzO8JvQjACWsJ
K1zpUqjLEOWXxmUACO8FYXzS0lFeIzp1KEjzGJy3qToOiQERvM1bxDmSn3h/4DMLdkebE+isJqog
D9KDviTRORVd++EfcwWx0oU6rU/w7vzQxsn0TpLTaNfbYF/EQ9n9/B9J7KEZAwbu34OT8xdjVMk2
JP6fl1W+W0lfCMJwSO4DCWRzyKvEfD2TTdMtdc9S+AvjuPClhOo4c2D0lgUuUT5EiT0KmXl0mubv
zi+Yyvg3rkF95WMMmkQ7YuxPHFaQ7g2Iza9m9QjlAmvpHQOIQp5I5gEgldQJtGb7DuqnbdijBJt/
r44tTnX7prtx2SI+X6194DjLVPi/jZVuhWo8Y8DJH6SPA1/Jrr5sYH3wyEUVkrp1Stp7OQkufu3A
SCI3iHJ+kicIr0Zoz6+2p5G2q9rEyBGZbATV8byC4VDoMuhRT38a+Gk5o2z45D7p13EnAPUTJQWa
An3/+gywSVXohsARJ6qXbjF9Hpnrhp2w1bcjCuXwJCle4MSH56i4xtKEEW/99quJa5Bf3vtloSrn
FsDHVhxfleJMXBQY2XBIzK6nM7cKewsjkC+OfwrAnHvF2gylXeAgSgdp5J3dLdPG4ywnn0k3rUrD
KLBcb587toeEYQ+11Vagxi0JdCAPOrjRDAhX095q+xOqu2OjvTwfkhayk23qZTXanvDN5p/tEr2Z
1nUy63EhJNLF4H9c6WBuxCbicXVElcK8coV/cEP7RigWcd9UgPYhL2SsZtRLxYEkNg83rqORnM8K
x0mu0K34VVDFhUaKOmrCUYKLFzSPlxAfLAzwkEPDf0lYRipOvwY7Z9uXwwX7BJKTYPejCEgY1uyl
yszqvqn2ID5/puI2TpClltMarXejYGQX02GEUbRU093xnVuD+pfN7038zQ9KloWSxIf0XnMMn22H
fwokDlAYS1dGjdzAu+awciICO1C3QMRFBnUY2vXw0cx7ahLEkPVTz09r/YVdY2ehAPpRAwgPUfux
R2zZXx7b+hNju/xHOyG+eh6BkbDE4cc7OGT9fNR68QE6mNj9VHIdiz4R5EzB1iDKsXHljN2py+jW
nBxYVSBNGsRNc/Xl4nIanIScJsWVkUTRzK1fP5KA5Q+lNASIi2WevavLP8kzDW2Mq1VHXyQAcFWC
LC1QgHoBRM3MZSCzi/IUl0P/uq3CtC9HGtBKbxTfGohaI4FOTEw09HQ87qZ27qxHuJcKkVHPzSiC
9D9va214LwxKIWtg/bJcP39otSq5C5uFkVc/Pn685BXu6og2km9Yw1KM02tuDZtPdV7UnkXPVvBf
Pt0UDHinS8xWdB5M5+Nqy5LX6ooY8PSIgX3ri9WPOCZG41hsuwd8s1UiBELmfVeUv3ywoindvxLa
eaLlD27hAsGA00gJfMrOGO05YyeJrvzadiQBzrSAYMc46fLIU6yehZZ6WrOHJqOD3/ADnZgJ7dGA
SHKoiYJUvr+rgd3kyyWLbbdw6RokoVd6P4Z0JbAAstXx3hcW64hbgHKG4zR2hQwVsHtommLkr1yl
k7Q559AVMfojeH7wf1yVapnXDul30kSEQGvHJLOtN4AfwBNEJuePQciUWcyL2cblcV5XWUB5NWzd
EsZfts3wIaVJrM6PBB0K3ltQc9zClQ/d6F0FNuwFCgeOqUtsDAcL9IrXBnDN1egfrl7IlD3abERm
h2MTOvgQe1flRv1/WoEtlz786rsd7uDYKBxHt0oKe8zwoetV2tLmpqiizs6jm0GFFqrR2CNZng4E
OrtiOKFVdCVVoYyx0CinqydTTVBK+tf/RlF1+5sduK+jUfKQb1qkIlPlGVQFADTwsQrl+oUti2C8
HEotFXMKxXOChGTArUEqNCT8WyA2mOZscSypGCo73pRTHYI+4Kot06LXBNzavFPoJ3UTkIZF3Dww
FF9mTRvLjeFA7BBwNnH9xQ7nzf53S4B3nnYPNB89xZQMMQHckHDomyKOzyoPEm4X5H+1IpPIA1PD
8WE7MN+QYwN2gMoScgOJjKnwS1RPTOxsLKNACSI44aXUHqL8Cb8D6KGuqfCvs8gOxGIMbWmnWTdY
2CNEemdx0mSeODPQK38Pnkx4glYRBnzQaXmpBuIhgPlsQUCfB7kwo55fIl4R7RxIYKYIYUbH5FX2
oX2RfwRHea59d39Lv1wWAhOv8MIBlGe/tOUOu7b+csW1tQkJkMXtf5ziSAtmcfn2Xf1mE3lpC6/b
dRogfkN7tDisJTsKYOYKI3PAX7+RqR5NsCXPnQhZngMeT8HDQi2bdh3ySPpKOCJRD9tJHef9z+aU
h1EqNCuIYUQBWV6fG+mJh+5SDOYTzx7oOXZQdODLCZBjM1DfGfsLzknnCTsEsPcgJ4EmuhTeKICY
AaVV5VJWybVlaPEgKrUM7KioV/WaWhGQY/LSQLN01haMDKYCzzrlnugyAW/w7J0yloswklTBwS3S
Uwzpeui6mgripFJedkYBasNXbFe1rrn0tU2N2TttnglnSXjCUtqA9eszknEx/U+VXVrSSPBrEQu4
4fj31u6OE91JTtjmHED5cE0dSw4IQLYVCV/tDS3GjFTFtTDdvEfAJasE+admylcVi3WxLRzoC3tl
1SDiy+oPWwc0Cn4L6g2mV3oeQ/3FcFagvhKKK8VAKBicQfgM7jNBUWM4Ekf2gdoVHFmtffycIdZ5
aJM/fPAOB8/Oh0V7yDwP2EXHZUJzPVNrsQwxcd4Jt5p0ym/jX2KYzYAKHCkq1MkkVG8x8ou5EsN1
5iMIMx+iAaNvHFwpzzDYChj7F+y1xOuoYVG7PgSNz0TTdgY3fBN1T5hhtfRxHBaUqqRKJIMKEVfg
QtUwFFonDZ07sREDDoY7KdTiSmAV5iQRDVLH5JBIEk60TElqBD0a4X3CJKVVzuqrRcMemKPsj0oK
r3Rzora7HQZ54/pJ8wGdzywtlSL6yHdx8mJoH5nHPp8OPNAGBAiG+G9OEcggcRBAa0W9rX3otGZR
4niXHVJP9zl9uKzvW66560ze8Oh5vncnldncBnulcWei8RI/+D4Qgxoy4PvSdVzEJcg5xXtrcacn
fwxap3sQTN3WqLiFJO/uBUhtUvwNL24qQD4tJkmulnFfWT6MZ/U/NNXWgvDWQqkmG4Gf7N9QePlc
1Be15a9eZ9Oyxx4dtldBJW/STr+KqepFTBQ9W+2cK/q2dW+RvNnVgk8K2MpmLJ8Jw7a2DlYfYHqN
h9+KfjDi/6SX1vm50i9N31taJzEf0LmXV8jE5QOn+J28Kgb/cf2k6xEvL/+4DwTjL7X6Z8RqHUeC
Kczd9a97cFKCzml3T/lsWk1mX0tfS4m0UD/QIl8EOHe9KYUlKGmAqLVFQuQvoEE1C+l+ssmHCvZB
jdzpq+WraOjopEH8aAaRx4mn6CRWPBT+ULwREUY7cpax7pCcHB+A6xRTgIIzjtx9STtLmAola1jE
HsrTqMTq1fYBOAN3OCrF9EIWuZk6/L+gBWzcHSXBgmDgPS0P2envCnlqDnR0i+ew0LqU6C7OC8lj
LDaiRXaBOWNEl59rabaP+gHiH27TUX2w81OKjnb5WqGMvigxwdIzyTIEjEfTb3HW0a9wypK9z9OO
b6NNCng0onAnDH2lLxpiNniBoH//q9GYG9NsOIUFow3d8qB8xzbHaqFRPAGlLrljQrSBIpFPS/iK
B1a9XuVc6svUgI4VvdHrnUHzWiy0l23QkaIeRynFViV+FAwt/YOxneFvkghazmwYCQvJ9Flthddl
D58l4X0hE+yiJLQAAqrA+YNi/c0EK1U0DY/pNX4c69IgVBvq5mqrs/lvm11u+cj60l7WQLLBqh/e
gQv3Zq07+oSMNoyx9AIOyCNrvO0KC4ex8HaAN3f1Ib4fP1jkBTKrKdp9oSKQhQOXDpPxO9+22dok
a/x7niDsbPzbX9T/FupoBQa0BtKlza8nx2MvvG5O/rFUKRKuEHNFeMu99zkd/yFSKIKWKNAYiUeA
4vIoo+JsYp/ObdnzzF1WNHtTQyFto01x/RHCqUj+uc7FK7em3BCPows1ssTnGXZSNKEdMtvy6vDU
oMZ6G+ceJ2EJkqYbf19BQVXL1z9mGkA8t9y9V52KqVl/nVCOT/KuiZt2J39kbmRv9Ba02vhv/yGt
geIRj9XfYayAgB56n0H2n5x2FVGBqm6QxyizaUT+4eJd76paZIx1FYYahMTbAV6JVEwzeY+Dfsbp
N/i8eopLdjnue7aNEX3VYQsfJd6gQ4bGPaAnF7pbVaA2Gf0ThqnIjL4QwGPUQcnpOqzIXoJH5lL4
NHs1fjcuncA1EBfnC+7xfA8rFoO8xXPR7LUrDnEREZwkdh0drTal7ppL1JLwm0xbaie2t4ng7tbn
A8G3NKIXvwiQC4VkI844DnfTA/nHWXRRHSQQVopy52U7DhkEaZhy5CUdUcrTi0TI/i1jhZeDEjBZ
+Dl+GpGxxghemT1FeUqkypzIYpSwpxtVoogQUeyP21LYWztJybeYxOHI6A6XPxhQZacQiSNdSl3z
PVNjwR+7KZF7lqybKP/+z/69fO7CUeD9TecPs71DDYszxZJ4u1cQl/4HpzqAlMFD/wxBoSmIUKiI
8AtwQPJUyUuTFFY5GNdDU3YbN6WiwzBmcnmeWhkSO9LMwNGcqkcjpw43rkrNmKRWNewj0GFkvO8b
bl9lBhPqiNGmshtbDYp8ulIEdh7NidWlzUOFVqt5qjidi4Pi+iu1BB3v+amTDWXr4ni39E5rlxou
9i7eX82BmULAwW87+PueCBP82IKs2BPajw+ei8j585hHg7+EVYfEzZIIGX/nuQ1DKYnCbkDMzKF5
7d1ZpzfbVrdd0qPvCZxSH6CqEJjEybi8bkkOD646tMNH/BoUXiUwq+YkcZDWzN7JSKTf3WXNPPDQ
uEdPqhj+nFpF8wZ5ow452jAkd9BXVEfEOs04npPQgD5QcLHHGml3qPFfJl2CxILZfYPg2S8o2MEn
b38KthJs9vbYhb/QHO5ezkYgZsI5ieNfyq7cKNhJ/3naIzEL7T275iAnLSANYMfl9FUmg9Go8z+V
v0FZW0SumcQ1yNfQBnliLWK7GRDpCRjF5gIbI5/T6QYrLUX4AUxjHjI28iHxtC31yWmyljXQ/uj5
JHCJmFq4g4PZgB3NaSySj8H4pU2yZ2fh5ycevP+tpvcsNUxaTq67cP3Sxu5c1D33tIg1FpqtuD41
cSoGQbxt7ZuDHwvCIOgR9RVA0PFmp12nTF51n/AfifG06Iw0wOPTM2Mcl3pNY7s2O3a33ARTRqyP
r98Dl9oA8zzBKPPj5N729h107Orjk+0r9juFqrM+BeIKf8UZFjFQtvnRFDfjrFjVhAcGjsLjHwMq
VRxQPvloL7BnUhlYkFBshv7dL4eNM8++AFmZ4X4BB2b53YJ+ehNRrf6bvTm8XaSx2QLB8BUxxOds
fhItrhBPrM9sUYTYLuDETL/wWylR5g4bN7eG1v4MogPoTA+2kokEKOAZpTenIjUtcX1tZKb8gbPL
WRwmCdXwTQubnp8ozRkcVSTYMkLCrDFDOY7sMGjm2H7IUeGCl63zWrLY2awRo3hqzooPJtUg5qPV
hWhkA8C357lCqL3QhtYED0tWn7XS3za8B2Fh1hu/CltGOSAm1jr+w2c7PgqGeQkWdPCjxXQufKTG
rhUG+0npccjwcBYTQa9UwP0D0FcvGfD+wzojL5wPg1IHHsPSROvcfH9C6nocWOB8U50L0I7qmBaH
cRe/FPDQMB++uKmHlXCRCO+GjytLuWPg3S/Q6foY5KGa6hZ68MtWIRSDlLpQIPruYUN6VOXV6mmY
AWMVioKKht5UEjF7DGc1FX7RPyc1eFkkZfg16gy+FDeV62tFD4AUBWaTGM4XZssdSaTipslL4yuQ
kK790H3XM5q4gXllPr6u8OQVY/f5XtQG5qRTgTcCkx36iy5vKe8jtp3l+B/sFQYZmwBvdDl4NFPp
4SFWU2EqSAX3xMw3vmspwrOeRX0hmtIHfWC2nBJ53ezzLBlPjQAj29UI4kMGM6v9G8W0B5sNH2UZ
URBFO/mQ002QrgUqtcx68gGz6L56hmbeaSUYqJEJP2mhDzcvWXbX+CNl6kO9c//vMGYLqIXZFiUU
MFb2+vIzT5w3BlpAkq0La7ioLm7EsfsSF28oLb0qD3W5HNOTrbh6wZXHgXuaIEx+/fZseBmYiGAG
5o3Ia8SI83zgzhPm3wzRFG3QSQhHcvRS5MFCpRZ04eR0NBzK2GAdZFmg+311dL28G9bF1PCz8x6T
+PAgyesDZ0q4DpiZm5gvdehPwT7SXWQgqITTWJbjW0oBVq1L1gS/maf/ibt8tyT2icRCjiexVGHC
8WxTJsPhWcfFgH7viqD7idlC3EbjYNGtYw/3pV9WK+lV+SSrHHQhCT7jG+DWA8DBPUEhBFztWsWb
RJFOMHbzoO4sNITP3ujaG6iblj70S4yjDLvUyCqUdic+IcR4hUigVEATKUVZNIwioN4qX3mV/gYQ
obnhYjKXViTWxDkSQEZHur4w/najK9Dqk6MF2J69KziIp6oQb1VT72iZzT9sXqQvjsNHQnw7IwxI
DmFwsOZE+Gm/SBcszWIZQ20kOipI4DGxXOj2FdouxXN9OddTNGIctc7S4W8pvrGDL3lX+Z2gaPx1
RErA1wSybQdIq7XnsUip8t5cCzW0pcyUs2fxb2wkyKf1H9Xs5H3TDvIfxZ3OG6Y2CVziBftDmtbF
c2VwpcPCezobVRyicXe3EGeDEkCd50Fm/nFWcjaKDPnPpPsIJa/txlgB5nGARmzZkmD7F/N4YeR2
5/J4LtbFrw5QpVG5ubk1FxqJLy8CQf7F57rIhcmxY5PYwQEFht7fbhzM09KGJ2Al5yAwB8NYd+aW
162KRplUNGf8moGyTzsJo1ZStKhyJqXfPvKDXIJWWBYh85QNkNuZGD1wchnHkCBTOD5KCJ7LgGjt
HWFNuL8HPye1ojGlo7lysajWXUxHfVKXsZFvVy/dv1FBQc9gTV9ycsCGnc8dWm5g2FlVHKAlDHba
dZDhtNQYAiNw1fytoCrlf5/M68RwPy3VlP4XQtHjtjuZ/wdZ1XPSumw3LkI6ZId9oKPP9a2GNltN
gJdt4v3d7OltBc00Xl7Tud87TShmXk4tAQxqFMsupoX6L94uzFojCuBYQh7m0zjtheHRfhx+g5d1
15wePF7BPMpdDzGsZN5vyebROjBv5QN+OwxDEoNtjAB5DQvboWlxGgf4vvpMUa08TxGAg/4ZgjvE
/VcrjbzeQLXc3i0T9XQ9orJo8kBuDP++EdH2a2LzESjNUL0me74Sbqz5zCSxugKu5E7FKi6ZcNbJ
AyCamAyhWfaD7p+j+7cy5F1ZWRizWRvBPmAY8LJSDYd7E/CEEiSvLXlUuMasf/jVeX+VR29gQ9WM
m/cKSn3eXMlrKCIN/2TbYW4rejukfFnQBO+tZmO4i4lwXYNvgG/zl2O3QDeMynTMcuuAzM9XwUSj
lYgdZZNKp5wpNFxVW86fGheyn2LhKf5AxnkpwzWQPIVCi//8x9VIcpitPN7gWPNh/nzEebSGJIKr
p616jVZuWMCmOw5a/CPsn5khXC7Q9ydu2hEHN5zHmoxDz+5i0X0MaQNioxbFHvekJFH5UgWPF0IP
XsgS5oerb0PFf2caHzHwPE5V5ehK7ljDIC7ZiM/sNlMjkrzpXipexiizoiF+I88e7tr6UErdUzOE
JJ0geJJaZDxBd3cn6UZfy052mJB/qtEkl+Df3DhbxpGNKSYrdw4jAbScIup9u5kqe6DnUlylkVmU
P5aWXYcI9hWUX6HLrP+2oBW6F0/T02b2rAb/rfhEdwuLiVLYP/Ri8QfpUURtiav3LhMP5Snqtvtz
5iI9jCebOhPIf7Jr86tm467k/8MZnaVSYCigh260d2U0Rw8IFcfuPMFb+xBj3A+BoyhUTzH8i5/u
ZHW51z/Lbaj4ZrpOakbjt6L/DqW1odPqf9rjQr8PfeLg+Osn8Hkrc/tYGgOTTa24A+4449yX+tdo
TP8A5aMMsA35+c3AkOrcqIreQ+l+BNxDyRalClAD3PGqhpHI6XvgvQEoJFZH953ftmMa6Prrp0uh
ev0IxfmInGShBnsqsoUSVmrxTYL3Qq2/gitVlTJ5gGE+j/Ms52L90JQcLMDAtsQIIUoSMnq/yPwx
eD9V/qgq1wU7QAQ22XMVV+aK0GF4tN7iVnhl34lKvOCOqO6tYyluiapC0yM6f71eqKZ6MXXRnFvw
fucoap/EXrPpDb1l8Z/ONkzDawd8fml01o166Rkx8ZY2I9twq8NvQD7IEDMRHwXIH05AjdkjcIhl
ei2gmLzEXua0BNaKaVrHhDP780YfyyklHAV+NRKBTDD8JBHf9848SHt7XCB24Z4QYK/sXZgLXrH4
w2mbxJHVLLH9PH4xfktSq4V2c7LkXhS180QWSk7TkVPmf62oqCX1rHK8JkYo+7dT/XMlZWVNHPz1
2unarb3GQno80lmqLD/Ay1L7f/nuhEY88hkUVtHceRQ2V+X3SaRjJ2Dix5azyDuXy5ZJQJejTlfd
+loGSIZ2Z7sr25BIwIcgwkeVt/kQ5QqVok3OPBWhGDW/tTtnwiBSmjWIoryMVPyebWMSQOKQlYQN
NfAxQFhDnGX2QqiOcq/7zpbqOIx5bq3GElkEPL8QJy+5jBVkV0vPSnpRklSY83jdoy93WPgsLQRe
r3eC1eh8azTqwEpU1yA1xJXywKrzrhMhWc5gXJuZMcy9n+Q1NxrF1yLIrRhnmUwhD0+YMU3xlF/4
k42rc7jVynsSiqdmbc+T3lgpyeUvN9hun7vsvL7wLim8KYVUU9TQ84OHHHDpYtYXxAucQoSBcMPW
XeFnzpbh1qVKMPZcvXAGFJrgDqvhvszZqelhGc7so+YkEMLCJq4nFo5Qxque3CIZoA294rA34QNS
oUWsHU5EsmGJEr5vCxBkh9D0AZ88AvE+PDVNxDR3bvXdURuhw4iRwQBg5F3XtDcNV798wHfP7qkT
9IPOC+vxtuO6GdeJBCnFQAPHKCqZlvAvKut8Bwdzz9x7MFR9cjmxD5rMNmk3nShj9frxZ4N79dpu
uejm1Pr+B0KlFNT8cB1MgRNmszA2egA7IOQprgbH5TQnaaCdyP+0fsNcQN9i1N/9a1OmbGBn59rK
2yu02eikITeemxujLJIZuV1OXLffzIbnfeMYQWGERFO1E8yogDDALIghqbq5QdgFmgL1alEth4qn
dAR0EbpDioxBXRn96GaYCXTuajNLXbNYJ5PT+MnxKI5UwPJciFHV9Cq9WPOuHhHdun+WvvgTAb/b
dvccD3fp3c0QgLPilCgGko4CTXfxOSHFlEhxKxRZQezRbLPZB1ctJT+znF8MGCvJ/Ne/dT7Q0B93
hKS2uaoqK6k6GWD8kTfeppwfsyTS9CZ+xZ8u4ZbS2MF7bhg/kQg8iUBYK5Np8wX6Qt+iNOQkqChU
ILYDJs+VBA2uArhg8Q3irIO/rzzesypRc5ZpdzP6SxZAhHHxK8c7g981yrd5tFGR3jelXPAmeRK1
frcWod5Zc+l/zcQwBku/fIXgaoDWmktsQYRUklvXYKXXY2LE6Sc84hnBC3tM8Zv6yulXtScgtonU
N/W0Ye2nH+rzrK71z/WWJFoTNIwsrJloaISdeUFAN4S6gxxoTRCIVLka9eZe2CrT33F/033jkZ1/
xR9lJv/NrFuou9J2ZcMKgbGurdBp305VwO5KnaGOOsYx7mvyLurTRy1ttC8/eiVUYSRcgEWYuGvM
wH1JX8kC3WOGbCboqHmx1MLFDTCKeMJnaDq1UaX91mDbYxNpbfVV5pcxBfe8HeXAo2IvzA80HGLi
eMKDZ81d4hqfoAWV1jn3rpNYmxsCTpAd6hJxH+An+vuMhXWRkhEWg9uFCW1KM1CGYrAD8F9N3zVu
Z3vK7flFXcEH2K2vr1qjxCqCybFUJ8NvpyYYwzOG9I0EFAVJ0s/JVcZZAjDd/m0EkJoES95qsEso
oygM4efjbIQum5Xr8RUX3WHIxkU09dcvPTc83fq7V7hzFIAJPdwAdXqRChJ3/hj25vOJlDE1t5SV
bmL9+DSMJ331OsQ9SSG/y9jF1ufVOOvlHgauitPcOnQfkSLDUF+D8fTPT41zXKptaR7gai2VrfZs
VWBPknaawk7ePIG+nxiHxuycj61CIv1oZsOl0tVnZOjHn4tx1rQY3MMQepba3+bzm+CEDwrkBpsk
DH/1sPElSK5ntHe0IWo3e01YlOTXpxmVyRzu4qx3vkzdzthCeI07En7Kows/SGd6/xqQ2kj3iLRm
kFbIqVIR+0TW4ibr5EjoU5zzMYhmFfzKZT/OWYLhhdRYmToxSoG6p++SK6oAmR0UO4pm2NrcBk1R
syI46cmD5QqjBAYfPx0N86IVuVLukP3bzQGtqBnvDa2KXYSuidq7fDRgP+hjbvES6ji+MaFc0Kj2
nTI8pHSH/L4cZ6iZD54ogqTcDH7v6KpUQHq/mfMOYoofZ1G/4t/incJUAbpiKbSqrI0vkjfglKpx
vLyuTZlsqDJbuQUGdob559DCnR3IPoROaJ0X2upIywLkrnLGi8E7GfHe5vkfx8L941pTWHS/S3Ck
UmPPnoikzbKxFjfUjLLFtpLilmzHVvQbtecQ/+fBB6iB2d7pVAoMpvDsf55wpXjnFV3jlg20u99y
NjLK+cq6FUtMKCqdhJqHR2rJqFdpUsasJn0v2qrQVRBFgCv7jPA5cqbsFZikS7OAdbMyPQTHXOzO
URdK8GxzOIWXjKUNqNd6QdM9YNFSJxRJJ7+u8qaa8ShmesK9tlsA9DuIQa6s5UfsgufI17ALu/Sp
wxsAPQ4QW6lmBsM4ttVnEIvI/3D5XyB7H6AQtuYrC8K9/1tNFkoRXwmczOAzbZIAeca0iQdFQlaw
kwfn/inIt1/+Z3gyK81f1n/Tj6vprd+txAr0AZhxD42FBr9rOETXUrxby8CHf2AivpWKxUYGyhdB
kxC2Lh9irqJVLqerBz/njGpvR+gFgZCnzlsO3mE/4CFjzzIB/q1EHl1D1G07b1gYpU9300k91OvG
Kj0hzaJG/9ebFBSai8AxVAv7GfKqzAbWjqs48Exhl2Y3sF9/WdkItPzZz6iU+bhnXBkijp1RzT5q
xb3apAH84gP1pmEMjOAJH8a3LL9Sb1zM0tfvLhrrQkN/WATPn08wwVxry/XkU7sAaXCUfuverO8n
YRa4SrvsxhjWhCY6VvyuB0CcuHQOzADqD6zx0w4PEFSJTHj5MQVEPzLBObkt+le3THgh2NpTlCIv
2opxYxSbNQcF3lm0mmtTwBJCLcKxX52sY8UcZa1dMcGdJsmVSN/D8NfPj0s705y8zPhYftSjxfGX
MWsxWDqkkWr/J//UQFej9rjRQAKgdpdHTag0QuGUsbtPvYde/PAWBZlaepaj+JhEuF42n0uFs7+J
Gb7+2qPPLHyu0MzKRiGNn5YHQVVemT2uKJXYf1r9bmQOGWUhBnZQKpeLpmk8JAXvZFEiPFnZExbl
paurjMqs1s8RAqxg8qEvjmrjbKBFshWZ9ACbBH3tZVbb31zw265+opB0tj32VX6IGqndWWoXyEtk
aPeQk/0At85hzg0wxYz3QWsvA54ruCuW+0btL5Ea0zQOGo2rb+W1KRmVBHgvQmonfuO9h+xub3TP
OEKqoScRIputuszpYk6FHxb+aRndG0815RL50u0bG6LBip6bCatmGHtMPnKHMowqThcOcnGbrU5a
Pnr3wDtIPQkAc78hFPJ6c0DPkLhJxzzkmqEJjw8HNHc4ARHFi+r8AM6F9P6/7qVpSoxdOhknLVHc
/510lb6y2vqfs/MYH2TNdrFm20DbVtmPwpqfqKvtxTEYASPkkcpaYAIBWEud+WJXunlmznVkrpmr
Bjn2xmh2APeYTvJg3OgWRkNHgf7/r2isPJc3oQn8fSkgA4wiY9Mlsdkq7pO3tSOI7kT5Gv3aV+kt
LKZxHxBY3hgG00QQ43x54X+7/NnCZTOLMwEw7dX2cotEGoDObK8cu/wm59ZmjRrzs3M75OMU3o5j
9l2UFnXW4FQYEgnvWxaTTYmsGMIjQ+uHilqA7aNNw69Ew91AdX/7JOq4vq8cAkhq5HcWZia+L45u
NoqiFimpmBbemaPln7u7l+L/kgVvnvidM2UGKj7FCpdmCSPLkJ03LyK/ThcDgN8DCio8brxHkZVQ
0oEl6pk1CAMOSbxWeEDLJb3xkN/MRAIs8gGcoXd8MakXddfVXX7kqmfd6qujTXVNylPDLgr7k12U
F3WUT+dpdnU2P2Me1d2BGnXael4BmWY4Cr4BPeWzd3czYbBZFBRwRoDKju8MAJPMJOx5KxfMZ0Aw
4LVu6I+OMSonKGxp6DXzZI2RJPITXD+7mRm63j8X2vCYVOPfJ3BplMeGNkF/e1FKQBxSR6YPerlL
yop2ge9qKdUpL8UbNrEOANJc2Ma9XL4sTqNiT8yxwvd7pJE6udzlLZ9OnkFh7V1ysmnlryE+JmE4
ntTVcubt4egzizyfiPPazeD/hoTNmG437Hr847h3b9CyEDDsnQxe6rhQcPPC3lJz6B5vNZvXBL8q
QU98KKL8fzwUYlDc/xfnOyHvA2uJrDif0DB/LWpwcU0fAtjcW20634YtMirka24kRkTIKDRiOZSF
/ml6vBG1XFZnsA9isobGEZfj/IC5rwvXrrL2YFT/JcusmbWbzBWZ7sUgP9HIsA+5fum8hVqeoOkE
r75bvgJMWo/z0M8lG9JaX4GTiT82hzPjhLtiMnL6TcPSGyRY04077LKJJzGAZ5KM3YDmMZP625fH
krHE1x7IRybPNKADvNAitOr+nOlefwqABI4RK/W3bmd0ArD3Mk1nGG4fZftWRTYTc4KkZDa02vSr
qnkX7KpC/Jg1kMAQDYGAhofsd6tf2rIcUv3EuNAiy/jKV1KqRlI5/UuxTO130ND1gt02VvMTxGRi
QahN9gPQo4Nx9S2U3fkxm+/W/ttidTv/EApXIZ1efKtLkZgrAmrYF/PBA/6y9mJuLLHMkUhaiGlm
Z2hJfuppPadV1dK7yVjBXPXyGxsb4zRdJ7AdiRBfFzdpFuu6EEi8u/N7ip3UUGuUp6Sa+7oUgs+A
Xy2clPHgWFkP/C+P5VeLMbgxOqRT0YbNQ0vEz/InMdcvC3nlhQutl8MLUvTaZJbWF35qKP1R4fq5
J1mPp8tbt55CMukrkPioaFTy+70qjN4juTEJaNPeHJ1RvqrcCpFHdWUiG0HeDqpn/Efu64dlz2eD
o9dmkOSviMOuIrYxYDCtT55p3FgV7Prg24h7d0Wy/8noya87aEJbQGcS1+o/m70+dNQ2I6gjq/XM
dGWX/ehhraAOe70rFjzEFSGG7RCxDIDg1gmnFMtxYrFjUgLiBF4UEbYDAryGav01mNkhA7JxDE6V
S2d6dVQH0exv3QX+wylW+ulU2CJvSwUAid24+zRlDBA2wke1Ob8+8uBgAIOLAxgPqW1xGTCqm/sV
JpgN13UCGCsIeO3n9466eUCbWD9F6lJissjnygJFBqc/WzbAUJmjIildC+RlK2wzQxZFPZ7qISx9
Z8Njmkb842vWziNMxk8i5wfIFgO3YrwCmZ5K7EAQIy/+h686vPaokyDAbQZQXVLqclClOxk+/Hpf
bcBwNXIn+1+YoBHDXAVU7b6Nw5Z6O+RcWZg8vbq/maamarFszug7Q/MAc7GI8DGHqESEU0g5+jub
VWviWM6dBh2pSWPImuv8mkr59JWtQnJInGDQdULno2TCfZmZm/DGVnR/R9BAfAVQ3LpbKUazr0wD
oryysiNwm04MgHQMOQU8AKOySV/H3O4ydgNE36JpwsliDmoPNU8PX9JAaj9CsBaPYFfniDs4CJj4
mocmd3WH+gtxDHWWk/nxDcwYTWg9xeDDzkAn4WUToYU4j5v9iql8iioEG9axYcqwCJE/FLdZ+sH2
e+mDHWz3QrddGUdu/15wzDwK+3YAmTfMP7ga4DITjZL71VERntnnP6OB5Ega9PDobnE2R34BcDvz
e1yc/BsWXevJLA1RoErEEY78GDucm+rIhe0ftpGAppvsAJQLghUzrwRoXi7wWQV618q4lnU8bpJ4
wHLSYIP+aBDepdKMu+fcFPIr8RhOywOhzZTVqiGzAcTmJuVpg6h6iDqo+6Ryox6U7yOscuxlIhYV
9HzFSapTfW8y1qea8ouq1P5JdlTUvQ3N4Xkiw7x6R0uZikJ7rC0R7dTQs5ScOOAF2dwHm3TGb6+5
4jO1vSEuWflqNITln0gyANvB+KUAbmVkJE6+MhKECDf79r/Frj36G2NATIXnG6oRllIWXizDWjwx
doWU2IgzCdd1PCCA7BksGg4gxmk7V+GPk6A5EIR+ub68Y/OFlax5gjptomGLwEMasBk+CH4w06e4
SFFdiGLEhx30pFkH3+61YsCvkgax5W+yPsvBwdZawtrzhq7vh5C2scHGFqOxyalU+EaxgIItjJcj
IoAz6m8sCXGu8a1+HJRFL5o0mCmN78ZWYxdGZv3fhh1lRLm+rLofUJVdw49VynVATIou5eFx+GNf
v89r81eFS1JT9RPcWPY/uHAFHczMPIBlLW+Ps3yU8GoFNTJsXj25ZdQ0vln5pZ4lpLQiaknbcHgJ
Zb8GfL6Ey45wKLsl6GI95oaV6IfGqRv0H7vR7MWxYNd+g6wThk+qO+lu36PtPBq8QSmRrsab7wsg
Aqi5g+zcQZTqxA6CoY10fcocGN066uAB3BwLPCP02CmF0Pi3WKyUY1m316fbbJIUyFMakW2bKYVE
dxe6R0TgzuNroIFQ09QniHfg58HZspRMXclPgv5mgIFTB0PY8VSdY7AfW5zS/V8Gnp+CnE768wvt
T6bXDITxM4YDuFj42ru54HAJvT+PzX36OLuUem4Lt9019ZQwum3MuRQX65ZEAXHfb5VDKW2loFHR
y8psps70hsf0OTrysifH4PW5Ni4Ou3usL82nPEvgN2sInuDSaJ3c+dxKgVOxhlUlVUgSRXueTLGx
MQwnu9JEfiOIev9PPU06cYWB08rWDpT8WYup8BRSlIkWWBrTHIgtoiLG55h4UGKJqKyV4aeAFxvb
NKRYIcFLP4qBkElblavuWbBFFJd0+2XP867Y8/oThMqWZDat5uYkoponbAlK6kxLGELuNoq/e02p
NCM5inRSpKF5UhoaMJMQbOQsSObBAP5HYRMall0Nv2MhKR6I0RzK6YgKAI8G0wtbkvuMaJ2lE5DD
BWMQ+xGzVorv6LsD/flznHzlFOq3Nk/ZItEbCsR9qz3ta8j99yhzhtvP0sqIXXLuwahtx/t5zA75
hxWqqvMV85itlb7OwxVLHgHd5wXjiv2aF0bfTGWW+O0g1+v2XzW2cGYFQbY72ctPq3PIL+H/FxCg
r1r+wZPu8Xqe3TbGhNJyEjMc1G0hRLUY44heu53srLIpQPMbybhhUBqLcRYPOOtalmsjDtzsC9Qj
2YCGO0OAdvooxyjaoAWpwbZ+7ATwDvH0G45+gw1b0rujamVfTdTIQglRiCOYk+7rRZt4fg5x60km
wbJTD2X4cK4zG8lSngKtfCpQErUM895Xd3OldRpsoayhUQkUY0eVFqyuP3gAbMP6jcjke13qzn0Z
ZosZlKnG3cA3rKC+PmdjjKc0gRIaIbQDD0o2vPqmsQ1IjY9K2L9zBLYsZ1+QnpopDHZAXfbYi2Dy
WW+ZhI+e15zK4EHZYnx7ekJLK8/YRmmLgLZA2NxxOcE9/uETuujVNw1GWgTPf2Z39do4FVblIVTb
zN7cKx/XTWTR49ftQIJEqOXP2LOyCE/j2mt2R8+/NrQLDgwlgasnB5+EQl00y+T1dEmZ6hDAJ+BY
aWoJcRZ+nsQD2vCfNRiTEu2xp/yLLPh8z6TvhnwHxgEr4mAyUc1A6DlISAQX6i8mYO3ANawR6Lzz
YXJF0Ts6bUeaaymp3g4AaG/+Mhy5AaiSUKw1EhYdpVVcJA8xzEDeFVl+GVwnnm78MSpZ+C+7aMUr
NjfV79x29Gh/CiI/L/UGsx7/qvNnk72McDApjq9xY1pBqw41ZIvGh/yXuwxEUk4uw3yHVOPZQbUW
ViEHlg90xS9hQfCk+vVJQ7USCf/aojr/gwc4SitiKzsEzBNxXuh2hX0byR+eMYL06nQ64BMULkoT
nqVDP9WqvWIGQMo2vVh04EYSHtjDOOpL1hsxiIG5DOVoyChDpPtd5z3qbBvRUs4W6DPMAjU/q/E0
3GVnBMDfgcZ6eeynSEiWmNi2jUvymvXyCmGAYPjCpfHoSd0NfMHlg5NACAZBXBNxMI1kT+1g4m3j
DtsnPpEZRmnNON/wIAVPM9/QMI3e8SxIREYqsxyEEW+KF7/u7kW5wY72CKFWvfBAnax27oXWs/pk
CxSKcFoJNX0IMCiyf2gWDn30rrBAorHTsIkD5ag2hTZ2LJ/4Slx6IbRDh/Cn6zxZR3p0RFjeaRkE
IrL3GB3iskJ4GW0YcoKYYIuOY3KrGELugJj+rG1kEwVsqk5HZCDiXeleKdOl4aU1b2HY7ppnO1g3
+LLntOGOTeHRTrr9C0INzAPuPuFRWiEeHBTF2JeHOzH2D4IVJthuzR/5evDJIOOpEEctDWcGhX91
C0NwCNqBBSNgJRrg+URiKd85sD0VJ7mv4r9PVFMHYoqnLtWXq8aNnsgEaLlEhsdFHFk/Qq9k7ggF
SzOiRRJBRrSA/4wlhb+GvWNJOJW5zfKhgphxgI/VrsFPU/7QbMxuCHUKJCJcWiaPKVAcCnnYKwFJ
ZyZaeHqBUmvwJq0SMOOoh3KT5L7SZj5Oz6Nzk1DwLffDarQD/AqF1idGgZxBdwTgjeTSMxFL7522
4oxdaG1ylp9DttvOIxNJQtTXkAgPiN8EHzvX75nRC4Qeu4U1L2HM5lgRYaGCdwAL6AK1y3o/fyEz
HFhf/dhN2iDlSuH+1T5TcmjqPAn2A3IswLkmud+ARkUW+BQSKrHYQ67kr6hi8HAe/9pKaJh9U3Qf
scuMEBv9s4ajnof1mc+xc2k01h4mV9BIRR6XkR5FMfWPHf2Yzw7Um4VTHT4uLmoF5n6aTUnuZIhK
VI120bujdOEWQqETpW7JMF/ys+IEBWiyf2BTh7O6UXSiVOCcY2aGscESkOM1Vs84goIQuF90kVhx
rDSVl0b5HLbq3v9iwmPVi94EhGuiligTNECMyS55V6jHkpb5QCr+zSFRx7wFm+vT7ax1NmMOeExB
e+HVjCCfk45CSX6OtNUxn0ErDUwHjrJAjBr55+3QX4o4C/aiqjcJlvYbAXyKl83xNCK6dfF1yjkj
stzmoiTGlaRDJ0+DUYayXnHBJelafSdwPD9/sFVBiWHS7MzgSMMlCq56pMWSr8EVvqPcybJdHwUT
yJcqW1dpo2sBxBq0oNleE/I9jrXmJ+eyN3TwkWePQDeOiGh9ebi9z/bPx/Ib3z5wRnMy2aoKYpkr
7nCJobCVmCHyL8X0ZmNh3QomWUwhd/0YqkWQDHgKZnD033NvjWRCy9SUXvBR/mAzQO9weuzExE5L
g1yMz6bk/Zs9DMhvM0EiHezUHpJiuqP8POJGQ2AZ2SUL4hVttu4ivNyL3G4S6K+3+VRkO0lfCD8M
CWBvMsLsfeVlyjFHVcKWWuIVBMN6co6yP6ysQlgBLAi9qtOKRpJ/QnqrcUr3IeRHWTMvIDxGCb6w
hbUDoMeS5uaM/1o9NKDxbK3u+GwpdB7gN0qUr3QgGIkFK3qv8UcO0kwdksSwUcNeziclLhXFq/x8
EChgbWaKQYr+rcWRKxdOPKWY6N9UpOtqPvs5z2DXRGMtBXOHx3VcDFrMw0CtIIIardU9+d2IQaCW
JR4zXzPTRqvoDe9EPR6x9amg0/qvrm0m3zKBp7Mb5F4EFhtsrsLQHgXgReEWsbEP6Kdt4BV0CZ4Q
lmDKMI3QBKaNtv1zOEhVv3YURBCRIGzMlYpq2GZe6EW2eFXrEjttPHpJuG7k7WXSaYUEqAdQQwR5
frgXW8ozYqOSRKib5ke2vxL3MuY/Hb6GIjXwsNszEuN1eVpyThkBYjloB1G+MIS9/lxX8nM41UAJ
LyVD01dR92rkMee0CIZIueW8DD99nV8/4Needn94OgNJQ13pNDEAyXla+7qKbzY0FqJ/feiNSLqj
GbzUQcya33Ydmw5yGPpemubFeTw/BHTTA6Rj37P0EZhlKJtKjk3WUETGdccO7yKsjdZR26mbyAdN
S9aowU8xZ6HYXjL3HB4l2wmOI5knAe8nvwT2VBdOo8MJ1g0U2x74iljqwzYcYMcAz1gtvGD7KPJA
cs3IGeOJYi6/BeGd1pRRM9OjEjlbzWXXgd3M0T7jQXEFIgJvFf29uQtsyDaZuOt4rp1X0eJNiQEf
KfVQA8unW3iJWDz5Qp3vA9w1wHu/wOxs1erY9VjwLZexbMycohgbxjxopA6oykcNNY+NPqwers1/
EKHF0jSXW1EcaSgrOudZO+Ai9wsrKxRXyGA7So0TDwNT+cu2LzSSqGlvAw3Z1PIndn+9I0knvWYq
mQF53jNwU4QOSV0+Qu5253HqUKSetjo9/ksGBccX2rlg3R9gOVMvAniPD+cANo8nwBPixydJd0dp
qS6qcAUeIGFwj0PXkqMs/hH1+A19bZA4zGSFJqfBAIFVJ13d/ZSd5MRj+Jap1o+AvHnh3RhtVntc
IhK/xLmsTeQmDJW1VtW+bageijMGH/QTbleimYt4USn0cnwb4QKuoXsP1mmfobaY+W5vXk5Ijf6t
i97Oger3k0dbaIPEaEtCFM3L11LUngqP3fpCCyyIBD4DQDmXEslq6TkhcHa5HXninvPjJRwqEVG9
hPXNUxYsccjaWXbfVawo0fSu/XkhqTe1pMT0w0ueXMoTZ4LC6bOwyYp2KMYwD4SYi0DCJ7d11tYm
cuAyWX58yKPxHsulRJF5jwXPC4HVB5bdIpHte5AM9WFVPv4BYD0SVmqQ8gPLwSVb/R6dVQU9qvPt
gpVMnil/KpVSOGwW6fXtS/i/Mwomf64NEh9w0urvHnN3vOWUst8QVsqxFBoeWsvjZkXElmYoXZgJ
E6cz4upBLEYcVzOziHkMfAOwJfm4Sg4lsmclAnMRUVHjno15F47T9Bj0S400i/hb4i7bG6KtrvtI
+rtqSGRMoAXHWMriVY5BlyKc+Zp4anDr3WYBkalXEB03Zgd11pYSkeserHpP5ogREkgjrD0cQR8x
OMY5niVbhivXujwq6Fc9OYFdRDFdQEoHFbPchlZORlk+zdnUwMe+dCPJ977brVOl2h8VbE1Or/Gy
gv4fStQDdYMIp+SSW0tZz3qXFWbgn2Hf02pmiLbl7c9JqfKYrngHoYb0q/AxvrXCQ7XpjysQdZF6
dzHlBdvhs9uljwh/4ceugEygJxBzwSIDLQ5iX14Kq2cPiqD106fz1XOsil/nlB+FeRfalFm7OqCD
81cMY9GA5Z0SR8k01MIFek2FJ229lCmZr2aSk6aJLLAYIPjdMsPyXnAX/VM3EH3y9J6z3ZcyGneV
+LAhNmA0HB45nbw/LE79U5KDCI6z6qIla4sQDl8jq8n6fbldaNR18QsvpQPawrNt2Fc7+Ls7ajeQ
/vCq7IvCX2/GGLfhCH1zzw0ONPjNSbkszeTBmCfspaHne9hVxbbYBaseOCA9VKSU/kIvTfQQd/UV
AWjMgoIkxQuoHDDwA3Yg9riSJ34CcHFAyELR88rjI/dMvzPqs+ITNe95MKPA7ZnBoATeL6QmcbYE
nSjaXi0W2VU5HrLCQeidGJxaDZlR06P8mcTZap3MORlvQjeAM7+hDRWg+aUiLYvtoFzISbjg35rM
MYEHV3fLXl/upgGMeHSWO4tFHoIv5HSKktGkHAc6Pb383i3wVyg7KS6D88pfCywUCOUNxdmKb1T1
twHV0cSc/DO3CUtp+MT/udXx4EU1cN1sHqbDTthLf0xLiplbe/XjTPpdsZePWFt+NdocYfNf2oKL
CbOOaX+fZ9CLADrZJfMQEjJmsTZp2fd8wW475FXf9WPL3LEDwN7C51iRxXU8pO0KBvtUV00OoA8n
V1wzUfZWqi/Scj9FEPlOH0NbUj2iW0Pz/6MDhJVv+FLzLqUfdb+XgJMiA5LYuRCSPMPuhwz4jTAc
FEiVF1W7VvserORaeCyucG6v1/2EvAcCmUI0jQyr9AS8dPsdpp3Q6HDPfbrutmfOX1MAwYjrl0Nk
eUZrXy6x30AilL87VV+lwMqBOI7RFIRnzPrxVf6GS1ALKFIe5fYHXv3M9Ull7dx6vV1Ag3D6bN0Z
qKqCRVXIzyt8xSosYM4xegCRMzx7Z70+p52yueXBZAW6h7cewWzLUtXHGg7jK+K1eiAqpY00xy9c
BgjH0hDPYcPLj0r7QlS1X4ZbmTU9SOgdZxi/K5GYaaWLkI68/ZxuwcVAIwpLAH7agyliZACKC+Z4
T8qYypHpGXLyq1uBj5JMtb945lJDJSD80DiYl7umqKWpAPukWmTa3JwTPRyiW7NXYe/95g1ezk9R
xsj9qfd/M5zinV1jvh9Z/YSp/8qcy6HIWnxQef7dExfjq4yqNpiduayy+4iZx/2VivGQBdF5ZOdE
1VfMONOOojGB6fuhn5jmwp9SobHSzfCVN2W6bgVXsSq4V7w0Ma1UJbXm3yx+Kzjw7Yn6YtFt8Udb
5ICr9XVQH8uTFmCv47SOhVcB6FS3oJOMADM4Q8UarWfD0kMwEM/RHzpXRznw9CKtQWqeShIINcef
7z87J71VZpBvfkDCPvZdlfT84RgOEBboObwvw79S5OvKIxCDFMkhpLHpMTNvPBG6XrTFQhzGoHeM
JgIc059hu2/3uPBGKQsY2X6mtvKaJKrXDX1Q95QV5TNOgJvtHIOnpyN043svHWCJ2U7rMje9s9jC
oJKcPlt/TKCvlZn7Bv5mEiWZdlc0zMnUjiYi4QOFTeTAqUd3ndd5UUkCA9XCyrZ3OFaANyWR2x2z
xRzlnx7YUXV+fscMUs1K9QKfHsx28qwBtDvp3zfPN2KUONzmTGlbc1hYXtft9zq514R1j5pJ/eRe
Qpeia+hk1yOvpn+szYN7/BRJMq94slwBzjYFm5x05DmDX9JuXU9s51x/P3MH4XmBuSqFORz71MJw
Eoyp+pG6yHXurGLL1clUTKZyJ5XieFC7rT0UKvxPss63Je8BSS6DlhLD6zi8Xdfe1NPJLBAt8wAj
kQ4HxHz3jL7uYw8rFSB3ZKqQTsbOid+l8Mta0iHt8hL2bQ2K56ALmr2wRexOFJXzIH/iGWHn+h9N
fRTS/E5chAUJD/0lYU2XW1bqXSe1l+81QDrgnTSUUevsf9LJ/p/Q79gt4dAWuYVO6qW3jQ90+kO8
jQfe7/vlJ3+3Z3tH9doI/LMHIz5Sx3ayMYR6UfKXp678t4GRerBF3/lkZrMvofTvuKzAN9TlNrKg
ekD3/2z1tytn3eukSQaAwqmdQi3izlHu74xUMevCKACqpz2/ctd858IleHIhjYNrjdk/Ihpri+JB
XYrLdXJ4hQeye9X5J8X1SqA9iFZfmvQPP7IakQyM4IZWSGVLZWxu3c4UzVY2VXoC0ymvQLNXAfFR
j7uQXiT1Nn+MfILYJvAp/F4m2w8dDeYGsDOTYCMSSVsZSIEOouFUrCaOze7F4yTyKK8PGVoDyzMP
ZyuWUXz6c3iaLXmczaKp/mcYVTucSOuzQ34TftJMkNu9Bv/6jCE6YPruOP2Vp9d3bTtF0vr2ybV5
g+gROQOKSm7xfEPcBqtRlERwQTKmWP/Wiu1AWrU8bx1iGji103H81H6Z5Vz1ctp6dkhcmkuMTTP5
8axzTQVVERL7GRVLTONVBkXyWnFtxPm25dGJFdDBUreW3ndGuouVgIfI7ijZHg8XFfP5VQc4P/HM
2Jl3L71f7YRQjqwesKj8yY3CRbUM2qQ2Lk0MHa86U8lzUBzMBd0LPoGAAQp4wywkWXjC4j2qsH/6
6KHJC8oHZjYcVSRAs/gaZcpOzbXWDl42PdvJZ7P/Vu4fGjsYPv0D21HwEYxc63XEri/V8xzZNFo4
lCWDticYKEeBsy4sJbIN+9N9Axc2ULSCFxbCYE+l/ir0asEshfoe5KNP7HpTsCsb1IUUMBLioi66
pMbKnaKGYiDV2bwpAH4wGJ8IXX7xBbZsGrOR5AkYuPUq+9FYLzv2nNNOrhDhuYX80ulgqdJPNvFY
LYgYZE70gCRBQf0HOn+BlRZVVgEF6G2Sv24xBaNkmC3KDVb0UnlAzGKYkyZWxKqRAyOasjPY61/w
t3ujGGlb8k+7TYl+M4RDi34YYModV9INbbv4IqvFYyIvckCZTklrHpIm1UpTSYx7QgFtC1XrCM/f
KnrxXNbEgJGvfCI7IRoYOGCSwd1yDzhwA3/AmV/u6HtyuSZH6mm5iyVFCWT0SXrrvCz4QTUJqkLc
iOwUKBmfZtHiL5KU9Q1cEnsr3YUwXrVsBPcouOF9zm6klm9eExeSu+awl1G0heVpnF6OJ8gWwk11
o/B73sbNtE5rK8braoNuUlwCOTJzgY8PBNHz8DJnLnP4JQIaWJp5Y/xP6ksKrwtGFi0SNHKDbP+t
dha8HYG2ZpIA0MkTtpmKRWLfD5Im/dBmUYmXed8rdIWGdWgdiHKBoVXVpWMI1hmcLZMdcgQpRhEd
phxljktOdW4xw7XG2u3xQuQxvhn9JVgBz1nsmZc2qaNBC8iwf1LyKWbnPRLOw7DZEhmd+Z9pyj4M
EJBpWoZdqjZ0im5DonlCrJsg3Q600WZ+Sjg782G62KndV9uZKECevX4CpV5ZR4K9Ifp7W2szZgq+
xjBryOr453gobayMj3qg13cWSaebgVLUItRtD8ns6+UmoXoiR9Is+6cfINuSE73avZntOJsbh0xw
xcYKpUIXrurdjXqXrMxk7BTZZuGF/keXvkQSKjLy8EJEpoAIetkfR3uJLfIOA5rmIXBWmFoJnXb8
ZJSlrLGLsFdGw8/po09RyllRwVvBSfglldu6Mf8z4mtrVOloY7G3n/eVg6j+TdX5qOBVfk23krBB
MzsX3wrCIO4tD/eYt5RGa1RoPMnjylJ5y/FEAzpsi5cW/y5EIpwQFzfK9qRY5K0VDT315I64IzBN
0+Zf+zzPMwFwpBVSOmzjYHIBjiysKw9wmyQZXuHZTd97B2Hp5qCIhCEgGVwT0ItGtTFSdAL4e4K7
roiO0Gablu5RfAkVl52wH80e6sDL0OXmSDJShcNEy9yWGL9s2c7acJDfk7Yxh1v9olF9XiRYmyVr
RmN3Y9mVjzXuSuBdp7H3oN+PAoRsyEAp92+3IZVJr5/tOluETnzE883QqLgVEzPkOfYZXKFDyWov
WtL2g/B8ml2/6BQmQTmC+5sHH44aQesyeZpU+SA79EmPlzheV6f576J02YcE7O+blZ4ROG1IMMb5
TN64CUJ1Qu2/9CbuvCxFH9DyIwUpJSYddr77V+rMIrw/rF8Lv6TCprRnnJNKeUFhOHdLn0939RwW
d2MZQyNm4OMIlGRtXJ32x6M6vNSluNd1sahgYrXzfDBiCy4DydQVGSQT/hoPgz0PUFX8OhxCHtq9
tewkBuDnfDxHSEA7oxdZaDYbDFA20P4b+xqCM/kqoO+cMoKUpAGf99cxVG0cuSiZYCc+EWTiBwxF
V8xwR7USVx+GLaGggz1R1Te7eqiGCGzvGodezZbVhcQoq2KtbKTePMpafxJfY/PwcgWlWpfZyKfD
wqPauttnkFqS1to/CYKscuMG89yte44m+4rOI8Ng3zf6htDBTXgmQApdvzpTZApD6RRN2yAAw4dO
GfYKigh+2w22eL4O7OldjYE43T6MFj310jkq3WHFvyiL4faw4kN5+yddw1DNKWl/4lnMZIRB5PxO
HfVTp46qZogomYBJUpNW4JhFi31+80dfNPmqbWQlulG2hLBq0e+wQlrKfv/UNOEV2bT4xPjv1uJ1
TfpN186NpLjPprxWu//KoifaiybHrvBSoAwlw1/K5V0A5s1T+gVXbkuzlMuB6YjnQ3BkQ3SubwRo
qCf3Gh9L2dlrdipkkG8pae3gp6R+g6CO4nSTKQwJGmm9WOUOX3sQw+1FvCdZzzCrb294vVC0t0oL
nLO4ctZPWbBmOcyUntF295U9MZNJh+1f2pVWH2zBI3gmmFl/iubcOnDOuKgNqfIIcx28lVpioGfw
mc4MFNLfobyCENBF0Dg/jZRqyUFDqpL0p6s2W4sgnw3CBinyyqfdME16dnXNXa9rudTLDPMYeki1
YcdDhtUan2w+L52bSkvz0euKnp6LfYy2NGN97vW/cgDnEf32y8rqHyu3wLP7hAVWmQY47el0bcs+
QvaGH3FSP1RW3iiIQZtSba3MX/vuvTj0TswCfUCmoE4p+Hwac0YYEXA2lTJmR6Ymp/ZriysUujBE
4zpRnkkCc7dOB/BRKxNnUJq6q26Oht0A5JTNYvDklSd6CdIfO6kb6aVnJ0YgP95T7Et350HgJvkH
rb6GqNFHH1+TtYvcj3fHTVRhATbiiL7XaQssQffnkPMCjvK2DpGIX+wujudfFA3L/DbaXjyMQE3j
ooIHq0j4dIkKDCTdWTKf2BFOybtNfo93IIniQiWxxWSMgzz51gDVh5y20+ewB7qJtOBPXryqO4JB
arad8vprXkeMA4I/ExBZjbMdM38S1uQGFxliWmJKc/Fq9/iaGR4yM9kYSohTZwWcHCwcqBwg0mv6
pP/MX5/ltFG2NGcLzA6bRg9LptZFntkYfrhdOusv+VVj2N06q3Vj01Y+E6JKLCW3tpMOV17Vqd+k
aJmbE5ZQZ8RIxklQ53l02FRThEzV1UVsc4dGWMW5m5R8Q4vjOfTWcqG8vYmefDh2GQz1CjcbYcT1
jbMcG1I1qB1Pfvbs/l23ecYYvH+5q0SROTo69ohg45LJkSGEIMJNa/GYwpnWj2wpzmN9IRbEb8v9
0NFJ9zUsyYh8ET2w+XLX1F9UQAoIDCFpX/fzNXs5URUCscBTaUpLi7KEgwbU2LylTWBbIEnhdc7l
Bfqytvwj7RHtEjr0L0EcGDNjzi01hcMtnBUo8nfL4wMeV1GXeFdvlucRtTTIcP3XFbBm9T3uHSQr
XtYbEaTwJeL3CnaM7u6K2Cj0EmggbeQMPBQFWgcrm16P4fAFn8cjO+gfRKrvaX9MFFc6rJGgCLNv
IgdYOzlXSYBwEg68s4kHygAOZ2ju6xeLmbyLriHGmAd5lsI0lJ4o4xX+FDSILYd+1EyfWSX+b8Z5
vjGfarfnad7je9y/fBGph+7BYK84zfcLClRm5xMQI6KTv8RbuLItULFlxUZkezvI+h47T9uNk5vj
2p2uyXTGQgOi30c3CqLRuBC3zAJ6rtEiNJ7Wws8oNhT6rPvnxEikbkOypTJWyhJ7UAwN5l/MKi5i
n1apTnKUwWbMaVHPO/NXI8l4t7Zdka1yKJe9IOth49cGaBPQ45MNFXhKc21GcxUVDbijHuNlGdDs
wXxuZcd5a8U9Y8rhG5CS3BYZa+kJuMa8zKXMouZ/vg98IxI6uT7P4jlVfDWi6XqTJNg/QAxXfqfo
0NOUAV+3SJKDrZ2mtFKJEYm+IEqKH9klmeV0HZLgxN2ibio9XsDxtb9/hZWYZwm15Xq6YtV8ArQm
k+f0vD3J6kdUkNxqGlou1gGx7h6Gx3UfjJqQDmboh+Li8ESAeXtIStME4L1WPYEtAU3CtiIb8ZMt
7VNAuvUqOCUWZY2bNP4K8q8WA1ECNx6BbmbDmJycmf2mocnlLKPMmV0iq4InlrD50Jl0KRRBrt3o
wq+YvraO6G5KHv7mH6oYx8sckSd5hxmw6KccGFKof9fsoE8/WK3IKVF+hIHQ/QeDAMAoZvaAUD8e
pu8rHD9BQgM64QaYiUkhLjMVKYzxlANZRyLzWm2/c85BZV3A5TBTdeo5V4VeI9xyZe1no6Nh3tYV
XbabTo+fnOkFbQ5BcooIbb6gMRXxWcz+RWeTCyBh8se9MIaB6yUG/7aAp4XLEAHdLhaf+x4SAFMM
MwK6ZpaC+9Ln4jtpNnjwQE9FMmKcZLkCzrw6Ev7qacGGtY07UQErULlsQ8TO/DdX1wtaMwmwDPcj
EJj2bq29Sr/PmrCpKQZTtJcx99Qbs7IthNADXnLGj5fXM7wcRBsWDZBRXnr5rfw/RMgSOvXzjCUF
4K58VuQ1kqP0ZIBE31xDFFCyYrD/YwVOV+vvA8ZY7tJ4MfYT3jdjjfS46yQn08QXJuaumfJrdsm3
Cp45/IXvre5POmAYfNnGdgsd+rH+h0GoiyP1vk0inz9QVZ34HrM81LgfqcI/q1mx35CcxCcQSncU
UUP61/z+zr86o5g2BHf4hPv2WoYtFgskaGEpHNcmc/RevOv4xjl6v2PmEgjZ3OcF8B7gKYCEsJu1
4fJram6z9ED74SassTB5F3aquJfY7ttYLpvcgGlHc8auMDZByrtMDBsWCK/MQVzYk38b9n6FEEOh
UJXueMe7Wx8ZNlpjDcOJk2TvSGALqi/jYFXt7PzXkIIRqsyNeJtc1Wqnpv/k9HMQYHa51+QySZwL
TLShrjXR9VUqJ3bGoUeaPCJnj1pCHXbO0Xne3Qt9EK7TITnPKx56rZ7nhoiesfAVNpLzrKu+1dNt
2j5s9N376QeLFY+7TlSFgy70uHEcpxDWvFXxAbm02T+7IiGbYyoiPYgZDBTouNZk+/Xk4GZ4t23w
i+ck3/OV5Jc386xoDBnnFqxqS6hwldbwKKTDE4mrmuU8reQrHM0Z6R3nxlUPZ848lOLAwqO+yfeT
xqxx4CyWKSeNmj2a/WAsHbfqZPyCyXkmYlRfnz8PeBWphiJ/dHvDNvOpuDiKlt+nQXn2o/LZr0ar
ovpVufy7+0zjsmzjXRGdSuUGyyW2OZCE4JuSxaci2V6/t37EHyYaQrWn8gKAL1/qEJCOOFB3A3ok
S7a1N+TreDV/GFl9hFpFn1dP1YoBz4wbjkrIEqRCVYNjZ8E8lG75BecUt3hsDrE2NB76V3CptiBe
KYcsOKg8S6wYU2Mc46mlhisACEj4zYV/atkULGI2HLLk2D0+Rja63uFyQoMUKme+EW7VRRHAZrsc
+Vb8Gsw4B3MHl3MhiGbrKtgqHjjRiyurtCJGCp1mJwHY6KKca51q378dFaaJIcRJAEOyrrjUZC8s
OhWVcGSun/GNx4pmQcGLDjU1H77qAPkIe0OIG9SHjeBlygW1mgy2bOyKAHQLvykIlKnoH7lJPuS/
KHBW0cRM5JPLprYKREqQ7I8WiP+/ob/mQLg/S0FvlX0ZgHPc3XKSOBw64OTDH5uaozTXUPIgmcD2
7SuF4ulk3lLh2jAX3YbeFkx/ExavQHPQqdt9uNGypL7Wcw7SW4EUb92O+d47jwLMXaoCHv0vJg+4
QxRcWyRgm67vOl+JpReJWNg5afAYWaUt9QtyMgtbHdthwVvTW5QCuMYpLK9NBmkXbPkesFpkk4bg
eBYMgMRuwEQgq8DmASvhW4WUDWOkc6nZKmoxDfn78BqOndLF1vXoRbRNrAB08iRX6Opja0yXWTtF
HZBIUarCdPi/H6RwRBSVC1lKwZ6HG0FLYV/RhRkYmgTahC+SzOLjVDf31OLG2k550zAQqA6V62Js
uvk8PXjfduErwiQA4MZrXQEKngHywMzETQsLEFYiOjrJC3W+UUUlM9yl/A69idgVd0KT2C5vwE3L
mVclgoMU+ykDTtmAnbiyy0C2iPFlMbkCtSbfbwEuJTWHls9VL1H94xKmW8TqGO0eDLYSfCKB8i4f
PgDAe37VoCduoAJuAWmgF8rrZYqKp184/9EKEaj1zmMT1u0DG3Fp7nWMKbBrx5fS/MRAK8FkLrg8
M1qMaitV1my8FerGDpzk9PvqDFZZK/uQCl5dzgiCOwmGQyFn5VkHrFUZoZV8DO1NS47BSkb8Xrhg
Ab72tcaSG9ZPtSlFsyBv44P58QGwLQqW9ZgWQfud+VTCYc3j/WGSCkb5qWmTMbcgqpKFCOfbvj5n
K16PRLPCtCgKpzrq74+q6VgfUw1E9SXSSKXTzDkunPai+1vCOyaMp+dRIOV3r3HIm1ReAz26+18F
iqs1Keuvd+TFQWA+QmCKunamCkctzxVc2HKVDkk7tMubWYknBMrPP/L8qs5Nu7Sr/oz5pdKmDuWW
Utc3lZMpC4j7wduaW2Zdhn5B0glfNHHrFqK8fylJ2Ae3Bd+s971lC8/Ha/SAX5PriIYoljgdkotE
jzSbw3YRfSQUt96HBbhHEjuysVzTRPGnQXZZN6+3ao+QeBeeryfd3LS9oSzYaJqdLupq3MQltwsT
m7/pyvwftR/71iRkKEK6bikrByWcrycvBzrjOrwu1BPUAQur6iubiQxZqb24R8uyflYu1NXyE0C4
aR6OdHa3jCWpyCkyoWUkbdV0PKi9UpO6G0l/CRm2mwF6UeJiDwCb3xgsAgTuxI53+oKfmq+al1CD
R8l6xQOjweESvtPl9aWQHJlsmZYV4F6Q9x4BRKLv0SsGyj7sDJFxyiwh8a7Ly0kG4bY7QVhUMnJv
yC3myOMKjPDRe9rQ2GOlbPEzI0NwiZ6XbGfx0qdGL42YK8WzqJm0EI1qi5DOJpw3UatFN+TtkdSp
Q36JLU5dsbwp90+XRtz6wDdXybHskkYxfxBkCNOHb5oBnW9JbyhU/rqf3AyjE2TnoNWbVPMMi5Wa
FE4NOp6juoH9JN9rremZHEF/C4R9qQluLVuuEaeVQDTLAEFDsS2R26DLC9HzDZwFVnOzA7MeyKis
+LFQSG3uorwwNg5rCaH/g5cpb3HujlXyByCakEPxhSS2n+ts3scFAF+tDH4SEFMWh9sS5I0QtrcD
Lb+t4vV8M4QCeTFobl1a/zJoQr4BRDHm4YAbOXH6IQ1Sof5uxD7+uvybJ7MCyJaSj5Z2DBwqCnk7
UhpOOcI7GgwSAVLth2JieFuFtgzOV0BQ+288T7IZzuNeEJBxM/7CaZYTESTIfSV/ZNq2ob9OoCwo
Tbz+QNXvkndgb9FAktakx+995W9k6imPY+IKTLWeDrkjvNGun6k4Tin9Acz/Cs43ZF081NS1DkpC
DtTTmg0e3Q6QhDxzBMmgDxW/XDqQBybx9/81vAQJmbPmmGaFIYJKR2s8nuPIYWY58BvMAJ6cmyqt
S0MMQqIMXz1EgOGLo4SsgAI2BoDrYKhNyLXSIh59T++SdDDVhsjXJlkB5+4KM2m3qANMfZLtjrHD
0VdhttjHXU6Aw4+Vqacw0EIff/wZzhIM4C+lTkQ01uSlEaS8ofwJ52x0+DyAwAJFlFPiEL+215xQ
XaK0gClGg3qq1DAdvIPQBJ530risL+vB6usbuYga959wtWEx7bnJRhrk/RMB6bZTCietc60zRUUa
EvXPspJUNGrxk4FlxwCRazC0Jwce+pOt85E34j7HfQw+5lcGmpHBCw2GSLlJJm3+PGQMBi+ZgIeH
tGfMBKjL6ZnuxVUNePKVwnNAAj3GIbPXVVZqI82oRqC1ouusR3hIhZTTjxXN1jHUX9fVua5icOOj
7yQXVStVRu4OuIUG0C2tTOelbmtHrYFtaNMq8TZbSVuExlU17NtQA2C7XHHTobFAj+qznuL2n/u7
Zos3XmKSv47DE6mvLjnjIthEMB7PV3fwoyyeCNo5Sm5azVXhEDq4g+yyFDBnMXYfc3cFU/rVaCCD
xoCMZp0zrzYCy5VP4FH2vEaQrXs+TBHNyB7pVpv68R+xGNqczGE8zwkiDm4jijM8JSBMLbht1Gi8
PTKInICuqMmiCdTzOT+tXODirYyh5dad5lqXK34nI3i8QhdFHtCgWwsdrwbykBbbpwUnVhUmaj+N
prgXkM13SYJsSYu+i/mYXeDQGwCV3GWpGMR9E+fsT5AArwjIJU0myN7cfSqJ2DaJrZcO1pUPWM8E
rNBQsLNiORMJr2JCWt+tQJhnmLVBgA9MmD7Qzdksz9c24fDzWcB5vo49aF1IEBmZOheqtJzqRNYB
gEo/lAGHHqaw8rafuoCvM5X36NzsRMHwsra4MJEqKe54atNj1tjGnmW1jYRe1kSydsQ5gk6GyVn+
Se7aFUC4SD04chBQB3rw0fDBWBSUZQ3CvQ/ZRJksaUR+45QEmae6kGxoUl4uYjoqxCcNXZOEpeVS
Osyo4QSKpSqXAxmt0aagBk2LJSvFP1JyweqGroc5w73/shS+nVJMXSFo6WgBmetv5lpoJ0/Y7cYo
eeZmsl67S/JgLha5U8Q0gnfomrJF1N2f01XqdnAAIK411K78iRimcJabBgMIn+meQoBYxCE0432Q
vjNiCKuO4K/wdp1X0FWic89LdHrx6BUblMMrs1bW6B+oIYtd7cHCqsvwkvGo2lqfOpnOMnsRtLKG
SLSa5G9CAw7lR862Bv6wnELNQQJ9j+kcB/esQBsCsciEHDjFxyOGWljaqjx3TxCanw5GXEHuJtX5
Hpi58FkItY+rPsbw4SfJIGCkCwN+74KSyG0iBRze7LWkgaYXTseWzSbIApLEZEPZrykyj1cbU61m
mh11wwZL6J89FgBqo8EkLvHip7gl/n8YuKQQsw8qOJuzaHSOwa6DOO2/LmLA75eeExl9spb1yEnB
eDGcp3POUWCQ9QRjhQGbz31WeDNDubTBDgNnUhqqmvVA6KutfSzFUe6F206vJng4H4pD7R88aMAq
2nbguAOg5OEwx0p3XDry61RXR6iE3waWsk3SNQfyrbDBFqvAJfMUmt9fE/ofD2fE85E7p5MZR7E+
o/bIXpZzdJDzSpTO9VlV5/joqSB72L2mYBo4wI5JYXhW5ifsOMfaA6MJP4KjHmjklV4VOMP253nv
3IQ+QIbA9PeQMQ/XvTjP3sV4utaVLdsyDPipdpot0fhfElse6v+0wHXpGfBccfyKIaeAPPnuPjUm
Ahv72YuoPV5b51K1+YO0HsWjnZ2XwT6YlDhE3eyrxeVmaY7bRp2Qoyr0Xja1VURXQbS49YZsDgtK
54LuAYStCt1vz2Ctq1zR30VML0Igo/TTCGWFv4CAO26b58l5uh+Fe54qzNNvg9+O6nPcvJj/emx3
wR5QWm/IXESiz2IJuVQUdQcr6hkmoIGnQXH0ghmSYvGzK+odD1RhHDIY6zXB9K9Xlcw5lnIb/iNE
A8OWdUsLiVsmjIXZuRc5aO0WPgMWtJcNGym4CyKDppx2HGSQmg03iABm6b7B0yhJWiykrIies/Ps
OyPQyyAa1sjLwgMxXnpcfzQ5m+sKkvTplB182YGDDqpq4YytNjX2f7c0xXUgPOl9XFrKuCVShoky
b5EufGXEYpev56cvbWZBpbqMjHkZG4ppuzF+0BNOKfqf4vnZx7AO8OlIq/qkaw+9zrd1b7eernYw
WlIYGHGnNIhPRXFkIo/4OQsP0xdNK5CYxb+D2VAwkcN1JWqfbAi2rUeM23yqxVUkwN0Cpz8mBZVA
nWdq1yZbYGycvuG5sE+QqwNdcnqTB8ZVcAcYZuUoohoivELC5rpMFjyn/g4N5/4sRoBw/UJBEkzJ
EtvQTWBrZHco1quoCnBB9e41WM9k5pfCONtU9i3aaH3F5imwBfnuarEcbay6jAzXo0VffdR4kUot
XAsj1v6CuK9S2KmdVF/Tzml2jm+KLn/IqI2jJiJG+ltuF5V5zBFtauk3nreepxGrROuYjq/p7vQE
iKnvArCnddpKJHktsC4yHI/WwKVeqj86+qY3+x34FV/oQxVPg415P3E1egfxLygAjmUEDYQ4ICd4
HFL8iKdBpuAYBsPoNCFNQOHUxIzBhEeDnnt+tVAOvms8FCs4a16gnfmoHo9+rcTuxWe0vpNr2qtN
RevoP8L3l59zhNLjuNbm9BEYElINbLbSU2MJB3ZOV4c9Xf8Hm1w9ziZFTN6sLqBQKNEnwCtlMex1
eQllhFivPAA8idkj9XnHw3okE06QaPFYo7uUSbxlm8+sni2K5nKDabGkRqfUmnY+WJx/yYg13VpY
iUP0iOXV68afPLv7B4xx8ZQkDE0xb6RgvkH5bnfm31IQUxA0C+5zcapHO7H5a/m9VITr7XfmZDJX
jgMR9TOrqNOtJKBTLQJnDP9IYCO9K5c1kvyp4BvG5KP4TQPjsMLEyk3DSaMsHaUxoK/YHAGx0XRt
hFrdNINY54HxnUKsUlzteZIWEr1b9aq3GdK1mknJJ8373p7ZgGKDKv+5DMaIMm0YXCwGJDlErTBX
nEp3cMyE2F93pJP8w7u/AahKE6szC87pQrqZ+Me8PsiZXy6yv+yEQmE0ncfXenxQTWVEYsMi7Gu5
X45HpPM0NQdCeG4yIgzPv5b7BHwxZXa6Kk0euZuNeHImtuSDw0oa9Hzi32EDh412aPuX/4rNMusk
3BLh0S0eGfTkTsM/CD+04/SY4++S+ASkBENZo4S++TqDyqu8AOE1NxxYgqdjQPFsV7LJlFBY6B+t
rv3S7oa7t79y+wKB8GAiC1nIw72d+OCZyS0/IuljmlTa1DH5100Cliq9bsvB/PYJasXCJXlCTH60
WczG2CuovPTon1ki7YglxsMEXII1YVd8d5QQ5Psb283d8n04159Nd+HXc39uEU+z4EP1wM2j0llb
Lrmb2uqMTNK019zCC1FVLDCS5uvCNUqWjpnZJ8DwszHZsIaF5KfwFZ6Gtddad81MW8GIAh/BoKjc
JAFHKbQpUud4iIMkwAKBWXlaIw2yAhSs6EqGZmzmmBLaekQG6FrHjrVJ90yFQ18LfwmP9fWQlDg7
GMUPTQsydjxHnciIkCgajSTsgjQd7XTx2w32mYHT6fWyXcSo38zpJEc8ujCbHfOdkRQbAqTc7s38
oUG1xU4jBlBmEl9KqWk/k9q3VmlHoF8t6GKWSU1hica1FnwXnTeU3o3SVWtYY6EInG01KusHiEky
HrUdSmpP8gRIe50KMlq+riESZ5ctbaNpSiroJJWUSIo8v2mGaYwmIYZVdF05YqTX5HzGUbfhy+qe
NvZq6A9LR/Chn1/3JE/MK0Kw9lScPfxlop9TCA7h8vCcOTz+uM/2dUOYJM9pJR/3xXvQw5wp+k5Z
h0r1f8YhGZJw/adVOanea0XT3XIbTiRgauMWUHlssr5mVKMSEZs4weIS5LK35GX6regCNg03z9/6
U5lDQdF/arF6Dv0L0LDxvD6VhiWrq8iuXd5rSBrHw+Ja3L7MOxe232Oqpv0v+BuF0kSxyfmHwuzC
TzlaS+dPzb5GOx1mi64pLkWl1c7snPqMmtlW95R99m6uupYcUEs8YMpEeKDcOHUv3bf5wd/ApbOR
/etnj+GryE0E6U51djEmkFLK1Z4JfZ2ataR4bPuSvNt7d5T3BPaJwBpOO7r/xUZb5medQxHL4u1l
LdlB6kj4DFNOCMZh6FtUpJJLfoqArDuh5y3CqBRyuX8Q68etQ2RidjFqacMSNMPL9e1NuBSqBOe/
y+IOxhayH3e/4rpgfXRQWeTSaZtZN5sxajf2Fv8JGGqgWuRDDgGwKCs8gw8sF0DcMMFCahhA/LlN
8X4tZqIz7IxVARz1YcLp9hu9s4sO9EYx9wWFz4GFR6i4wp16q2eyQ4ZELlp36jOE9xHIbg7IbgFb
WtvNGy+ZxvrUL8U/i3HRuY8XJw2BOXPDWsJBCT7m8KsPXXGOc+o2fGmw68IQdLSFlX5b05FDIp6F
vj4AYjEA3CB9lfeJEZku9PXsT1du608g4E0CVv+w7ATlbSf2/9YJqbJZlP3K6R7/N5G8O2J6HVwU
5mRbD2gdPqOMq67AVBjGLzdAhcuBT1E92L08Htwh03n3k5hdNcgxlSfydT4ljJTypfITBXAZOeYi
d8YJ+x/SjhSeCX/PYI7hq8qBKaLQ5AgVi5h59HgQGGvqPuL7aPCbP+oiGTFgCF5yPNIKWSgXdLV5
eqdxVBytJE0o+6zxUKkIfFjX5Uas3AF5aLqW25ltuTf95NDZEJd9ptckABx6JOt5BA5KeeY9md91
4snDqGWMoQVZXv/kF+olay62+MvKw4DgqwQz5LZ+u13kpfXgOvXen84smb+xBHMnoa7JQXH1QBN0
4YNUkY30Smgq9bijKLZCZHIEGrmJcKfLGgCltYXHL6rzgsySpaH+u57cOkVh5TB37/tRrZ3SX7KM
lEmaQNU1vV9kQ8n+7+mA1eenHkb03b/NxPbS/rYKrdr1Un00g0e1L45rXxkcZ24z/ULjQ93wvAyY
JbKvrnljo36LjRJI3VenoKA5fzRda46Y1YnEImSrhwzVTh3vZNUUS1UtxuasJTH9j+VjT2sHVNUj
YCeSejHXXtVF7ImumGIRHeB51SijfDSD2Dx3Xr3ED5MDiVsFTskoUrP4A0QI8vCI1z7tN9dkJItP
0tAPo2Ue3QbFBA3952mUkQtnC8AxDNxOIVLAIz9RosIX6GgGrciCxDAwBgH6eB5dBJxy9SbvS0xo
hP1rFsSDDVv3GVkjn9sH58qobsIUJD3Znre9OQ8Mo9o+J1uYvtOwHK3RJ9ESTK6pEt+mcLgBMmZ9
YZOZTTzveqd0QRuv9T2ND0kiJxWC89Q9/guCdOpaliWZkz4T4WJU9skV1VglOuuNNM7k2oBv4yMO
uuDNUBcqPtGB9HsnjYETvIBtItj1KBs00nYvCAVbMoqXf1VUnxD20mNzCt275rLHqlGR24U95F+w
Pcjh0W8A1fgHhQegq0crky1Pur6yRpehm2gHG4HAWdPalA7i3Ewv+k6PJ7FM8Q3gY3sY2I/C3R1H
gb15n+wPfdK1NMyllph6FVPTMejXM4qgKFU1YRF4PTGOzko85l9CG7waYOOW+EiO9kt+rHz4BILg
BjMd45f2RvGwQyxC10FYXfGFQjPuP3zxzS7fhTXb+YMv05pvTZSs0YdFwa0GHphlocLzQDYZrmYP
yT8H0htH7S5CqybNlwDwNCz82T0Q9FxOSqFplGdVPi+dWYKeIvDODYlv3Itqj0LJUnORZbfTyaZY
5dAYYahTKPoCjjgVqtwF4SdushufjjSfDz8gYrfb/u4CQuIHjly74+oDc9dnJEbkboP4DHkgNngI
UCwt0RyLqmL519GtP5p5AT3sCfgO4AY0+3WqMc8s5qW93ceN/wtF0BaBB1QsPt/R399TZoaBtsZ9
5aG4cDt/4tBXfraGD/XwADOGpxlyfkqIQvKOryBz5VuGwh18XH7Rv8bS2k53U3DkvJTXsMrVVgna
kZWX0brbyae5QlUcIoHn/3Otz3cc98UoDUPKRIn9t4xHc97SMVqBs2qIz1/D+5+5FMMGv1uloRsB
Qki+uIxJ1BMAh7v4d5EOm5cgfDZlPb8VRs6pZNS2qZIHBTcxSyiuQVWSp4x8VLz0TX+o3gx4xqev
9maKuNVfGJ8jr8a7fmlYqWQG3IEB5iUyYLG73WHkZEjHUUVMIQiZrTczpnCu0Zp08jCKJHPUhgpR
1DihLUiKcaUtThyi4xv46sFiQMdsdbBrEmCA1aFOenUdQtVjUcvSSXbTuJg4b3n2LVsBHWB6pUQi
twhjIcoJAhtjVHizDAM8oe6E2VjA1o/NDj9EgKpoyQN1p2g71kwlivBJrizkTfS2cBQ+rGiWa+UF
ViYZULYMEbhxgkLfulIsqgrjW5q4oY0uVlpnB/OoGzzrNooEiK+3QWUAItY7Zbb1ge3ZksDK06i1
UvETl5ZjBDS7NnimTQUw9w5JB01CBrKJ9DCQN+kr5tu0hhsu4fN4rqsZcUwy45lHEZiGVBYvP42V
JrSDsBQqYEXwlIUlfbvDaJ3JUnoBPKHDF4xuaM/fjXVTUe5A2shIfdFoBCbhxvZjhncY2D6L8yLQ
Q68zCwhQZ6f2tg1oc78MwEzyF8vjzpcJEo1cv91u1gPznamF0R9Hx0gkO+Zd6FS0VnwbbpoIxIjt
B7qAcpWdgSwH3c4JtMqAN6xBJ2jC3qqryx1rZuWxuZhVNNG8OxpuB2ofv8gWYVhe76xPqGWQEaEW
VG8AdNsUCaddWt7GGyD+xFx3KnyRV6NE5axwkXinC1/3+VhOwCbYXrUJ2W4qDxho2STqPXj0cxyj
EyCAzFbfCvpb0zv3cMP6n3x7jfugxL6oYpd3jKmTlKrDTc9smBl/noLemJMjk2DNBvrRuYlbPR3C
wTNqf2cRsnKpOADLGseK7tWxDueLVCWfoCYTridwwl/AvNqC44SwIDCjBB0O9eF71fOtDXvHp3zQ
qFeSiPMCwJc3OgpgoTNJk+2kozfjP7Wr40/Co/3YnBwBB1JiGU9BqXPx/76lzB2eowPpD68qx75T
0H7EIjnImTzF647CBOlYiwOD62ep90WUnqSxXT+QL6VuHfqWefv4fxnwYQRxLmuuaump5wi7C0Hp
1N/pEF5c4VpfBvq8hV3Bh5/bekKTbuxqqHvthaAqbRBs6ngY6zBaXMCdrc+0bx4OmHL8pUzB3uRQ
XhaUW67kunLG3uKXEBCVN7kT232al2lIKiDitqfPbW0OTJN2K86GOF9PhV0EhuAZYA7o6gncF22h
c2odE8jYuhkyrpXt4zIM52wwYbuH5zRQb5SCvj+SwihdthEpD2ByiJFR16vfCiUNG3PJ8tAOBaVj
8I7bFSTVk6odvkVc1MnAAa72FibEuDXqsbeHs5LaqEKKhgMqTWuOTvAf/lkRXYe4PRRCBvEdLFuK
DCQ75IkckxjB11Nr2T6W6JsF+nUV5QL9VRbM0xQ4ervDXwwOom+Kl+W7S5sWvhXEu/5hG++/lR1L
ou2+qfll0+nLx4S99yC6Soy3FRbU9Lea6P8zYwPmrwQrEREDEKSRZfMPWfdrXGClRs5nsSF5jHNL
PN5/NTPLejGWc6w0EKzSJ7GMqaVsAiHjcYtRpQUq7I5VjMquCSyroYo88DgPXYY1Haas5Qvuk7wu
kbM1/v8st12iJW5VU4r1SRWwD3tTcAXxP+rg2/w6ku6fXho3MDi2gcsFbYv+I3Snffo/SsYXUi5V
M/BPQdYo54/2Xm+R1OiBUG87+JV8H0v6VAKokYG9EbLjSoLqr00VyFqtxSD6P6TR65imbEoKz3x/
YKxgqFee1BT3hEE8l7pFS4NOM9wRkBeGr66jPXuT++JqPWZfaxdYkex5vqHwy8vvj4r8MCd1bAvt
6RLA49XgwzG7361Kzg6x+VJrhBogfaavI00Y45L21wcco5Q+aKupPL7qVZrpijZzLP862p8eYsq7
/3q4jqZ9Z88SUNcD6KN+054WpgkqgfSua9vcqZU09nBQDX0b/5MkOmRprXzK4kija1Hhgfd6Uw2l
Bpe2LbV2Yi07E47z3teVlUnX2+u07r020drg0Ibutft9z2LwF+TOhjWSOU1FcyUZt1IVhPDe+Mwm
k2p2n0dPqquJW5AMuF2krrObDtlCnUpcXYgNwPuCUCbGmbOFq1lberEzHRwHaQ/NokXs7tuEn1r1
y9+6Gmkj4x7dLfeoq2HZS1J1A7lOI5YUNMfajQ4/O3ceinbMJ5m7bYte4yHnzOhVwHkqVAA61YXd
JJteHCY+uCMomzmJVLX29Z/U6DPKLRNzpDYurWK8rTJIkAPUehVjPowL7/Eyq31Yk7t0ifwAJVmI
oL2klv9TNejaCKsvi8pOw7YbmH/L3+7p3OSLHIWff7Qx6DC9aUWcs4+yK3QiaGIzkPYoGrgnIpEL
sSbiyJh8qAeaHvi8aVNJ9rRrGAp+fITh5ZRQXZ9YilR/BUp+yIAi3VoQF1TfAFHrV2iaWuMMNTHy
IzSmPbjjC6SOJ9eslfm224EKwUJJFh3KcIYuxX5Uafrz/FfHNXja1RTcGSXdSBt9OTPaxw2aBgnV
8mI3yJC/CQvp1A9G7GlTrwFeQUsGApsZ8dfbys888qk0GHIJ5hHscTaBm0cVggQT3t0Kp2cUAtIG
R30Njt26YdTYUmI4YtxWHGJUxe67gxpHkCANnGNSEcs1V36Ux+mWtP0bAUcOMUpLf5fylxEjSZP0
VoeGE7pZUjxheDCJhz3uUw9S+oZVKBdkTsM56uHRicLyR5yStkaH+uGofYAXkyMXftdzC+y6ozQ7
y78WgKnNXfYl68Zinr3sloZ5557eMF/hrA+SAOnJe0/+i/p6/tLMTHADZz7GFJQTl8FvRJkUcT+G
nOuF2x1OmdKsqeltPhZOtEcagksnSj/DT4o4mfxVU3Ekeg3nenZhmmiZjouluRgJSp9KOPBHVL5v
WT9HwRLzOYxFhJyy7jqsNAIN5pZ7xohpNWT/+AUIubq7Aa9J+06lndlA1pUB3AK8wGSVjNtnjLzw
qEMVvLXy+x9UzBV30aZFtGoYnoom/98JoekFYw6JjD9ZbKiDSj/HWdq+ylToPjk4ZjTe+B4er7cQ
dUyIh15k8OEdlzkiHAltqxRxb9wNvo3JOhVD6szHM/AbvKieOH9UdUARlMUhOhxRzH4qdDLq5Dix
7RtXp6ZIuVYzNga8RFzHyMXqvBERJpSgEn5CICSB+NuYcrwmMovbugKPpHQ2YZ06x1ZCe27kGb58
BJ+mqTuDQO6Tw9AeDptOIJyOOMX/YdydiNHwqsa1/V5wzV1F6zVNtm7ygCKwkYh1g0XbDy3PQzqB
nfkPkGBZ0BTptjUGGOqI9ZoJo3oVdaZUsAKkX8Ha/9zcdDpJ6fWHFVoFiYxGmuDMpl8NpOaz4PfN
G1cUespPa+CIFk/CAsNgcKx+jfG4l4hg0S3XzCoXhzxTjbhR4dPFmRwNZfCJwx6qH9QS6JrIDInS
c2I9FnHkew1XdIQ3fjnQcP89U45PndjKInBudV5TSqwOL9Xg/vcY/vQMsStg1F7ec/pXjUdtGpOr
myjzpxyOmNL6t6PiKm2qnEUiSoBy+6fjgGtwjqC2dw/EbOmMzgYAMWItqN/kWw/vaRcYA0Jx/Nv3
kPn5vPVa8/N8hzFwd6Jbx/2Ei/mn20z/Cd2aXOZEwNehkNS7e9zlMOhT+FDCqP4T862047WoTMMg
p6puOWL0HHyfgn6jM10Lv+j2MrFvo5fjr7xtW3pBWwr3WXGevthwYtxHxf/zcPS5D9ctzaR8iV2d
gbnRJWQDxSCmc9ZTs0idyIWLphXx4+A/6/aTiKwK1Helqk72oMT47W1xRo+lkZ5aGYytW00jFF3u
/31xFOit5TKoZxCVsjlcdnHLRyNbfZHupH0ipqKjm4wt6Aal2Mk+e39DO6WiTTaLkWCGq9oMShU/
CZUAgGRn1vjU0eOCN3YQdTPjHTTBsbmEma25f4QFlozLtitD18zTcgpbT4Dp/VVXXhDDR0mbaeYo
zpWQ9j0TNNkxJFMTIjmbYH/slSMR5EJ1bKK0ywP9SuVAp7EfCas8P6mhYgsqiPnb/7p4JbWKabBq
h9y/9BDffjBjg90ak4uow5GYyXb4jk6ajg0hSuCNjyKMn2wFvn3z6tbyTO8pQmRenKP/k58kVb7/
xLS/aAszo9vzirjPL+NyjJMOOb5sFEFJJnyZVXpjIJFzNS193LJH/9SXv/VFPbG+M3Y8uqUVFRAw
nXkLpBr8mq1rxqWLpqPpwb9ShWREKQHAjgL2EG0fqKr5iVwcDZ5fcambJ87Q8F71LcvBRK4siZLG
RuCRhltNK6Xlb+7cYGUkWlUUTcgYdGrBz4tWmb9VZi6k4QQLwybs+MNV/mhHTg3s1zJKgCS6RuMB
0+EaS65Uz2CAQWvkxd4n/iVqagh5FGGqna65bSOt9+fTZmsoxKAdEX8bNbiK6TDBgIvpkTqLhmUV
B3Bjad/IL4k9Bb3kowM4eFcU35Ny16xaXlJeK5ejxiQUzPB0xyg8tpKMpVQ2D6ALYJu/XcqJzAP8
2js410Gcjf2ynkj72IdXp3QReLqSbN6s2drhrQCguo4jwQOorGa2+bQ+1O0NeTBXxZ5DxhOKCPE5
S8gjRAXtSF/uBLiJzPpr+RA0g3OCHPBZXiQ/DM/nJtAuvsJ25vrmrGyr8ohoVRUue/2Vvgu5Reyg
ILoo+g1rnCVtXR1qpTMNjQ4Y24LWs9XnwCKVKbub70mhJ3/UGTvzg7VA3inyiUx3v/k413re4JUB
aR95R0ax/bAbxBuu4GDeLVCneeztiYuU2QsBujP7vYCH6cNM3agZy9u8sPGj4bCNtE18ddnp7IFZ
lMalTTmHmTv4KCtYRqIEz+uMmFbzZFmsooyJMCXBnmZcSsIkSaYPPMp9V9B60AmsGMjbq3heAaf4
yEBmmuDiKawXLbCPvqMwt7CLoocmckp26GT+BfN1jXWeIZRClmdN2zLhGSBTK7plfWf1twGfCWs/
M+PMj63hoGY9YeY17rCp8VlK5pPAKqUccXTeO8Z4XicbS8zkz/L60LYtjy+edpmq15bqv5gSx2tn
hhzwW4ldCDuMzLEqb1w+Ir6+LEWzVtsOS5F0AMTYdpp+Hv/2+veE1Ozr/SK0T/BZH3zqD/hw6RAT
qOmmNnMdbd2CPsM6rpT/ZScAbf+EwIMXkliIc0CiEAXeZf0nBN3tGAiKwAoeAsWvhb+vaucnp1ex
NDRlWx7Sr2jriYuykIjVfTNeI2Je9J1Gi8xcg8BmuUfAweMQjZj6pWwOUxeKbOsdYRXSRKVlwDZE
wxC4dpewijDL94yrsQZQmgLonVh1OXCucfFr596ntyinYafBI/v4fC7R9lX6NcjT+ZEQP3utodF4
3y18KARBsvFK0INaCoQgdwTDWPWL6b7j6HH+w8IWue/ynKQCDY0z32D3K2FSHCkIDcmNE+CVngTK
NepetGznzssMmp1wpp+cqtO+SuYePTGyVslk7n9Zp8+IpEcORYfwn2n8PGxFcQyXbncuz9QL8Lcm
HHL9vM7N6N/W1RnNPsQULQ31JFMG1VEyH02JBrHWwygea+Q/YBkGpIY+09J3q2X6nBPVrWk33BFF
BPc2l605vMPx+UkLj9aCUAAhF+xZsNUPNK9RfsZVSOVKsI8fWhGQUGLCmbGQvS6pi3RFSHomNeuG
CR+7dXuLLD//qvAhEOXYIXghg1cQY4LmG/2zrKbQ6cs63euprbO0a6MBPki0hwLp0Rezqr1123zk
QkfYXXA0SSCbjzlX4AdqsNg2zNv+k6//OrHm+a56qmrUYOXSJOIR4OulnEMoJbP2qPwBqGW7l7Hr
Vo8BrG47rQ70kVN9guSZrLY9oLcoaA5dNrEOaSafnmCAS0fAfBrDmJERU6GWfmGbC8s9ORpxpmZQ
Sx9YVF1g/jvfiGfIv8No390oPlJdqOol6tJJP9QCOBMXXCQy7BNfxu8L05trdC+1TWoKA/77kpAa
lMwWsP0znLd4zp9zeiStQeS8l4nxFG62zNqjOczxig+7wX1yYSC/ycUle7BfFjqePkW6NDDfBLrf
u/vyMiqLXiskQGWd0yB6hH7q1TH0nIvE9d7kyaZnAdZvJBjIIcciny6YcyCpyBXi/Tw8fPVn172c
il8sOBGsWyM6AZt1JVQJM1D53/gsov8zDzbUKRWY5Tzfeddn9hQKxIUf4sNilUXTC0rHX6U/C3uk
oBx7zSjZ+Gbd+LGlCI02xyEXk/t2ENqVohCMkJay3626bQkDEX8Ne5EvrWfQL6AmBZpcz/qfsg6E
jlMQx7Ln0AxphuqPTY7fo5j+2wYlcAFyNxS2u6aFrPw9WixH+03Ssj/pYHUYtwp1rot0WXxDhroi
S9NFLrlU87fkb6I/D4xctMCF2JNZrYUUhU/b3yV281Qg9g5feXwCA3wgOpVAuqv9lI7pmhmL+vWi
P98MOLiwo6eoluADG3sGaD8PJN0Wkym1EUKlW3nwvaHrFw2jjnfmoKyGi7xV9/mah0kWZMkMVp7G
6MGAgxFqarl0mN3E8o/O9SzsDxbulW0ZL1ZToK1S19WUEwwAu5jTSiIbdcQTi5EsFuIINVmVf0hq
6Ynqktz64jQy1XVp5pvy6wxTr6Du2jpmtWXy8buKf/GkAIz5zQKuiWfTjSgQX6x8lDrsF2uWU34T
AS69ihouL8+Yyh/48Jc3GWUs8SW7EeViLj0sWJGS1Btsy4VUwJyweYQvc/iRNDKO96twRHWmFMUR
0dMENksXIZb3CDP2P7/V0iWGFsjzRGJ5vQhS4I3A5k/prMBSXwOjBzKdz1yHF/PDu9wa2S1UayME
Kt8QL8S/L7tLGcaZ5ncHjqm+9W1OKW9BJwcOnqnjm6hVmGg/fysdtgc4OB7BoDezH11e+zQw+qnR
7qoYNMcvX8NHHOIKqeM0Zr4ynh2oaHMIeLUQoXPr7bL2B9664oA1/ZH1gKT7KjeiZY9BLs7pEwJ/
0yAB4XrAUS2fwlEBfXU+AtLni8M1R3bAPUV4nlEJ2Q15yI+z1hZxhfVr5wVFTUN2NMscrPuSMveq
VmYh8bhnlx0b9iI7Pj6CivyUVVCPFaAe4z0Ply0Hjb+wL9kxIcm7a6b/mIcvxoQNsyFc0kPVT/Mg
IGVE8DzgGj0+n8hnidPWG7mOwMw4Qz01QwSZzP7FiXfJa9NtfEhHfgvV/e+pZVQXdLYKaAE6XY42
4KuygGLIKKMFr5FR1NBmVscyazZZyUB4xv0Mw1CqX02qqpVeJYQdPmclVOSMUvlTpJF+m8tRt64I
5hgri1+rs5dbrULx8LrJhLkRJHm1WBwqyZ86c3W6bLIKJ2Is14jp7BnL/uoNtp5k2BMztQ7/v2xV
sydRuex+oZtYZOsQ37orAOy8z6HHyizBkj0JsGs1ErBEuKIdqFPCSwOY60v+k8fGsuLB5R6qwCkE
7guSJFfgxnh6bgbu5Y2zG7Rl84Xf60b+b29NxNPZW0owLb9XAwItr7z1iwz+taoHOgcncBiVWopk
9DL7iRpQjMQKKvgX4Y+yh5JipyR5y2qd1Pqv0rznPhM2KOQOa5d7FZveneUTUxQ+fljHUJP0eIAA
6/5T9U1lQGCJZ4Gu7yv9eH6IMqjisJJsWn4a55rg1lsU72zcmHrcD65BpGN+zJV14+DNf5nt+ESu
G0Sk7gufZvarlzm4vrrDyFlZzu3WHU896WAMOcMuzxHtPPzh64wAaWLZHvWRnNCxZycZVP2qFWMs
LaiRRTi9v8uhPnRQJlBmIR9JkUV6lklJACXm10ny33v279vRBm8oN2Ul1/HsQo683LVVsy7dj3mQ
4txkbKen2Jw0TyxBB6mxNencyxfNbHHV91FZACwSAxa82OYp7HTUVgiJ8/YtyMPdXMZ6Kfn+aC/8
mLQjlAZh5r7c/tmfSuZaOVoK3jkUTYeurrEH2R6ujE4Iwks1Z+jkDmMTzc07/rA6srXh79X2+IXU
Gyj3KpT2itDQhN/Z6NQvfeVsskmmMS968FKaXb+kxtD8g4OWEJqYyoWRkmX+hTBcq0jRyc5knLDt
4ZFwPnphuecXhMxNcET7rijGwrt+qUh1IkngIMmCC20rCgmQie/CPv7P4cqRIyg9+lIDT6jjdvta
/e2knGS88EC5VTMdr/V6tvzNXsfa8YfdINR3AzYby1w3EIyAR+/8MicqcQSFMb33bFfvbNEv3dFy
3uymqp8bsSAnKRFes1IzqJmciHW/vVhSddHsfLY0UJCZMYoCerqThkUviYU1oehDH58c1phKpv+C
DXRH/Gyj356PaVbHUTe342VE0VUAPFJvTEAN3rKsz2Jtww95QfSsoY0voEYMpKUXsA/c584Poc95
rGkI5DmrbpQuLQbl3QOHLwxbSWebeCRpQyg0UM4AMpE7XBsmvC+7eIcJY7cdEwc1XKwVL/fGLw3d
mqv0tgPyb1JL4MeBBv0Wtd53vhpAcBMMDxo9yZswbcpUVfcxSNx0SXBW9pnm/4O+e+Ykbi2uc1dc
T0g/p9/ZeCLZCPus4R5bF+Tgz8625vh5Pk+CLDf4QceHlSiiq63yuXUoPUMPaymwVzUzt/0qhhuq
Je9TGtS+8Ozn61q2zcQr/NG8fv9FoxquqmXNPrDWMCFnxVeqs7NVnBSCourE7fdhR1lsuoBSnVne
xQmkvfNGGNPMlp35/0jAux2WzuwG88gGF2XJYsx/AGHQh4tz5wUFje3ZptMNZDqr3QjOq9WYdqG4
QTh71zy2vSHASYFaPdDrPRScEUhVQyCGRS6aUVkuhO+1YD/6Fhtp7Qy95gMM82HhuPMik9nauGvv
RWIbNaJAhpaEZlGD+g0D3QGqCMctpFqrfUm4lSE6waCxAKM5xot3378q5mAB3a0J9ei9rA1l5opN
ErT8sHLQ3HmCLipjDQRU614yZe3kTPpqpJEtvExz4VGTJEfHMaC1jaxiendB8apv917iGVOpV5Yn
DYarCCsjqzlj0kqGYpw9ZZKrE8/aLxHf78fwm2/hZpAgbnSLgcigTQF6H+CDh9D8BAQNEQOB4NP4
LB1zJWBxi+nhdO65jUFOQSzZCR71/wbvvh2wtrrpqy9BHbk4fXtRqUkP2rER8iYOhWXTrzU5xwDm
NijQ/3TE1Mb4+CPcqOLZhsQpdEr8Wp1XbXWJiY5TpT1uXOppYIqAg7c+rCah5FZI93CdSpQBTJvw
+gKcgUqXHvvlhJc75TM0/QdKjblxRYiwevkIGlm1T/WCQ6EN2jKll0Xr9BjHg1XF6D/ots278/Ya
9/iXLVBHbDvkJj1u9epKVckeaMGKJniKSnfm5h1vncb3x1ekDj3Ikg3alnc0KfGQUnzvwPSIYEdU
pm60sxPGc+qx21f4S0BWHJMmAPzw4Z1UaL7WCmjLPdYAqsLqBQZE2Rs489ZFJkVLYyLZeUmB+5ar
eXm/555+8gC7w8VkunTb1QrcgE8UZui22kdQ464AKwknzmttV8mPz3foIJJh+8jP/Uzztx4vl0Tv
F13hU0zvsfvjQRHl5EYmK8qWTRwoym6lhZw4ICW25PQCEWHu3FynrbEXREx0anpBa1osNXLcOo3Y
CtkfDRY9xPNXglzEph9ro+1h7JyOGXZq8mAvQ7n3mA+98tS41NEEkft3s5JmE30DYCGAwsJhm/nO
vpvCkFo9wrpV6vZUt52B0I7kjULIzTbXQ1brf8quWrPtceEYHkGEoNjWS5sXVIxdvIVHGRSf24Wn
oZgewugWhExZIxMYW/uspK5e3GUfcMXav+Q/5GYmOhdfimoQaaFDp+R/DNEHc81HHGxq3z2Zj6gs
elFGhHbF6g2wFnDHCArfo9DYBlbQzV5lb56gUMBgOt0tagtDNCAbc4qBVVq8S9cwEr/8mpBh1mIj
vmc4NUhjVgwfjENP+0+mXKrUfeZMP/JMxBOBiseSiIje2lUifFKkQvX/6oE+xqViIguJtFNYf5SF
gmRfbQe6eIRo0EJ6t3Prg7VQ9DZQAHJk83jM5QcR0Cd1xkvxd1GUAVUvnO3M59nEb9PwkDisZTuK
XZ1XAAnQyFJebnkluVPZ4WOQ9Nilu6sYI7tEaMFwIAKJNeDQ+5y17XAhj28WhBriLkSuLM8P6fqy
vF5xJyVJzX1/wPotF65wtTQvOgXZgKl2tcg+r1jclT/uuqh74Hxv3ckXass0rdQVcNFwyXVToEqt
RouU8rpN6lyVk+CE3mK1WsLtP2HjMNO9Qn5X2rsDehvOcV5+gZ532jzZcyXMuMm2qf0gNF4W+7hf
aurRBAQZi4vstfK9qzOguWmP20XX1X4T/D0Sh4o5JomnFsph4LQBYb22IeHPLDzrybu9cX/xzeNd
BaDOx17/MNCIk8kobxDjvBATgpao/YFyRoZBokfWq4OY4Vtqsgh1zrg3+uvkp0zmJ9A1NhxEy/x+
W+h4sY/TIH4KaridF/qNhq5NYwv4Z+y9G+WaI+5nyYx2BA4uy1q6xvg62xRr7Fm5auI1MZQFopld
zGWWM0zRL+t8qi2zfPZN1XQvqsE3LGG/34TWPJ6pWO4KW5SQ/uVI8Rwz0zXFU0HwcJJHcuRyzWBp
gNVVzzuNDwIFh/0ibpiuGTV6+zwsJx0Yn6NsCTxcLTHj86t/rgvSK+/sVYvEPjq5lCzbdBVkJmsZ
anZRmZIY3IiZC7TaK8eYur7gcYt2fEmgWG3kGTpAdyHz2dFjUnk4Uqikjo4OqYrQSWdBxTGqDQtV
dXe6h/tiGSgAgIFqu59Fv5GC7XKtT5BkCyHHokI/NPJUe5F8jPy8/kjemoDQtNTgbvA5TXuN3hhS
oOHfPCvGWKyxr/pH1FZNEXMq0s7wfl53jjdmQaY1K3hQUX0abpPuBdZv3dRDPLkxUvHu6/TKJIaX
p5l3ZIggdluFTUK+nrfy/hYnPz4MGaBP4ELgtPIhfgGClZlSnHLUFRPz55c3KeygEHh4eN+b6MRE
J1icOJou8C2L8Ict+FsPb75d4OJpNduIW4q/YQcbq80CZ1yjPosywcEHwPezRu9HGBbVN5dWDG6L
l4RitaYddwEB93fbCB750A2lJOYmewlJuZYz1CVB+IaT5AiQWZMta+k0tnWI3m+xdymwxgeaCvpu
RfED39YTvWyowxKxYuXPhtwMFhDBYL3n1w9ZyJc68lcgbHVoMGcHiL8y9AAUZI2YHoKjQHz0PbfX
yLHex6CNeOwpqMAGhWRQqcbjGvU4U/CgzY7NhW7rWKClcTjdre69fgBfjogfZGSAUmhjuJ2MC2UV
PUQ5AEBRbT/qXpPUWkR+Y6X5qP78+l7EyBKGWxPuLN42NuWSmzw4TRAK+AE/4pgzLzCHE0bL2St0
iVXk798DYtpgKKYzxCCaSy9RZSWAlfL8oyc5VN7Dmu6KIkd+qY+21D02izf5AtdfaL/yVs5BI/Sr
gs0cYFGZy2UoiUPJFt0sxzkwQ9fWHrZBusuuBonBlLnLTFx4oLUVSOtPczkpgD8mIwwPJauGFmfo
vvhdQoQLkZxr7C1JYf3zS1u63fr0vSMCSv78LxLLxR09X+mA0u2m/lPU57O2rvz+ofmTKC/NoZ1K
T1pESJTuK/NuCu8bVWBCXsBKkibb8mUarR/G8xkanB7r8drlyQTcJPieB1GkKRTCJcqh4LX2R7r5
vDIWh7jRFwc3j7d3dDXyz4Em5aAIKKUWZdFdLGqliKVoODba3MD/vGhimghdil6zjumdxZYEKqoc
6RF0n0ycmDgRcc1moCHlE0yiJplQLPjuJau/8eIOA1Dg1esFl4R0pjFI5U0qd0jba8q+e6hq3G2Z
HPpmnw7dFBdtTWVwgLoCMKdF1oEsnAli5A0daZZNf3pGU/BhYnn7A8m7G+vNB+EK2XRPOSBTeQxM
RCuWu4kI14a4a1SMf/2C8GsOvA1a1W9hVyf6bojlmDXsaCv2I2p5VkFdbTe3YHm4Iyg8MLsQeKPU
zLTj6+/avYGcHwGPdnCj7oXQWuswtDdyIXhk1dcSeokEx3pWCdtjPUxqAtnUJ4D9J4s2ExCmpKGl
yzTnYM0evJIKwYnF0W/DZuXBiuBazPCUDroq9b/6E78+B+htqjpSzAM3z7tYFOZYSJxIuPZ2TnCe
LmB+mhC2A/VCbSrh1166a6VcdUCzajyvZqjAvR4vxwsoFEuPC7uh7SICtKQ3Lfs46v7JfTLWLoKV
b8GDEABa6fbS+xnJvyzFY2mDHYYTRza/VXBIRbdQL4g4SlxZMYZZhR+JtBVyphGj5qU99EsTyQpN
1/MNePmSMh3yPGw08b7na1GYDFKCl1P6zj6zZGZL4uBcSsDY/zLxDmCbpjSUzpLKjHPC2QJEkIm0
QbZlKWt4lHWPdiqX10rI/rWEuCdkCfDZnN5v6nM7aI3KGN7voZ4q277Yp+kw07XLE8wXXr52SZ63
YOhW7ML1P1ip1jN2Z5qyrhyC8vNdJh97NA84bLiSj4xE3E55WSmXe77BV+TiusAcWXXyDkUJltp+
j9NdAOnHAHQKprNmnxkeFkydcgEHAuePFPQh/n/O7dltIT6l8+vG+nhQZA7HvntsTk4b2dhzIdk/
nC/ceQy+blj8k2U2AXmxmsGKLjV3J74IilrR9YEgHDJQYQNvwTC3QqDQeqx1chipf3DtThostmqe
P/oEXzmBGlyF5Z5X0URw8qZaYq/2HFAtWXoI3+vtFfaX44f6Gy6GsrWZCOjvz1woge3sWyymDhgr
IeKGm3uH0biSOuEtf/Fp1HvD/t1sQkNgJ7XmHIoBxssBi0JZ5d4DOo/FBKG7DK56TLqEvVvgYaE1
ODHuqK3dvrbKB2++JgLAqVUG6FB4hGtX9PNJ34Xf52hmPXe2wkdfYFEd8+jt2DF4nUBWW9E2tz5N
xE5F+CoK7kWjl6oJRVx60Tf9/rqpM/dzFe6pHax/5CsM5ME6cEzY8hvcWgdUvty/h8mnHI+tZPQd
jG0oxU5SmDrpznMi6sHTAScxECFSL4/zOCSlIiYESWhCLXymfqHw4xrM7Wq0YuWxim46zc5cE4ux
zJNkFKRIK5QTpex31llPc7ISgvBBDUJupgpPnaJmWhxE2Bg0Wc7tbMCUxz9P8Za374bp4WBw4UDN
RmZRz/jUaFnWkNqhfB0hUgIHIM1W7Pn9GJISh3RYpIM9wZJUhAy8bs51EpUGkf0eBbwZ/kjBJVJy
w7yPrJ8xFayPIIi4XzCW892IOuGyLtWIoIQhsZvMVqDg1p04sfUrKMk7hexGbwXnY4YKv9F6xNlx
ESkz9o8XoWVRlQNmizg4upq0cQRe5eJA13GFG/kfeMCfecf6SSZvrTyAn2hd6dZYynxsB/mUUMsS
iNHnQelVVRO+Xy3JI2YlfggIfJBtsIPuMCaC0UTkYoSj7L0P4aGgrC2AenSG7WxI/uQUWejGeIXc
wZlnVrIR4Vjj/da9kuYfnodOKhoya8iBo3org+mNvDf8WzWkXZqC7kTFgWmNZ64XVjm9ZHtq/bG6
bfOq4vDDw/VeULQPBzmXXzCkB3DYy8qSXsZCj0rw6dsw9oiE4iUNENs/KKc3YHkjvFLML5kpYCt1
1aJkhkHH+o+Cgjw01y/7vkFY4WevywmG7mHkrDn+9Alt0ZYWKJfQYkl2SQUmPn8Pl5USQSeJ7piY
KGtGx+8XoZtfyU1BUjEMcdhCwx8x/eP+HrkNrb/g2L+Yg7NauHyZ1VBQGquHwS0OGbdtdgSj82NV
d1Gf3MwpMDJ/lT/dHuDg+7VRdiYxGH3+z+MefavFNey0OGlmNtyWfBo9mTMyVSRC8NBVb3+RLhQ2
oVVKCvRFJRqGZcO958afGYR7+s/FM+TzhPm2+sFMhe4Msbyu0tLL7XZuvysbxQikMK9/shUWuZ24
Wwpz6IQRwcuNFWrMoprYKJnrrZppcCzjW2Tv1eoLaj2jbNWEhR9TfR6hSyNsK5fYEwJ0Zao94AA/
ktyM3AREzpjqkvuTMOUu5eHj8a4Jp/yeinmB3EHCJChVU8qa7uPQZTvc3l8s3mdspWOHSE6b7CHC
sGYf3O+0NZjmAKv9loIVcCG3ti9Modk6euBOi8zbDR7KS/rRBs12sDj6wipcAljPWmTs6eWIuoyy
Qo0gVQcNadgxIgF2TwiAKnaQ7lS8INEFXoYVfbHd00stgcofGUBcaFHQBV9NbckEX5FTH7HPcTu/
AQO1Fc09AVG1LC/VXYIe137ARNYZw1FQ6gPFsPCIHcqi4VO59S7xAosVZoDMYjd9b6qnFSlSuBBI
Q7/D3qnxaxyVCXLALUzt1dllhCwpjPLf+aEI6wxLmFgv5PoxxaS0Uvjt1eog7bTBy2sgsmy7m6Zw
o7OsT4Shf+Jo1qLMDjgdGW2LyP6K6x6YhmjkiI/n9kV1DAOHQSENLHb30hSGaD/3SuEc7RZWTczk
qHya5oTwdTAgoVaD6kmdlxzzIKcfokGdhdUN/ASrdnBtqT3CIGHmQ0L/6Tm7hHKnkocb/SpnLxio
RqWN+DrmOhRJMMGpP7FSY01d7iY6hASkwgaRRzefeuS9L5RMslSqiiPk6UtF0bUAUjHLqGNe2vOR
byj17fWnFXkG7MfkVyzecfENluvCtq3JEnba2JeqB4oF5fxF+1LXo2sEL/wHwFnr8+fIk4L6m5Z1
i8UZlI89GEZZsRl2YOzC0s1qe0oePPSZmNbiZJ0Id+9KkZ/Av3cFQANxkEqK4tYkEIp0KYvamPyi
4D9RoPukrf4Y+vLv+3JeFWgOunVHT8S8aepdsNmE1tLgBHUq118aQy5uzE8As/SXVIKcvNhZ05cz
KcNVmPGOQV9xWuRxuJLFQQKlplVZQlTKu2jv3RxSvXAsQ32h6jeTT5TxG46xaNytnbu7d2TPTMd+
zR2N+s17EbUxLrB1HEvxdj1PjIRd1uzb3z6HhFpBvruSvcieRco/jf4wEE1tCUBaSFA7q7gWQm7y
KkrzUxGbEqMhUNFN8FIuQKCF8Ss1JRHfjsPKLz0qVWeT2g1msDCDWqnAo+8pUhIO2KBRr1TAYYYN
rUfDoIqTIpLN3UwPbsMFWtN10grbrKDTmfRV/kPXfArY6UK6I3v/O/6/gsfgtC/2S3zl8r7WHWu6
QYcNHnXhlYkcQD1M5E64sAvOHAuN8UIhQM08WD4azhiRBs0A6DeZvR9A9QPphxl1sK208mKcKUxS
wmjDZNuFqgwAB+ek0uZUPDlL8c+3AQ/L9IWJ7YY/IzrGqhJwv/UAiKWXKBVajNht10T75Dm6a8NA
48NiF65/qSj6tiDwAQ+XotG+0exmQ//qbKGjIE4MymrgBS6BMfnyRTbnYIaO3JBMXbjwYr+338jq
IucfIF7X6Y1mfiAA+ja4I/51By/uy6M3WXk3QDhzhqrGQekqKmuxYV9+l3xag/A37rNPcavwU/hh
5O2gLFr9H0pZsWwAB1CegLTdcQEj8RqCbbhGllb8Xtxqm7v5uTJdcUpSDwYYs1ub1vXAN35S/tpv
BOkwEW0TwvvelRkol4ZgHe+JfDVOLLbkDvW1NsaaBhq+y11K2zpKhw7chQ9bT+i5oZf9f+AiFItQ
eZDuwgacAApsRknSrKvOh1OlFVw68OjaDTqkXEZd2db9oc/r0M4NxU5n6D3pc86p7VSKvBf47W6C
ogiBO1UUnwQWf7ILl9DUweH6emPkIuXD3T9MGIKGeTTAVNWwxPue+otN9Q/l4yyNHFw+bEJOeiCN
nJ1MBFzTN4lEAkTVebKiIiSwX9FRnuhC3Jb0xqTLYdWCGBCj1dvpHycCo5/QvDGbVig6PvlemdgZ
prZbrQkY5OKmHckK1lar/2Kp9Jng6jzzwKIT/3aSi00cEJDXN0+Ns1xJXuOwPrans1KRLsjDEbN4
J9RwoZPnOHcHGDMubioeDgllTZNNALID2sRFfkhhIWYb0aw8QkefFDSNJXiE1tBzNoFx3CtXTYDO
2PrgTe2iR8IGkFXtAG7+03I58m2HEGFqVudfQ9T1sf3Za7kf9/j0nmpOrMJQa32oBRKrcLjLPb2k
U1FcfnnrHk4D/x+hTVoW8MpQA+as1jqfcKSxGSPvYK/gUCAHSxTRPg1rgQLEH15QEN7z6qyIOc5X
658q6eeSabbIgWdQiPrs0TSQ5zVj9VRvMHgRDlkspSYnoMaYioT4+Kaf51PZ7LZhneqHwA1F6mba
SWJgPBfhsOM+H2FDk1vebiAaxwBgWwJVOsRYfba3oIjdPsKf8hKb4TN9g+xizuxxph8Ol7yyahLy
K0kCM48ruaixS9EUqOZTLFLbUiSFwgKFMsPUnnteHnDRbvGeGTerhY2BwHboDpQy7D026rRfdvjd
15dUkK9FdiVClWqsxkr8C3Iyp64sC9GJB1qwUyviROMf3x+qaecqdvRcDeYQzAuweJ/+C89kz5dC
Ey7J5LXh2kgBwU8bW5GIpE2OWFVfUFmKnZcX//uPtkP2wsHdhY7PBUxZGvoitwoE7mPm72rXzpOp
R2Jt6d/0loQmWa7BHbP9tIDXXMIwo4aziXUfp6UVnUwWZUM+WGnDAy0NmDoe00B7k0/lIHbWaMmx
U4l2m9G3ZFXsZPa+pTcjmF5sBL7sunfoEgqNXrvTFKunptj0jHwt3NNZPUmF8BiTg9oZuZ11iBCT
XrXUK2GJ0jm03eJrC0McG6eBkBpkWqOleQAcCnzNjyJzDv9GWXTJRUjtJpXnPgJqbCTHilFAR0zl
JL2WtpaPDia02N6wz+BgwqgxRKkzYe63XvVDATNCRGZnfX90BykHf+cdG8s81mh1qUirX9An9HzJ
M3vRkNDZK5vYEeDWpu2iSYrzhk3cJjUHGsutBscH8YmwvHpMq64sWUWc4YPbNtE2KfnjZvLMGUKh
omWp1A4zgFM/QYyYgJ6Z7Piafqqa4JYNDpok8EfZl7tIUP6ib0pYYlGoWVQ/jEmZ+gUEUwU/IQh6
hzVrmQYNMFObcKQLSSDYXe2uhY2sqHxtqj+P4fsFP+cnYxrcqgAvQHgyFlhIXLvIjmFkbG56P2+G
1+oW/welVhkLHv8+N0Tldoe0L6teGAZuPmzxote5CjgbnXfn9aj+TnFoTGXMhOXn5u75DtZyXFB+
xpT5ivW3K+PQ5Q+PcSMLqQwJKj4nXBnPTeLYcSORiLH9Ws2UuLvpLoqV1aQefb+Oo6E1EhaxR+j3
ZbjXb1dZzBSeEY6wtwe4SQEL9QJIyFGDWqWVkm5LO5QgFcW0adwNzOgZa0OZVkYUt3ZbWPlxloZq
CbTNaxyU5F4KtUje/ZCCaXJ3/j0BER8DFcrMVsqVuuXGp1X9KBjMLoQyFZn3z+WUrmq2sNnhUnsb
OespzGJlcrjq9ABWA5nbfvCJI8sKZAzZdBg3gZ0S05boKWHNnfjhpu63LCzQ+sZblY9GdPmMTRer
Z8J0ke4uvILVlBcJ/WH55yMaYJCj9uXWojkAm/2pDp5y0EU/huoJHt6p5WXY1LtVswzDFJxUcKGz
687zv97V4vTsLPF9ENZuUoAOOGTbDpDAG4T7NOo2m4rWLQUW7ofUuXAgBxWvUieYNz0codQ6dNJr
FdNDSYxfxzg1/E9AvwxqHZqxGtMbrPgjlCysb+Varh2evcV/oIQva7divgOzOVPHIfplB5N30SRl
ZE8Rmp73Qp8Ll/MNTWulVqKtxqcW0dzL0X04J1tRFdVFgNclS7spQ/+rNtT1U6tnY24j/eYmN/DF
BsVnbwEEJiqvAASwW3EppMPQtFPkOVJquM5/XuCiAxU5UGL6SWlwMVrvFIZz/PRUWattBcJ9D4Te
96qIwzx3mCwMbRUl2ahsRysjLZz2TMcnMotDIhz4+d2jrbD2xmPOzEXxv7u8qICieTQm/8u5Ebtc
iuBt8cVC6/gKfvC8x12tuuQluKZEKhZHbFymApjg2z8ru8oOLPFdqlVxPvbMKcDe6i9ri6IjWvJ2
JjpgnGh304N/T//kF8OWQ7RAHKTP/FS3oeYHUFiCqOvo04qhFLzT0AzeykPv7j8oDf9pfeB897x0
ItKWnj//RmXLR77nA/5msNv3Mi2XVW5NtKrtB0ABB47WqUoAdzgm+7UJNJypoALNUw8WReJMGgEd
HymbNsSX01P3Iol6MW8Q7PVpxZwd/mOqOQ+us6XsFdA14mjgbXCpWe5jHV73jIEY15CB+JZCoE1j
wB1nmXA43AMnhxSKtCY0Lq/PDG8CFRK6/ZR18V2grGwsTh+unYynwubMUVEfwLN42PiWdfllApwk
un5vaB/D6cr5QnYUQzvxUU5G4ruAcW4JoY1SH/Tj5HvEZj6px76zpwLWUQ8UXJISLDx95nBX2oOd
NwHQPo0a11KTY1P1LvGi4W1/zw3mMVDS9kxgI4bOVLlOAfi06vfNIeSoLPa7gnIpLrrMOsBl3JUj
8zMSAoFWOadcZG99PFOghE4mjWTueFn90ZF+nlcpkwgIBHEBLoQwN2rp4eb/k7BDs2qX2zrHWJ6M
iiwKEljH12Jhnu1BvktHdMvw5NiyMWowYeyS+/+nBubTpGxsmvIIAi/TKYhPxl1F2vgMa/1sSs5J
uoUCO+HsDLkY0Qy2JpdIYyLXLmPsv4wTFSSEx/QVQVG0Hjz7qbhfvyDPwkyeVxsUHvZdQSzJR3p9
vFo5pPdGUNXE77WIzNmOALkXKAmJCA/qeyZxnOs4HS8PGBuVRTXIQuBJ8S7SxdGUkNxRFwH1WWkp
X/iVuysDTi3AeN4RLw0GwVOl+v64a2i0/4ly8/3Mq65/4HL5vYsI9Yu4mqedqr9KH0ukeQo44w9u
yaaPIeJImlDy2osFm506YuAcl1XW/8nKc54EeRkCn6MxrexyF00HUBA6ZBSDfCyfOFDTwchpoq9V
7dzmHKYfDRdDwICGGOLypJqV0pHS1mZrCyT2GxddcO2nTiwdrAWQcMbQmBkaX5S0efXGYXsJUedM
gnMAKqrDFZ33qg5u8sps5WhvovnOTNNCm2HcsnMvqL1IqcBVQPtZU6gpw5jFy298B4Qp1kmIjrr3
4ioMycVS39YL8IvQrKwni0/plzSm2CviecLS5lX9nNiXrbGs7aRVztf9Sb1CmvvI/3O3Wp4A6KSS
xmL5WBDsTOIkvaXXg1bFTabdbfWWhV1Dtu8yplESfPVrTVi/YAtursFR0ES46/zDMDJvRftDPXgi
waGansval4q8cR5tq/tf1ZKimKVKjq+SOveopzBatOPNzgCSsNYqiq9hfY8V21CeRiNEGcLGQgRX
f5LDC0xhDyO7Jitt40wpN6NqenfanjeJTnp0L+Qhlc2w+myMAK5X0L1rovCywgSAxYFMPsU66Tgt
lUNXT84NPGOHeod7NImu0JX1CYrScG8Q5In+41/mit9nui/Yv3qGT50dVwfTZ4ylY7E6T5DEW0v4
55iaanXQJfc2xoSs6H8N+dtebmMCGZgZ0rJ136KzdOGXR+V8RnJiU6frFA+777e8eW0kx8prl6+t
45DszlARA+e3gfiAX8+F6JrRl6n7KTFU3H6GI+13ITyFunJ7lTMwOsfGV233+S71kY/5Kvti1BB1
EfzPCPBCbH0rN2AB0slLdIj+3iCZWEIpoWRNYfb4wS3QQsa9vB3NxmNC+4BtRcsfC0q++DEQLfVM
B2Z3f2RzeRyV3h143Tc3lYmEzGgUQMAZHu4MfzQRvn1CuVwBssz9moF4j0m/fEa0PJiyK/R+dBCX
psL4xZgIEDzYtpdsBQUXmIjV6zJTtb7pD9Om6HpM2/uoXGO6oMQzPiMIflgVF1AzbT/DpkErRQog
vClz1FbeQL4BuaR+HPkUwBW/JWIms4RHeWV/JSJV56EDYCrRiqzeVO9pGl5i3yGIoeitqp7H3z7L
Hlc0VZ2Wjb4hkAujUdCAAcYsR8PGjIldh4suJo1fX0gNnoF2lRdmoSFbTR0uQ7HhUi4LCIXJrGnb
xgi6cW5yV8yORvkv9tK9OGSDDyT/IUgN/GCLa547W6V8/fHI5ostDjTK+K2nekzqVYdhtDmB9JNJ
D1F5VUudPqbh9IJVFOvVvY+JfUHVT53sxXL/L80yzCa8JRDc8J0cyJknP2VHz6SyML8uw5ohQ8SQ
0pQctPQDOH1QVWGTpv4Rys9IkydzbYgBIPsWl4p/+/z0QNxHMIVpAD520E0gZu1ScDf8OpoyrC2u
P/LIXXuf0zFEIj45yU5T3UW7GYx/u7HR6EQwv+WX+GcOEzduV13eS6i3Oietg/BHsx8F64aKa3OK
+T1EiEBNsG4qkj7wzAr/1X+fCr8zdaQCZAhkOUgOJSsOUn15f3z4lZb1aHYvdDqumtx6HfCsCRT8
3Ygu3/uBQsaKvdJn0g5P+uamnrxw7fcpR1MW2nGt1DKaUhTY0sCHuNYXvQ7p7MacrIr5eAVML6qe
RhfhVcBjcxQlwgm473XWqjVu/fbRnLqS4AKed4aROAbj4nhFETk8h8tDKduBPATKzp+ij6zr//CT
IxjZC2d2dB+hH/Ck7xSPv2JNJrEEEDKbeFQEr0GVz3AJTL07zmFzEJG2IscgYXTpQMLP8Aqp5xIl
CjMWloGjRrnPu0JtfIysxOjFEcod9t2ReFDtn0gurKay7yBhIuZW2h9Eva0LUYjfQna84Q4wwGQP
Rop9yZNXjb0C7pZ0rLjM/NW4d6xBxdnelk/gCDKFIc8Iw0jltsRTXrcCHtbnXnalkhNs7nqsJdx4
rwd5diiNyEf9j71m3VlFLIBmk6BQSQkinOerR+vJYWAN6gPjOZ2zGyVBVLoVbzjnsT4FXLAhGzNm
BYOByFZuY5H6IR1QGbxHRouR8SgWIjPNVOJmOc9b+87wR7br7cWFYOfQ4g7Q2AoxNQ5xqefG1wP6
afTKyAnhz9hmg6HaktPPMpTpaDbD6JSEqMylsY6PoXjUGrAQb9ZR31p25ggL7t5gPA2Zen2xB+sV
JmVfmgc4OmBQlQGgTB+/IWczWk/6ysvbOH5e5gWlrcyNpzLBa/vVC56XDMlY1e55AAyUy1fKtybt
xOGd0MUyitqPQK1nmu3b9Vcb7HctguKwCjLIUhOnZjYWZN1DJw8ZAmMPIEtuxHavDK4FFzYu1i3i
QsvVeFZkq4vjxYvAyYjgjd+YVafABTkdmnck36TdMm8jCB2T2PIKigYdZme5EhAc5Sf6xOS5plNK
0gtfxjvE3wZanUdUiepVo+k9X8Z9eBLbaQn92+TPE2FFHcDwv6N8OClFXv2/q7dniARCkp3TOm1Z
QVpO686/h1BrmMd86UroRnMUYigWwLLOnApYeRU5JznOi2oxl5napULMWWN+6AdEWOX2a6um/Kih
v204dVzJ4wAjtGYmwQM6/z6CVQD9dEQIx+nATOH1rA7li+6eG2RkOGCVKHxQ1LkPC8A0P37Tq4Wd
3ZMS36TQ4/DdNb4Q7rVrNdRvdXteURbHhbh4haT3nVhyaAgfUbE5aGBGLT2AyAM/31pqM7817gzF
FM8z2IBBCISEVN/JVfURU7ditvSEOWuNMYzth4Tn5WZ/1DOFu0IYyMRJBMJrgbFRenS5d9ggPTrm
mI2dpIq0o534wX9GaNR3BC2H0BZNincBHW0SE2DcvHOiH0zzzxsKcYypqhd2UOk7sq3F9ZTBwXbN
T624Z7shAyhig5mE9NAOyqCfynXt2a3T88edYitcrbqkG7js831TVBxNJ0Oic2sImeXPIwdFiUD9
NvPg3QRfbGhmqJt5I60MX4xlPxGMSW4fkQ2z3lUHZ594G8cAu0YJXfbdp3IO5fVD22gXMKPRnvrv
6hfdHurqXd6nf/Wdok0X6fa2LLxPWdyy32oBawlI3RFntGttXTK713aF7ytHKDvg2qiwfaYdvC6x
6HfOfOLfTnCDdl1Mf5HTG5e6Ga7IcoPn3OTaLVhnfcY6NpCnppXawabBDWSo0Pz7RvA2DzXhGvQZ
FF5JXqsrKPcIDbLWEVBxTT7mTzuZfsH1En6sZYwyu4QokX6VMlNbVLIYdc+A8aZeBuSOrvhWmlYb
SNehrmfYJhR5sD+pS7cQxLyG8dF/TvRNlMBHBvCsqJfMY2tzIOj3nagnEKS1ZcnmSpoxtzqbL4ca
DBBkC8Y4JfIaVQG1rKIok+GyeG/g/srTSDoFmkUpRBvaHJ+J/Gw5N+do1yqafKH8BQQ7MfunYljr
4VXluqaaB30DhXzgb5Pt2gEf07vxkZDSmnxK9LmiA5jAWRN4qYqL4+Om97UKdAl0vHim7/uo4l0P
5athKlzY/HvMQGf5J46bJVz8ln+dKBnc0d3eBCXmqTcFcm7OLOjmJjALSzcL2b3G9lHbue8x25AB
5pbyKeXJInIgd7oO/Kt7Mfaq3ApLOo4tORd11unvT0+zpTuszFh/GBgxmunahjNOTg5hhMRz2uRw
LxkSROy0BJQpQ6v7k0kvDUZjOirXEjhcT3PuG7hPZxmSX3oCxe3XoLSNwONCt+ZDv0EEXJXnvIVl
Jf8dCkXZPkhbizk0lKrN7p4djF9bUdWHmyxWCQW/OlZV1Z9ITRlBvk/u0ztOar4gttf7G5PsiT3/
aP2FoFAeDH20g2tupAIkM8G/RiQ2l6uAkPfmGXPTQOqM+2fb0i7ERZ37iaFhWpC0gOZfzmnyRe7W
RuI3XLWFatqSiZBge3726sAxxwWfxoZ/gc8mxOQfrbjXtT9Ipy/pPoFdsQjkszdXRZmBMMDBVKcW
77Vf1Ibo7wnijZ+1IKJjmQOIfmCdpXXGnqXy6sCCs2/YTC8a02GPGoDzi8g7EFjbsF1MVk3Xa/fB
yhvEOjzP/4nFnx1E9gDHMtvaIsuPmcuf6FPGOGurIGYRTaBlss+JoEgFfWmMb3MjuSXYbQH5mn6v
J849iSktqVobCkVWSpN9103WLHg1F5UyKoos3wNd3Aplp8zY0NvbEpT4TENKa5+FnxjqCGQrT+tx
hu4X2pCJI+FhcpiXsMEaOXJRvfy842yPd8TwhQlDhq26f4YB55ySnyqobjE8fIW0e+xwImRLrgVz
YtXlJeXtcFIYYeKAgqtI3LLzh184Sp4j58NJ01AU4wR7abAsspiQDD460v+ivpZt9iecC9nZNWCJ
uDPO3p3x2fdqAFZDl0Z/FAh8+N4vOfRpuxugVxiSkvpxbXMDlcyrrXTYJPPRf5qIlxkZ61LRNZfm
pEi5fdDeYPouilNrIofNfPlKvk6TuUp/qvtrxZ4NL3EoQSszuEXHXmQI+hoRa+tILPU1A4uxW7p6
5beIO2mSgHzV2/G6S4v+SQNmkXiYAdCN4bHrjes50kWr99cdVDXLpDMYTA8h2OFOxSl/uQawhrPn
3WthZjf4GpRXtas3L29rHn7oiYs1F+2ap3dUNwhu5SMqWZT1EOWwN0A2dLrpWs0aP/nHlZJaSk2o
ztU6Ktjiy1lRxrrPi8YiN0TjhHK2UVwvMyzDmjzSinSjQbf2UkiGiZoeRqklcvwBC6Ad8ltO7TOW
y8cEyQtQWdpjg2Rfaa4LKT1EFNdfyNUmMViseI7ayCZs8M9cOUD7dzwl3FDC3+8m5DMkDibceYSG
Azx4LkfqpM436V6doAbE5TmCUTzojUhMua0mDyZL2xm/4dFLsN7/Fe0/58SfVBDfiyVn8CpuFpIv
7Q7MVT9FaeEA1f6BU/tfTPrlycrZSjHrhJB+X8rv0c7urdunRTDlHgasf2EZzjotg9zBLclNRD0g
9ZkTyqU8uqSNYgFG9Aoy5nFO8Tl1cHJI5FwLAC2K97OKdcZ7K9uqA7zlMeqv9DCdo8cCV8GfH213
iR1xz3KVH6z+Gmq34rtwv5V4DfKVV2Mm2ZaR+dJoEyL0K+PsRpj3Jr/SaWctpdqkcvuAvRQ8GFPR
heONKdQG3FvZUVPziH08CryuaD0yaRTDBu9SkXd9UDz5331sd6V32ReD7S5G9xOjNPsmY0aIVGnG
vxI2heOBxtkLA5+t+HEcwafsJ2TVxMkLkKYdzS3XweXLrnRV4IBfjLjDWTzUCsr6GI1MuhfdllZ/
whvSb5Sk9uj/K0l5quALYLPJgIqFRA6CU41C3M44FQnAm2QCRxNDFnOUIQeJAP6AhTkY9Eowz9Od
Ik3/W88F+LAsMsSeL1xoW31UAcXNTiOZimutcrCb1FBl2gFmTxmAyxqIy0cPXVJGRIvJx4sEY3Cp
GcFS6aZnt+H5Rze/9cYzbwAAqEnFQBxcVSMxduXNYTGs4iE6Au3BwbWwiIMqd1+dOPCRXSvYs38W
94FtDLQwaWmjLNRhu6JLj8+pPjAtYpfysGjtY9SxzmGz4lHZLdSrdfoQmYZPpnpaatKkKhAMAdeH
1w8GojJDatA3CGS6g2Kvvy/Fw7+wZlMLal4soECxf1CBmWL0Uz5QxbAmvYEcp9F1K/FoRfi0wmyR
u0rcJfkVwBIdfCXejHquqj3qpoM8cb4pE0hYZBr6viMJLbmPodG5o9S6NDqK0nJO1eIxxN4OTOUD
c2Eb+xix+4qJYVEdXFRUOSobXSVroABxOuziihczt18P1Www/z2zNp/MIjzh1NmpW2kfJeBBMwXv
Kmpxqs4VgJ6ntOke6KR1uW74f046WId5QVevZY6RTUSOLgESQez4TFPVzOYkERwstbT10z4qpeEt
47I1zoStu3q4c6V/pJqcrjnPrfeqFsxwehU1J70bUlFktEQpdkCpQTvn1iKMz7QAjPNzDakE+R4n
lki0U8M00Q13us9/mRnqIRWmPNzkE3h/KA7cTgEyklwOp+aaqVyVSS9HZ0PgPqydl/ghJgASc9OR
yQllhDUg8aC+IiRUfVmQ2oaiM7lslIXg6i8h02cDV2equDQtZ4/3oVTu8iX3LUcgJ1/4gUrbqN1d
3on4HntkRMYZGuPSQPqQPUcN3zzlNVuCHPMTGZktF2D+0Gfo5thIYoku9/jZ3uUMLVqiqQ0lTH6Y
J/9AK56FCzheawHAFQF86yWmS4yWUynlUGxMhY4XHbtMYPl5IrpGSBMgRVZtebLjNR8g/HdUaY1W
IjOJ3KmEQSpjxvcqz+Q/m6JAtLYyr8GTvHyEzoAm6f3O5ujMPEISUIt8jmt2BvWAS3c4966lDhze
8fSUldobPIgMjx3Hs1n+XEYP95MyRj3Sd5KkZ1IFzB/hVB72jF3oWYxmJ1Ld9Wq4TPiHlkF9YO5Y
s/Cyi5Sp4/6iUJR2yPnClWl1DUUY04dmTRGl3RECTB345XuGuCgg4QeHXzIgZ1RTEl8dixSuvA3d
QLFs6hu1+kCMkgihzcZmCBMg0r+Mm/2nA/kJCTjkn4fFYL0UY/2eyE8oXY+cBj4YVI6/I4kPr3Fl
Vye1tP87Szfa7vhPNkyzDLGtwVIOW3mat1PC/o5IduLgxRQz7bW3CQhEiWkzaXYMDAQlhCNQ8Hox
ftJrOeLJMUiMcPZSO4TqGW4DSUTHzODQFFy5YjCKeedHBhKPsdAyLSylZ66xc1uNoOAkK2jeLFj5
WMPAXOfqsr8RLjUUdg5mBfw4S7BKdZKtCFYmqeH577Iq07n6+OTY9Q+wvKkdnoOt8tim4GHUahlO
hiK4QRGAnHUxw3wYNI2KIgPzR6e1an4WxltFVLa5bWs2Xo+baTLHM1I+h/Eslb9rAnOuSJjAFXQA
+XT4BGnppLwXz7h2OQhECzRelbrCTr0GjU1JhlKfm1lmVl2QqJII518o3L1Tkt1tO/4wkrPYQjmW
y2PfnF3M0dReFyTx52lgnwpwz/9Zfrvb+nele0Qp0cFblzA2BuZN/9UmW4NDHB49oCiVcODoooC4
llnj9iOpvhmoy/H6yzwMt588CJRZqJSbL2XlIFb7eRxM2w8XlBEp+7DQpbJe6Ae/5D7XXPT1IR1t
FckvGaLZ8KDS7lZMkW8dZV2JNs1LYIDgVuMgvh3CJ8x3T4LcI4gtxXBILZ4YmYlMKfWqm2k/ZRyy
rdGmnrHvbTcvGwsm1KpJzcFNsExsJYhOIY0eo8TH0CxTHfBhuoywdde4wU0bQzR6VlXABsk9HtMc
usWsc0tR8NY4HfXSg/X039jfR1DbwR8XFQ1pVk6noEB7hrCNlO1nzqmhhGarCYV4zETFpLJj2HMe
fhcU9AlJ3UD3JPs0ttq/jTMwf5WT4D/EIRisw1+eyCa4AleHERP/tw6+PJxonkGqNSwHRpJyk8nN
Qr16wBJ15GZTJcqnOYqm3KmrIaUAmjNxiBL50yeg9zeeWw0ypiTHjjWBPs6M/nhSvmwWjtVV/DQw
b6sdcc0/yXcbXhnkQHoC0mXVFMIUETNjJOtmw6GgT+n8agtW2uSKHVD/J3ByDd5/qDYmPis/Ahsg
feFm+J4QVxCtNYN50zsBK3qdHjZM6NKuIfxACH391i4M646VRIC5tXHlXnBO5TNAd2BDAU3yANIm
y5GJfZjIQZxhR6AiOLumFtGWLsp/XMeFPtYC/ktTp5URnhBHH7Fu257RLDwOWe8bZB6lpENUqOQP
dEDQjkNaibQzBXJfUNyXoQo4WiUzMNz/ijBdWbytU9oXQ8Cy/dtCSnnNANzn9UPPUvIs0IRYtey3
udcj9lPJQ0+4KC9cmWR3o2IPmy9tcYPjxdhTa08PP7ks14htA4z+xzmHil1AUMOx2/ygseHShyog
mDayghf6PktqpRiltVFRxb/pHTNY4o7G03is6qT1Uf+V+UJy40z7zYHz/WarJyYOLSQRoEkNQ14x
7IxCPxMMcQgI/9LEWkHjjidTwds59S43ehsE0aHFNaQhKY/8bhuiSG64oaV0teIJP9+GJxcsMQYI
hxk31do+qhF+559JnFK/hzuCCr0L4cRgtDmZ1yoRgBkGQqY8MarkI7cqiE5g/WVfsIz5TGXyWEng
hgb2ZZqmjOjv1JHaN9EE/hIiz7OuXFE93KkzSuYV1zUDGcRgCzUrBk0slY2FecWa5Hw7bNqqYINc
v0PS84+HtODpEzF0MmER9TZ6l6zkEHt4xR2AmIUAgo+ccZJusGG9Dy+Xq9drYAwcVW/PS+YIBgdR
Ie2hFUCgpL3HjBKOnAsH0DVTAWNzYHTNNWFhpUzydfD57caihGuzpNGQdST2nqz314DYfXt3GxXw
8ePYT+KTDZbuI4VSfGtUa9MD2MiDp3mcMgFoVSefiTCX92oSDbf4Wl1EEfKTjJAKybWErgc2WABP
stgFzh2NpHNmM+zBdJMI0sHFrpitzMspDB5XuT9NmXKfnXH6eRVkcfjCTCp7XiseaqeFu04cYVUP
1OYzAJR0ro9yiOP+rmCMtWNPpwjVfUI232u72ZgmPHgP74d+3p1ofdF+zkbt3wnCbN+vKH/gRaaL
MNQf+SzH3JcZ6jfr3pv6rrvPYnys3uuI7tEFf83N3njtYhyAUx25CI/go7XOT50mdhX3C3KmnQjJ
IBsmJZqwnTp10BBpGmtg82ZYjSTbA6OwWG7DTuWA567Cjz6nng0eXxBGLD4Y4jEGp6pr6oI1F/Ls
6fUQl9My5FZe6TXh/NhyYlwO9igmWGKMYIyGdPWT+I8OJ/SKGSXI0SVObE2Z0/zHIRFkgpYKDY0C
fCAMe6Cpx9jxPlLJFN9eC0xlFCp5XGTmiYWEs3vGqpwy48xf2sBYjke3JslAmCFJCu8tSkpvZpaY
0+Uf5aKbqjKD+5lK8RAwrcMs21v9S236KMiJI8mx6ah0wkoO39Ne3XRmIhX5V/FRAefDq9BX9PLh
z//EyFd5kLaK9juAHez5UckyMsfcturgc/D8v/fCZpMOloXL2AaEomP+zZ5gQ7MNIQZ433ED1Dgu
W6q2l4kXxs/Wq0kIp9XiPGSLl0JAFlLz/zDsGwc4eHI54trXs0d6Wng3dIQUT55zHbXvbBqOckwF
PpYriK8kTywH/IRa2jAmynDDcVWQl/zo0QUyJDLwPN2fcq/o5pu52cOE3p2ICrTiIcp1MwD6wTvq
Y6kR7mEbw48WfMSxnOOhJwCy29Rm8KOR+Rw83kCmW9eH2ME85YNCF1ZDZaz/JRnqKFOh/z0c29QR
wTQeQ6C3RFqiNF48CwF6LIXZQVBN868tDPobNKTE6AqUooc2HjicmDH7490gtSJvLarZ5gXdjHJB
EMCrW/rdpCdTCBRRJJfzreROGkviwzpA60bf6guY4rsgjsIV/Da8BkyiCemLabKdZ5YfM41OClOs
yHM4NDmiPYfO4ZRTVUmW8SEcEsYpg5xNtdM/qYCRY5C7/Dc9ztDz9CnDWkJaD7JdTDI/Ao1DudEc
TYtxgYUhpO75uJXrM10BBYt++xDJL7IbOcKGJD8zOubDpmPf3Uy0UJXlmCt7aKDV0ughdie9dFXB
eeGoEWaE9r+pEI6D4RMWMQydAqBa5rRmh76+MnECUHAmU27euXqPf+Fq7aedMT+vlwI/WSdR9gAC
yRQzwDemWqtW64Kteu2uEl8ADUWmm8Ip+okc7A1M0Ry9cMh0aTltY+7vyrVBPI36h2TyCXNY1u1Q
pHydZydYieHxV19PuziiZaUsRPUbUKX/PBWkKEFnmOPKvusX72MLZVwnueRpzfd9IEMCG0paTmWi
Dz2U0ELpnwY0UMOhXO9NJXBqJFYGiIpkjNl5/k/warF3r03hdVHfQSwBZke8h/0/2cdOHoS79Tiz
1684x7dkmct7BZH18I/MuO10STc86a13I1xwNTtdcldL6Pg9SynMnKjv3yiP5jpfNnRyTb0pBJei
cg2yQNfe7mrTM6+jKPz1ENFZ+RvbaPejBkNVrnkvcxGJy2SWNC/0e9b3k3/OZBqoFrNw3kBxabiR
+QG/hAbGwsZS9xl0oYLhX7qYKO6Aa1KnW0DyTn+VXidrpRW5OIEcP4FORYYiXIFduHauowW1y1kJ
rDoscH9vEli9zgn+sRervGEKr03rPdubmnY8uDcjcNBp13VzylrRO7X6Pojjv/ruz412XAqXjZV1
9DoLKE1wd64FQz8KkiEpLZAjWosqRpKnOH38lfeeSmiJW2Co7bmTeHALcF1BF90Sg3Awb3bIuGFJ
5jQMpwoJGwji9IUCpJ4O6RE+/kjgbcIDpeuuOUVl/5zZh4nOASlxm5egMSnGLKnhMn1QOvllN71S
6ijj6cBTI1kKvyU2qqdOfka0IwznZZ2jeB3hl7hs/Ib6deJ7a6DQwXQ9MwTBPRkWIsDd79/ElrnP
wdYQ4Fyzx22pOgXk+dlrv4OTYRTTnWNNdomoj0ELKYjHQ3gVInHNxs0NDZ2xBkQ5rwKEpPOBLX3N
QdbqYR/+6edQ5w1WGwgUmWa7w9WuG/gIb/WJgtASrE0Clb/rKBxLbqbRhtslb44ruMaObDnXEY+Q
1rxDaAHocFeLcYjGE3U3eCnoC50EaQa/Eeo2gGaOxVOBSFve3qs6/y6KB/a3pyWX/I7XBe+DuWDf
7AAlcii/gf9OcLOiOObDl/UpNJWWMNTkvW4Fo3n0uqIglcnpXuXizVEpSIx9kL2UTENd3WXUz7jQ
B3ihEVBUG4p5NoSOFy7NIeMRoHytI3CrELMhQX0XpdRVpmpJ9QUY3mlj5Sn4kdCB9RqkyyzPLFGd
KIgJibJa1wj20ljc9UWVWjSOjwa5nDQ/2NetGasbH5wAa0PVJ58lZcihh1xn5TvVE/wJk3J/+Cnn
OSP8A8HiGPyfqyX1A5SKgvvrN0NKyx1iJKBorlHA8ZmNFDEEWfkJNGhJJGQf42TLd4TUIY3BwTXE
oj6jLS9gutR7bsicbXx0TF/iXbSxCD/VX2rKBRP3N4nm4VC3AFH/5MAPG0rY18CAQLcc9IQg6t2y
0+Xl1txsyssh1GqomJU363yRWFr6avR+N/jDRjqLB/PjxL3Z85Vq0G6CZy1BHYHTlsyz7E0dr89X
WgprAVOnqqdLwnbkln8TXjvEYPgT2dszNQxoUTFGtKRJbPdOt+vPhpi5kSJ7GAl757l6+TmiNqLp
5fRU9ikowbOFBTwWzyEFnAgp0dvoFAAkFixPxgVdHo4dMafI21hi7EF0fBE9Bha9v9nx+vnyBVDE
rprqsjCC+BJXUGPf83cTc8AxzZUsYZvMGkECtvDcnALaR3zQHjTtUzLFGbjOpx4LraR+wXxOFR5Z
2pQMLk86g/tuVE53uLEKXqX9+USy16wg2SNqV+1jZsFQrBhykNO7gHz0U9FGsO/el7ekYdu921Qe
D6YqlZ5b4yIvh9ouMNrOoH1MWUXIEPe2Nnaav9uWlXUpHhz3D/aTOULw0Hu9itwsD9iVSvhDtxs6
4dHJ1wcFbg0bI3f6kw2hBm2Wqi/oHvg/l+dcd5Wu0OdCeiKH1mZ+aXhHlLIEqVwIj9OZzuDsTSkH
JojOeg0Lm5BjyW2QhLH/L+1dC/8rje4BWtMGX+xbuzwwN62yN2j+NqPNy9W+JSPPUmkC8pzXAcF1
gfQIqGoI6+prOCkgxXp998YC24FOzthUz5Sl2M565jgjpd0FqjyQzjuMIj0VbsbZwTM5C0eM+59A
jFl6G00Uj5xiJISJc1V4QASHKdtYqtOhtAOehfM4+KBUIwBl3TNw77AOjLUapq0aZs9Mz1wBMyCO
AwJ2rgmt+E+Nt1DBnD+0IKipqmWBdrFEgAWwihC9JLegqbePn3icH3uEfBNI7q2ExEr5tWtIWlxv
6x/wd24lc7Sv7l5LnCRecNlV9xmOq8+EHJZ8g1d4znlrxqAHMUU7LLw+0m3a7wSmZ5JkA3Q3TM9e
ROP77kcMjypQzOIw6/lbYbgmzYbrW6w70PMXwG5F44ibsBwRuXfAWeHOwGr2LNwRyO1z99L+Ta9a
XQ8tCUjmAyEFmmM1lPa81DJbDqU15upeFkZfNm/Krr2ivft5L2jiKbzp1oUFG2DVEPVcKsGbopq5
nGjipruHWk5OEfLaBg9SXp2GO4j9gzdShxRYyQyBRW57E9ALzZ3PAo2pBDd9uVVbRjmOkFD0hm0S
LW8yOT8sZ6eI4PYR1/vMaGp8nGi8eFQqSuRU6rjzIwy7FthyygpCgbmo6qQ7qgIw98soRMgaPPJC
rtgIzMap+6OblIPq/OlUsLOZvD5UfaFgoTt7kwRyjEfpFWxS2URAMvAYOj+rNuM+New9+fzMHvgL
G+QLeruP8RThOeYY8DC5h7K19F6ec4BWs4+Pgkz9TFkirXthE8EMDOoHoavdr8Eh/rBsQV6ARWXY
po3pGc9n3gi120FFOBJ7GP5LMfqMc1kR6QwYIy9rH+w8mzduug1I6g5VqvdTvOFLRek1TNdGZjZ+
XPo0iFYehWVVFJ9BpL9bRir/b512E7yTZNkG+3dHgTFmfPbrA6cJFZathoBw0jWA8aMaBDJTA/Gd
RgoCfnBnx8PA2voTlJi7ftqwUwnZLnuZlP3FEv36bKuVfFOe07R+tdYVDl1Fl8zqPlfYhL/2BhA3
yb3SOigt5V0ItPO0evWD8QVP1bBsddKld9+7TMXksQq5MMwpfvnEh/wkn301Wuj/vsiaqTyjJiDK
UXYDabDsdDUSC2qCjom4Q11+Kvxh4Alkb5a9q9KMfolXue+ZLEHJyi7kR46GE+CBCdCR2EJO4UB4
RtVIuj4wLAfc1Z6bTvAAyxD1Wi67dMo2Wvot8gb0xrAHsBGwHNJK2Ba1cBJdcgSElRwKJAe5rsAD
RtBIS3DubZe+30xS55BzNei592v4qSB9isWOWgRTRHZwT3d+6Tt6x+ijM2QyXsZ2xB25TD6dw9gv
/HE2qZ4RmvrZ7RGZiMQPOCCcIdhhaZm1B7dC+nG6sKcHLEX9maYdyAlV0dr3jHOeiagET1j8RFeB
ADFtjz9Kb5bjdLxjfDPv6SVnxaUHM13X9neLkmb7eeVonk0BWBSBx5FZnBFx85GN5nk4gtNocCkM
AztfOwB+v3zMnSK4C6BP4nfZxtIptIuEQiBA6LxLPAVKSh3V9inc8xcNDh2ljbg9YDJkbq5v/XD1
2Kt+0kPRzJwdctM/xdAzuIrqbc0FE4chjjPMSP6nDLJ6FZH8UZCp1ofLRjpgpklYV3qbMsaKNBA1
yZKXUk89AfYybWd6j6amPdbwFR/8eFP1bUOWv7eLrmYAyYeJWxtJ5FHcdZYLLUF+W3RUVqdEQdLu
P0YpC64NVXUuAYHVqSP/oUYY5PpIEWjAcEHdPK7yFz5bcjKkTyOZMPjzF/msyqqru1JqvPJXRuJG
lYRaUBAemTLZkuEuH/5tJ5SOncqbJwlR9QC4+JiKwViArxSYChV6R9wIFSyaKjvouHFnNZzlcKCk
R4BVixc1SPdBU8pk/VhttuTSsA4b0sFcOS7CzukVUfjMop8tQi2GpaG7wA7tyQnn9iRgpaGA55Zj
vtO8bVqkhdXBOGaTh3xl53ssMiiKjFg98voSzgrVz+vD36w1BhRLbVEpEYhB3Ce6Fd5bm3Dj7nxr
4SbmkIy7YqkREpDiTkx8s+lqJnpCZIQPskJJVEQIJbtuDLIW56lMVsjIpkukz4Qe9ArVxCbqTfaf
qfg4uguOnFFChSULfpz0YbdV1caFUrNk5Z2AgDP6xnJMTkmxFNMBWrRIHU9vDu71OaJ91VhB4WIZ
6ZVeE+IskKhLk1ZTr2hBe/K64qY0wyNHZt0T08JdnctuhNpZssPZ3dQ009O8oqGzPZ2kKcDuTY9o
DhsWyZVZkE+RR6tKxMdcGXgauz6sWIxnSKitqcub63iSh5MgYSrkAGNTUG7J9mwv+LkJkXxQcZTO
P79JbkHlhHGQi/td/f3J6bFnoo9nxmjEvW03QeTKdIg3DB1xh/z/oADHc7Xg9c0Wh74nW7BJihbm
EDviPbZB8fgq6lb7WDVaTIVvMgtAxNMfS5b6K2KuMb9yql0UzCUzKKoMEwPJLZLJdP6Q/e+s3sLb
1+q2uFwfcRI17LNDtKyx+XMBhmFrOFPQn+BrF8ejTTNbBVUsG/s6y9Kw+pFKPDgt+PXWPgx72GLI
W7yAvKpNdkUBnrJle1+TQ17OCa0qBaG02mCQ21cC1ALhEbgCzsL2+A/NGTdSmFr5IZ4rd8Ty35zM
+sjOnyDvq7nvFLRKdSogoV6OAGnazmCdJJXrCzoiPX6n4dLhWDh5fMF+8AEZGjR4hvcLd2God+sM
6JTQjQ0aXCQqx9dlIKn5Hj62pw0Uw2acy8c+37oW/9dNLNlyY6hPSoyQo5KTWvjb/GHnKLCv1Un0
dUzM3zyB5/+31zqX03c8Z/lRJM18YOTzvchxTclJccgvpFQbBsJjxq4kve1YahfzaBHj6zFUIDwo
d87QexIrifxs6kN5qsitCNNNhnBFM/ZIgd3JlKG6flOWA3uQRwxxvwURiJ5shUB8AL+/Zdthwxe4
x3AcXyGFjWE4GZKYyeZ7Baq/+/6I+Dn71iXJbnEg7d03fI0KBG4OCahS+0KGlOm/3BbcNQu/8T+c
JWyU9pITFoudOYlwbzDHLxXrylR4TTNIOIok7LORkk09isJl1kcQ/r70wJQw6GFvdbp3HhbULawY
xabWWFuJFyhsvYxWeZ1hwM2HVyWuo39r61JRDLW27MaW+gQwocIeBdfYy3TOlnGWHLqHVU4y4JxV
sCG9D/iyjTXCKdtK340alBsmgr4nJM54DgJGXhx3RqV3zg9clc2y1Kkn3pD4ugU69FDhS2bbc+ve
p21C3jY73rxp1KndkMR3Pf2mf33ldsGhYqryHWe0G8VavCSV4qOf77yQwSit+pox5YXhR2Sf89cY
Gukeg0+9efsyN3hvDspn5rZKbx5oCgR/6qISXPnylAPmA37kRtJArIbwEAVaxzbURgne5aBMJoQc
5YvFHpuvjDaDB50nvZuaf7ugmOHej2x/cmz9hDUjd0owmyMnTu4Lt7IXMfisLxuB4wXrvz91EEIk
epriHhCSPh4v9HF6zvccUqUT4TFDlt5JrQpUb8a1PMhtXGGUCuxbfoAnt7MpWY6f4kQPU4LSmITK
BTPUHsz22+gCEC0QtERARu/iFRzJ8UAdu6T1oIF9jo7mqkpSjCSjdnJbTIqDnrDbsSg0bz05IPDI
x3CwPRGw2mOW0dWwnF0dGOv7h0RBlWTv2LKFCUApTLIesXT+BrLFZK3wuBKdlFVc9Z0as32xw6P5
Z0U9ed/J04dsMRCfeCRu8lAvQB/43MmIsZxhIY2LCoOOM8ZCQdh/mpPOz2GBgi5kki1NHOu1XSLu
yXmQBk11K9zObgJBYZrouq/YfNBdNyv1SFY5Y4XxvKxvhD4vQkjkWSJ/MqjIMd5RqxsY67BiaxN6
GVk5HI4mJg0d0Mj4JN8bpLwx+0S3Ibnd8+gRszuq4Xc3NS80d1gig1tbANgSDvkEZTCLGKWzl0mn
QVJFBK0Ay16Yfb/+6AA3No+TKJ0hOlPTvZIA+/u9XtfRl61py0XIWLfnsVYkXv/s+SxmK1Im4gad
HY30zGfuzI/Rfq3pH6eM4Oc6uJ7ej5Cw4yLyPfrH/YW8lTGszsgBHKo+3/wy1yI/Gz03cP09LMI4
VBGY8gOPLp2sUmAgmUE9ZcFCZAVmRTAWgCjdguoKy1kcaS4xKlh/3vFijQ4aA6oPMDbzMNm98fRN
FcUVWHxJNTJfW3nUlMujjZszjLxzM5pZYiGHMVpP73R5riEU9odLph0lE0xlfWri7rM4B/bT8JiV
TmO0D6bLIn1CVqHmSByTPNHPKtWqvzc9Nfv4bv/joYML8Qm1TjjaNzlYdSdXVXKTA3SEHih+iJJx
AR5EnIX2icLYTbe23U0PZpPMox19yL/irr8m5TSvNp12mpANOHuhznm5vKCAiOjgsTzPyh2yrgy6
MQ3RfTbwxM8wnX6o9vocjTNRr2qVvUL3R6x9YoRq4IBRXfREn+u/nGHhMGBNYwBmGkfU5KDN5+YF
6PGKcZTxhiI2xuhO26HIgnS9GLMRC2oQBoird5Ul49UnT0L6Toxbj3ytBU0KMv2fZ78o808+rRaw
meOZBKheURsl4FLUKratBgZL7AR2VC7XBcVVg5XBaMcXqQDxCAqfjUXQBAaLOxDGPEgqHv/QbC/U
uJ5/+ecRhJ0ua1RuZ4NbpihWVZzvWs6c9p+GI7seqSd1scGaVeac8mY5DTl99Uw/l0zXNgmiko42
8REwv0tEeIoTVmQ6fgCO0MtvDjCUejn/YsExlBq3kNNi3PnmlybbjE9h0HOceKJp/Gmpk4/Zri/a
rBv+/T/FYWVBmv62mg/7YMmifPddWpyKPdh2fwAr2W3E03gN5BKxRcH3ECe0PfpTVEqwXNJ699wO
zjFbWKplXFBpf23cGDPIo9xBbTDNXI+2SRAFDJDZE1QATsqNojRbWZ9XKrDObpQrcykRWjHCDYTG
zw21VRcp0nEPwUyMdbLA8zOzWnaI1gemCvKA1Ed0bJcH6M1KCSpl97H0/COga/zBhX7x7dNdNSyl
Z4HN5VfaDG8UBSROP4Dq/TgTaIT5l1opts8c91Mug57jgVROz42TZORQDwbUpyIRC8O/JKBYiR9/
kOwvr27WawSK1eBZaYwjqODZLBnXUgEp3X2iUMpQ5WcSyw07Jl7lf8lNqXeYwp0My2REL7AB/w60
rO3FrNPvtw//lGUEZ4np86BDpYPc8yAets78fjnfU4pIOvWxgHy0fiw2kLABXT5x59t7zTucHIzH
/KleZkWPCuyT8KZXRXBrm2xYgKra4ubbrDT15V3qkDZ9XzvNKgwkp1ZIg+IQdicbV3UHrTqhCdt1
30LrFklYiYuhky4F/Qnkm/1zYw/brXGVX3qpiGzWWs1xHIdv1smJKf72/AqSPQZMh8z1t4f6MU6m
E9B3H7v/wcHi4SzUievc473U8CdF3zD4UMLMsxR/14CVjULu5C1BhWZoy/D3D5IlIlPzXWjItRcX
kpLV/hw5qfNnO+3cgoiXwjFCf1MPfiSslIa+5tjZi13oyV7RIqIJLwaSM0wfCwUD/+GelI8VLsse
KJ38uvbYty08SsVztvosDWiDgWk+1HBDtmq45Li+pzd/3928nqYkPT3dZlvVv/QDSHm4e/g8Lc3j
CSsuWfkjjmo6burMJT8KbEQLp6Ib9jMDHbBE20YiP9qDkUJp3uRZoxI3dWyeSqzEhR1B05Bwzw3b
PAVAfTllaDcZkWNWq7uC9OdLzA63TXdhpXESqMMygvk8Ivf4kLN3hpqxvfqfNltRzxFa5667/LvG
Bv8W9kHcw3+BnEZ7SdQUklpQiTnjXmAxfHjVwN/ABBFgF4Wfe2LLB4CXzkoBrqeqwhs3VFK/nJtW
Q+33WDCVqxyDVFowx9OpW98kku2XEO2YTnbAodgP3/WCqKpfNkJ9MuuXsQwaEMtCXGMDdXAhNiP/
Pk7GFasj8wv5Od6bJg3F8MO7jQw/0Fk0vNrxfGIRlwCDNKgqr2wN3OvZ7mFo7lnAIJffJHDxOtCB
ZlVHDmM5lN10H0fYqdXb6lcxgfRZ3JorcOX3WqkHI1fUsCbUwM322ROLR8mKNU4zdzGYL/cR7R1z
zV/DnmuX9ilT0e23DF24XQGPgi91gSzmxj+O2vh7B7fU6fmh5TmitSkjHJsnfUOgi997wkMrUIYv
2HVdIKNYrr4OzPqxT4Qe4E4p4X/8gx4d1L7vUlebS6mlQKhj+dR5JHFDBjbSaEKnpZIB6vm4sVit
6QSbK4MBsMGnJN57OR5vAVKcsFWAGyni8ytCpSUYgQRkEB0eyvMjI+XPbxE2yJmyCqnpMxd9Stl3
S5/lD2dAPTQ/LLJ/WRXw1Funoe4oJ4X2XZy5X2AP5l943BRZ5B4xNmlhp+Ix0kcZJGSlruHXciFu
3mgegLXNf80tH8dnTi6v7Cup9PL56GmuTbOmq8h0uplcwkpvBm1cC9zAUAqP5Rtezf9aGOIzPVlA
5s1XY2sceD0lmN/DqIgCOwnIh6+iDJgKC97T9a7uc6/MneF7vAxqPbuCeiR29S0KPuARbEZDYIcb
oVkUnkNj4ug26pyGjgKMHFbB7Vxd6NsBYhPowXsk9sXG6nNnJTuZAZMLHnjjkPAklwZrBLdajkfp
ig3yXh/4AmYb95imlrwvhLIx4SRAmwiTAoP/JSUJTb1tCmea3hb73cJCbXke6EJy+34iG90wIEfV
zfU5OhybA0fDsxgB035vqfkzCc6KKOBB3RF77vaA9UumC7EeDz+7YXYhAcuF8NLkXi3FwEdq/B6J
n+ilRx2y5/VoffzVk4dC73MVjBYGAVIkTy27L3klifRBsHBItrstG7sdd2alWVdIMlqcQnBjax5b
oUrQ8PWutwdWLesBCdxAJE5V++Y3WM1ddjv+/VADh7SAMfWuf0Unncyc1oGFwYcs2HsW2SFuG4MV
5uu4GJnlNUug1orq935ABJTUKuIMQRRnEhKhYVXBzZf2Toht9In9Ycrf9NqcOfuiKPZ34zeU9AcC
z6I5UN9Z4xOht5uWe4TgbDVCoCpEDC2cGCoHmKy3eSFimuJNRgJ+J6yqYw9tKy6ymJ0XjUiKGoF3
RWKdLMmDCbnhXEAGGGUmbIYcgGlZknAolAmR+H6tx/38sVK5LBH6OU4a5O5SvHa8l73skkICvwf/
ZljSeR1EuJhI2ew0ZS+84mpROuVSf3waADPY8YSnudygMPo9eMW+4nZmVH5Wg1tse6XmJgseTjW3
W5h2nvGfRutrSxdxMrKw4xHq5p62cnevYEorB5hFPkUI2qvWwIM7fvDdoRPTyg3SqV2CTF/JwfIG
OlRhbDJbbuvRKphno7aVFyP+g7AonM28uUzx7DrtpYREfBxvDpnXgAmoWHxRgQ1b2s3RkfOlphsA
ifG+alWdpFuVN4GyrukWlAogcQiBQfQAVe6x7F+277aH1SFb1xzpcWYtWSJE1mdNVlNodbxQPiYx
mMSiM9DcGg3alFJqBpMujHISZB4WpuulR/XcRU1KU68xrHq0+SDN5LfJLSbKWQ9iHDB0BaD6o1Jg
6loBsSOGLIXPnOewLpVM3gQ5bE8jKbJWXFNPyj5fDiV3jhlf2XJb3YNBeiXlXCLZMCDuEBl5aSmq
TJKhkmIY9gCCD8pRQODH5JINwPPqlth6PWdScY/mAY7sfPOtBwH+qGjH+N1PHuVM5gF03tlEY2NQ
/wCuU8UU8iYo6fur8V0A3SSIYSAliGfSHnN45sW7YoxvFaopN8+/dhpBHaNdBQTPvCOmXck5+DhH
TAMiGGm1j4LHi2QvKg1S7uSjHAba6AMkunbsMwpO47n8+Xp7HH74d2HkoiAhw2nBam6v9nxYVVCR
FzlOEitXuc9jNVZCPHDJukbxyrA8pU2fvj9dOan+p8M2UaUBsYLFaTxrvsrvXPiWdFKxHXWQ728P
4PCyuovbC0njQBFEi0d9nR7LRE6g1GycFXtudkntrG8Z1bpkly5sToP4c9rS4i6GvDzMbjhLYa00
AKq/DLxTMYACSrgGZUN02J0DdvdIXDx8U+wlYj6bwjDFh3GGjLWHGULytma3KE+Kp23dayjuhFEs
BVqM4yvNGREZNmD5PX0RkBwH3bQMG+nGK11la/AccwHYjPZ2I7WH3bd8YIGdtd+LD8M12PxXIchk
DmuqBWMCRmOWJR7Pr+XDXbESt6s9uLi2f9RWfyiChY6jYHXfGiRNb6gGXNcCnpOnHbIlFAsgB+hx
gmz/yQ/KseaUtpbaJFheyEbIbO+YnyzSwdbsYU7Bmi2kbfD0v4lvovpC6lcJkm+XZ2DNZCrwG46A
NluEYYXFRGetQzM27ypBzmkMC+nA0RwwELzA0JYz2IVX0MskJKHLch8QjR00QLHK3ur9LE/30tda
zd8rr6qfj2FikTr0eBiI5NL35ZGsiL3xbo9PUUC/1nM/O4UWB8EbwahUq5PhieICJGA7tlU2cdEJ
hfDrVeldqDg9kmVtSWEunszcdzZh9LJZZO6tX0M3PosUh0/c/qFWQZ9QES/xZxv3SUAHCcLMZQv9
BxWpMvjZE/BpXRVWjd6ZDq8qxubCHWLdBHAqlXKPua/byYiFhGu/gMpUYACYRXHh5SC5yvuuxQZ8
sNFLkLdz2T2QMm6usnp27yZ99ade4WVaZFe0VKx0R9TXCTaCXIayRsBQj/EYbZXW3IrzU/hP9NJB
WFbK/ecptL5jRICYsLoO5bKBqEE8ianXU0dLkq6tMtGH5al6f1xR/TvDMk2Z/3QA1KmX48DgZJgP
XtPSEADmolKz9uViQzn4DLt9vk9d0DaX+yhvoiBK3UpGicnpJij2CiwvOZz3vNAH7X3vEx6TgHsM
WiI03VvBB2oxFD8ASI4X+kO4gDkoQXdyUJsSAXigLIN6onAgdsThWMhn34NAvYR5QuXjMpD5b0rf
oLYGncGdTMXNVFzplcYM7fp2WQ3uHeZ9+EzAQMn3bVb1EISLVJ1kpIfWLwexBzbOUJgjofuQVLTz
qAweexFtd+IWQ/WzL6QnsQPH0OH1fhdw5rARXbVzS//52ObPD9DpDGaPlOMtPhFk3yi5V4JwM6P2
93K/ZI4Z2/YBITMwLfAlcjVYVJNIKHBt31osVDWlrG2O32O3l7VQfswabRm3/Ng/xst38ysK+WR9
pbOANNfUMUkqqf/lG09060dv1zunhdV26GQYk7V4EWU5z8HqxEYJFtY4oOpZbfnXz8P96yK7T2Kw
AuTrB0FLs2qty2QxnD/o6Zpqvl8lYrkpqcmyAKO+k0ILKRzmHjQfIpiJ0uI9e2y4+q236jZ/eq6S
SPIUH8384EKUX/VcCIl0QdgmWevRHLjQt7bPQNReZ/Op38deBt+B1mqwGQjYO+xaB2njdwhjOX4G
rJuYr8WG7sIWQdQsH5X4fZvKBZI/4N1lB/zljo8/B3SNL6H6cRQp3LUvrEMDGX7zpeTQpwwGe9fv
dlCIdQUEDHAR8Xc+jfLxHskl4jmUQUjLmdUSkSv2xPb2rB+l14Vg5ZQlu2qaeH1HQjVuwQnKrWcG
2N9hsDPvr1Ke3xjy0ZlJOyuDMVK/N7PTFQF3pxXVrzuY1g/jK4n0qi9yrhxTzqLW4k3uVy4R4qVk
gAu/AYm5TNt41uWzYUe7rkSz3cfm+ZsHKSt3eO6vSm4jxASk7WVxqf5D0PDBvThQx9s0GS4ajNo4
FMWqLCDBNh+j2iLE7wKXsoXfxegsZ3PKujx+rNaoK8llXEOvWBfdZWYZlHnz2q8mxd3ferFcAmit
+Y8NFTr0Ii2l0FrMshrPWTIlcv6em2VAnWgDAnMeetvmFWvNY1yB+hOvT5pO8OjIN4GmYw3OLLYu
9yOtEu0mN1aWEykEXl1cMC+DV/ePt2zd+lqhi3Gq8bc7MccVVL9xYH1SWU2Rfe3PJZrFBWlns7I0
QsaRmeR+k3DPCaFm0tl9EtMo1NCxAEG4OJVBynKgfJ4aeW2oRrSaiGhaBMfRyvuJbyF6enhnbiRL
3RvbepqPQbSris5a6mpAplSVU3PuAh2Gu7eir8XN/flt/MeX7NbvViFTe+WMDUxntgamBor+4z5B
Pa5Rne00+KD4390aPqfo3u+JwogbUF8lqz8V/ZFZMmBeu8X9X2sEJfUYGdO4gZLVuejJFlCv/ZNM
JHMUkQoTr45zOx0JbiZwFjTov51jEhagljOz6pN/o4/s/7r4n/pX4gQxljdmhRT7lDXjjztktE2I
2Q+Cy2orRK3Rf+1H08XQDmRGE0aaCDIBDkgXHnVpUAkIjpqosqZjVbn3Ceq4lnKuMjmjzJNT5tNo
mkcq0SoLHsqDJ6jsRw0ZAmeRzcQ4fm6yvTyBpY3r4/j1KX9qdluazTdg83b9e5xHa4ANSykOxNYq
G0X51J67pY7XO0XwU1xAYZLHCQGQWkEh+3p7+sjbsubgW1/bRDCfGlerri3cRRO+wSKVcEhi6Y4d
9eIAbiJOnKUX3JEdZ0CJ7LWFzD9lQnfBkVFuaamQdCsGjDlse5jDGLeGU/D10Ug2L489zaHV3PQI
oy2a2ehhCedI2s0TMtmr1gl1aPl6MaBhU4WEaIttHxzygjEQq7qs05Ex5bby7AWnQZ8vlIynhKDO
uHiXkxhiuGnKWO6OQF+suSpNaB6gzddZYKIScgyymX9OpBm/EGcmUEnrf/XXyyB8F3yR1NsmeYa9
eEnfdIDcHqrwOy8f4WmJ8p+aD4Qjh/u/ukFT8oFMDNA/xH1EW0g7KbAGpiazaYVewUQeO0QfHJUC
euDHcCECOYrzjG9c0OQUrLTFXKN1uxWJuTCYYHeBr2rUnpjlnYIX8QaEWec8lFbAs89BQ5Dau5T/
Mfn/ZSFWrs9Ri3I5JUat/EzK3SynMDZPBgdKfgIvcmVEHDzYOh89NLdvjoP6WieJUpi+gSSHoJgY
wdZgU6/Y9bHq6IAHvsiBuYeX2M6i/Gdd/weHcrMHaAE0maolh2ZicyfClUhg91sk+FOrs/yKXwt6
0C942+iHuHlwA1vaNBI+DRTeZQQH8tj7lRdPZVQihJvmuoW540vD2Nx8dazMZ674KNouhf+RmwDs
Eq2NakTW3Q89s8w+C0xCu8PBu665CjNFEAXM84pDr7Ifz1EkX4CRdmIy7QHA9R5fU9HFBfeBTqXF
3LETLZ/ebjqumIrpSuPjFYW3pyHPcu+NvLe3yruecUzQ16dK3uXb7rkqp1F9kRSjMAJ6TMrIwgmD
YCVMa1A8XpTRLmNdUnJDaCCLiFzrepEtLaJJ6FTb5c8HDj0atK1l32XnixUNCwPyGoaHbTbC1d24
/5bjxFxuIJHplEhGHMNslsOVHP1qZHJypWoNVUvuLXaGBk3fBJLKVw/Z4pLFf9auvARB9NKOPoaK
mcSg9T/B3LLT2vtfHkXdlZBJjjxjwSZsgKV60vAQBZvswARnh1lz8HgmSsaZD6V2trn6us7qw2tN
pKAo08rcvzpx05RS4EwSOD1UaRMm4nKPdQDkUUfPP0VQt4xeiA+4kr+i2ULTScH5SuNK5kyX9pYj
T2CGtJ2R7tnHo+JUi5StFpwe2ean0HVBl0mBZHx5I+t8l/Dqu16G+Z3CCp1vaibyfFRPrbOv/RWJ
fC8QAyUirlVBgIe+PFMG1D1TUil7VtLV2Et0Y1GidEm0It4/3GtLDOk6oIWV88xQODKtE0hmadFu
tf7BkR9Sm19A+gxSYmIFKu0FUjltWnl0QKp9/xn3pgo0KBoSwC8ADszprf2f1Nv5eQ3pcvB1WLMm
FqaAikzrtj2qPjjSTmG9sMM9MlXPM2U1ajQH5urW3CY4RRjFxKcTFy4Nedo4DAVBHBFXA2ckWzHG
oJJSjLhA3wRe2Z0+qdkI66x5h0PZUeqRR+MniPj0FALADelkh4MtXqoMnY6ctKRhvyu3hbHAUKLZ
2yrFaLWWspGgsvi3SwQ6LQJT/HiGE4LME0O07VxNALbAA46i5Dp3mp8OMB9isJeCoj52TIRNeuaC
DwjsgdnH3nlxFb5cWZEf/lbg6y8YIZa0jbD9PpO3hbnUghpOKLBJTYjm2jYa9UOVpDcnJ28lcVtF
UCzyY8XeEb/F02ehSAAIL/PVG1FvTrjDi3JHPU6yE+YdDre5ogGpgXoyDMxYwdcTO00Rn+3OrKTa
qs0wr6f+7D1kBLduWDukpq4h0Uxb6YklGVih3yWyKRPVg4zjPXqbkIxe+sTziOoDM9Y53DDGckoT
CvGOjyDv/7rNxZng9n+9x2QwTFFVQ85cfZflxzE4ru7P290zqW4XOVy7jMLPLmF8RDEGpbgqLxDW
z/58XW5zfE9x7QhvKYSgEaeYWJ9UfDMNUMKHhBTJm1LGQt8euCs5BJCZgtWOeJ8JChlq2gMzHVcQ
pzFK9YItRj/ZKwVWtoUMOCjdMjKOd+R+wQbeUaxMII+/7exJDlPD4mV1JyIUCrU8Un2q+a+OlG5E
AYJV654S6Zbb8n8pTb2jymRyeBmkT6uZ84DCuzSQwjq6eVvkKFSY0ynjVBdgvNa94DkTKi+FXlAB
z4nTJV34QiVzz5ACOfgZq0IdzvOVZ1m/hkY+tfVcT3EhQotjjuHWdQ+NEfYA8+PQ2vICtjYlDSxV
MEngKBG0IlQA9l4AcNzMoEzqKiItvbp0ka37gDapRidi4Oggcf8pWc7eRBiNHfD0vOeqrWK9ch1j
VlYr9OP2mucTjQKPh5oqkiHquKRzAT+VLxBiTlJbSV4OlFEzK50eAKggirV5T3Rj2lNyeaRFcMQ2
kr5DmJu8PLDHCxU1RRtgroXz4wmR5vQenIcFRXoXk+QdyiI3Puh+QlJgK5vDMccCaauCczCHQI6d
mlBM1At/s77MhZ72lku7N2UMyG/QTVmNEZ47lcoHTXkDqbr3/nzxQdUb8pQQkaeBzwae08fc4O4+
pIsWz8899E9/MqAy8+o4GiYu37b1nSrP2ZW36s+Plgpy80uwHqbZujjecL3QEnRnpPvBBkt09q20
cHINT3mnGoJHc/ZxZwTUDzQXcHFSMZYrYvOqyj8PyoBI7ydOqguGYqqEWXScso06wYBm0JIu0TWa
ZA0GPvcRu++zm9U1DPpxcqsJ9nfzlfBT86Ftbd0oTYm8d7Ha3URAPZiHLUwb4rpBkXmchDGCUP8H
MQRvgV3ZoJssi7QoL1ZKgerfDYGs0ltZ5rJP5qhqq9SFFQGanKv4rw441py+4PMxY0F8uuPvw7rv
ynuHHy4MloQD4BykpMMvMLpVbx0/ET5g00YXWT5lZ4D+l2IZCUCiDL7ZiwPGbtqph2kcsqGmM/M/
rLm2ejNN9EfPm2Hug2jQRzo3C4iL/SO1HscSRUEDIlBJFTNhJAFsWRIR3eWMZgMJG+pN6J44ncEv
MJLtVumGf+j2IQINLc65hmA0MfPnBCn3RzMsC0Sy0vTGHv+uYnW9kTybWZEK/BozI3JbizGKEf1g
5EpNz76RYHomOFLmFoQWSCKJy6EbMuBgd9vbGGHK6//QtmnZMcI86M1xt+onkgKNTFTXFv5ckPS4
Xz8DNQ+djz5pCQ797467acDWNRyO9pi6mOvqpPfVn74Yp2fVJR4K1y/t5Nfh2BzPLRWNVXBhF581
Fs2Q6vEHUvMUTHDTdCwXvJI3fUa5XkpHH1N7qiZW3cQv3gNTZp0SdC96tW+0vSmzeWxOkV3mD9wF
XlMaxodOpqZYihFP0RKc/Lm9mTjip19o1Gdg1H5h4KH7Bn0dJ9y23cH4e5mdr+lGoLBr+t8kA5eW
ephx5GSzn3TwUbLMZ2u0ysXGhb1lOe37Ed0rUpnoL4HqX6ZgSDjeJwCsPCDSSy95Xio8EK5VOAvY
gNe+sdrj3aNNQJkfcZF8ZI1GagYxYvU5pk3eDoLhVexJjJtN436DQ9XvGBjsZ0MUC/ZJyk7qkYgS
rm4q9UpnL2xHNKA6YyLNGBLFOQyWOQd/B4p/H1COg2Q0hzhynhanTsfuLRv+qv7DOlhn5D+Y0DYC
FupY4UOcSXo8lYNHRAlUlMy6vfzw8RfCKFgVUkF2TbTket+4nUdP/LTlV+Wbp76dF+jclO8Gj5FW
YU8tsEr+AORpQRBVYHMFKC1kWGUL1JRy8te2DK50bEJtkD1sM4okNVluUKr+culRKSN48BeCoHmi
/lN5jh3qmutZhb9Snc7eEK0xajf7nB/t2iusD2jSAfwabRWB32H+QeN1XtV9k2xF5f4GUKKSXsQ/
0KqXgVctm/nsZf6gTo0tbql2RkQ/WYkHnFZXAMsjMuAKwSaQ4utY0vWRzvZFuIBCHdxQgwwvVcrO
DqZFGdsIFsAUer9aXzLI4jfyacG6HeTSWIdgu0JweUWrBZU0wSM6pprFum2Zr9VtsFVAO3nx/zi0
gQuacZN+CK9pq2lPwqKt7OIZ2ZaNR9MEUiUk9ce1SNjpBVnCGui2ETfFEJ4DqQdJRRyoyeztL92a
yho3ULbB3K34pRZh7NrXSPD2jomhq+t/Xh7Bhm4YkHyibJHolkcE+vYIc/hlEVQQx3wHbKxGLZkt
DPBNFhmr1kfVhBYy1wih6V0V41XpHJ2oEcfyExq0FQ/1v/7WZ2cHV5QIY0ouaPTFvZjpc7S/kPG1
idwj1N+aRhHZoCbGjWcnfnvXx9gGjiNE5xeiY7t+gHbTapZ0XAwH5ObpD9vZaUlDTqypGA2zlNM0
fM8z0uGx0hfTWv3+0wJvAELO2WdFOGUMXAakmp3lDi731Bwap7Ix3M39BNhCAYXbuAhKyt2WR6Us
5JRBQOR6dSFTUYqo/d6vGrDi+mN27hFqxCZjunxig1Stb1E+36GaQg0K9lPVynJPG9fTbvEuxhCA
Qy2Ej+mvqhb30Aa8ljiT+4OBTyeyjOCY7Rn0ZBkpNpBwI2elQUSxE4n1/PBx5CrpzqRB2puTwB/e
N4vXpVr1Jm/2okSTnwMN84KfAH8D+FewOzMH5eT7CDML7FHd05fXbJX3VkcVKvpmWAR8rEP7j0g9
pMg35X7zklyh1RJE/ahFEGdzzrluThZ0jictI48Lx2bSZtmEzcsh6S7SwOU74t409/h8Ulvm6pEh
oTF0VQNmKBFpTSBFuGYRksTgRDciPYRZWf8tc80n5rWgBqRNCnzMv9sHd7SNdrYBsIUTdaWMvsgF
utYBHZ370C01f7nJAuD93sze6mVlK9T2Sr1lWtYnBjEMDVYDlSdM45E1M7VJVB+HYCt0RzqgMFu+
K2Xq7vKCgoI/mm6i9xO4KDkWzTNuY7Ci2dwzHrusuRg+cpzzLK4UGTYisaicxDKqukoIi/INMXnQ
0aSpGpCAOxq86xVA75xbF6yEBQ+DiScmyOYJ4OVNo6N2WMfaObSusQSU5Wo3t6/1gApEnBkWHEf1
2+xsU8MWpU6J6s80K+GTJsztXcxYdS5dYHNPOFGU09Dv/i8BZjfgvw00VtS0u0WuxVe29Lr/m9jf
ZYjt3lK5NIpsa/H58E0DbHa6g7/Xy0+cPwBqg49foWG5jUo1hhbMorNVuEqTqpm1+n3ujGZCovMD
Dxwr+3/9ar32loulLlNl9qmK/4kbOM1ANXEwgoDtuK6L//dydV7Tk2mez3guidUFuMdk+8fMQAWm
dOnSKtHrVE3s9Fyo0lGzFzrmzRJoYe3yITLFYJ1yjk0QT3V589XjwLKF/HMBN/7WIMxd5d2lzJAR
B2kDktaU901TX43v0V2j8nzBMLgit1MZMlQFueaNC0fEWRhxuWKsacS15kdrVDdJx9MRzfpbEAZE
g6awhNx0BSDuHPoLtfvXkiIYb4+VrOlmAlNQ2zgLkNWsHA7uOizbzPprwRMcMwkYXIY2LLDkqbL7
ulTQO4ZeD6H2+Ic2BaI6KmjV0WaOZH1ntFAWt4jqVqO7j3inIZBDiY5iFqzeelfIMa6GXJ+YU7gD
yArYNLxxMne243DC8q4RlZ17h55Q2kiAOC3nJQRXmDHO5J+GRhuiCe3HRRrqyX0PZarggFVttZXs
uBJfdmx0MBhuF6UsxcO2hiHpXchSd9PJvVng5Ieu11QCxHwYvPtGCRwLGsoUioPBuKpGfbX79LeP
YbAsTKjNzsjtqJl3e90C+ju7MBlNTqt5G/3Bkb+GGH1W+gTCXqSr4auPhOVdHmjnOcLPzTbmDGT4
7cXI7eFjQpI9RLLoWq4m3G8PB5aNcwG803OcdHC8e84Cg77S3MyTbkHycUl1dZbutxq6RVdF7mt5
gEtXF2QiTafCE4TncyZAaqONRPvvGFOk17EnxXvKp86m0MogoFBxZhy7RP3JX83Zz1yW6nKkMvOj
3qgudkS9dpyuspoO6iKy2vxX/gQkxXKIRlp0hGA4YO12l7NRB0XlOBN077fOd/ybdl5RtUiZbI+1
7d38eoLaf11CBv3BHWbdN0wawryyFyaixbv6AZYjDJiQO4A5+q+hqS73G101+LFJazS7vBpeZNl4
ozbRohyuIRe/nEiO/KEj02S8U1R3BQPEZup19Zg17oRRVT8SpKGzucU1dHfM1WUXk0w+OIoHZhPz
0OdIpm+UJ/0l5tsX1pCQf+oFC09mXXIwintYSXj+H5zhpl2vxrviyL32cAe/poBGOIJaOpqAhLCm
PN+LZ7/AL5HzMpBZ9uRwdhxL2BLSq/rHsfZJ0EltXw7j5azV2fDWlHrEOVVZ9OwwXttUkTjiHEBt
hqw9+srP9XH5oMEXe9VPL4DdCE3Z8uUth70PUPAG8lEse4iJJgTcsvkPEimXjSOymZdZeKaBIQv9
4VCfUlKE+gyvgxhJHDbe/ZTZzcVn1Snc8Fe6Kzi2MpqDyBlLcQohNUe0n7JhB0+LUE0ayIeCkKlh
+IjEAEdOMWsfQZ/IliO5xW0rxTGJ+ODpNoTCqzBy0s0X4SFlGTSC9v3WqLsovVIH3P8AZh9gh3fH
IW9v4YYDER9M96gmAIw6xFu1pgwX+76JN5QF2n7mvA6BtlRTSZEkgP15mwKSRCc+Wr7w3KNWkFu7
Uet7pAm3GTmNoYFlpYp5M+IZ7R8MZLPOmKu/oSVPLdCE27rI0pgtPKSbeOGHeFJNam8mxIBFq3qa
9VtgdwgBWYkxV3z12EpyYxnufhQYjUMwe+8+LmsXx3er5x67O2Dg5FKDAUxZZdDm0N2xeSad7y0O
CgQYzWbRJDbdGIcy1dOFne1nr1oh1o7bTsAJuMTwmpizqlG1eQHHWg9U65p7E/5pcDpDkOAl68yc
1is4uBca4cIKXbWegnWQM4++PU18iFWmWRvILXbnmNMs7VPci3zHAy7NPlnF80X/VKh50aQCer56
LjmVnnH84El/S0EY0NzO5NaasRMcg8+DIELlyKhuM+ySjjDTsAQNObSIto339mOMMab16LXLrHXi
dipCfRGQlJOeGaygyeFChQ3oZXxa3dfkKSN8ArtRzPfbvlbCur8je6/OtY9TJdRCsWVRi6diUkNN
T0p3PK4mlQxrpJQlKaqJoKIeIGDl3jOArbtgc0QBpDv/vEEGnDwfPYe3pkOavnxalJSes8596xTN
0+3huiwj0fhObcOQbd47MApyGw4JKb04LpgensYcY5VOWD5m58CdFRL6HhEnHJ3IXyDgw5iiieAr
ZOVJMsT4reME8Diqx9nfZj37DFtyToJMt6SwhfIK70sR0aND4XAjW9wH9ov2Ich/PJpbI4W2KyKc
eny7g+KpyLvnMgJgtj7I+hbE1lY7ufXPyP6DLll+GSn4U6xHqRnpPjFGwLVMToB9BC1MrIpV+VxB
FGyfXUY7iXvCx5L11uj9Oy+zwMJV2IONs86UEpoSRo0atg6kFdCn53M2r65lPzZCKQ73IeRz8TjS
MEaq7r1g0REjQZ7LUsPSPwENZAnLBlnQzQvKLojn1IqHtTQwGM0g6mjbkfbQ7Qxlyh0ZIwORcZJr
qpMQQm+G2TOzBAHRdL/olc3tFM88yzX06QSIRYBxh1dg1p5VeyK8+Y1qDSdY+I8nfbX79sEHOQZo
nAeH0DVEsgOWY/Q0a8l+NSnGOXbsWukhg6YeE2aSZz5xRaypH4cBpYm3uFqXJqeH35b3mg0HE0r7
TXWu0DLdqfmPriTVS8GFk1SJk/70lIn+DcDHyVrXB8gdbouRYDBRWIhETvUjAc3PejqvxNLfuHuE
quG7BgYS66OjyWrllO63A7iFepz0zc47Zq18eKiSWAPXxpXCZzSc8tCMrxfrT9rTHb6v/4elV+ne
+jOJpl1gJ8frHdggvkxuQ6+ZWBobToM/q4BX2g/qhFfIswv0mYMaxGA5h+AXsd962IFXYkcxQUzl
rwTnv1Y7gnnD6xTem3KWREy9Mc4ZQO5ZM+06gKa8xr10zIvDpQkRACWUDI7L8C0oV9HPB9g2dpGS
4ZAhcYMPqUHSfr0V52ZjB8wW5ThLzsrPDLhZ0u7c6k6ffeqoO4pLFEZeGKIVA7X+xAc/XK91vSSC
t8D3lxLUSNcb2Pp15+7ukq/DfYlDvbo1XHBfR/W9XqmDkOnDjiJag+r1c6PzudhZscDOV0Zbf54/
DhtZT1wHGOuhmWE9vYkYyLVvVWBFr3rYZicSlZQWvkFmnVPkpfERLlBuFeKVDpVD7lIttBfC73ys
nDvO0gXAw91nfBegGVlyyFTBhJQcYnqicwbuRKg4L2ChAhabeOvLK2ysv38vQNGmL/ANt3KW4p63
OM6zUBBrAZDTyHqITaYOShLjYVgELjrdwCgFQuwiZ3TrGgm3MJV/3S6wdf9DPrKCp5D+lCYK0t8y
9IkfBSlkfhH4EBQ/ZxTwX5G2za5F6yvGIKa/7DMk9Erz9XMly5Ih7faM4uvTBOTjCKwGcsZOhE45
EUIvhoUnq6WOIqZljTXSQ7kcwuEIqT2N30zxB8Xyb7SVPh8gFBHyTCg3XMGveVTk9wAYzZD49RBb
D9Zwxq8HEEpEVXr+JjUYfgRVk0frVKiUK6Bm41HMBCTcpUESto9AUK1kF9jW9E/vC/z2aucqtph9
emhCJpGminRHN5lP5pbXTWQAr8ghDX4CNyVq6SPkRc9eHU4LqjytocTCNSn5PHkNewKOiS0KZQNF
goi+uX1CPTY6vo++Hyb+J6qAcQQRDoPDiblfzQp+GYh+3jN+6eJJwEnruwvmo+X+9eNuy3TsG8gW
kWITuO/6C5avGCCKsplIB+TvD3vyAdMWQVrf4zWX+V4pKspU76r3GLMkwjkrMfNEasTm4dneaCQM
Hk+iPDWTEaEgJFk4i7rV81iqlMvOMQbciqDv+bwZMCZEnJVMkugzQ/4SvLeTfCcybrNgZ1uifZWx
KDkmCNfgXweCi5F5ndvTEOiLFi2hLNIeUBvG3Ryc95UXP1CyjsKCjDHubWfa0AsRymAc38q5/qPT
s7K1p3nTj1s0Dc3YAOzkIQ60WJFPuoRcqBlY4PbDHN/WJ5p4NI5kVmzmSs4VsdRwI54ifO6N1k1A
fEGL6MJ6p7CLttbnti4hJzOaFCoLjJYVGVlEnl5tO8Rz2km0t8kL5i+GOcrsgT2U9aCC4RrhvvDX
e9DLGow+ieyYi6FMmmbqdlsJayxixzcCJllQ0TSSDFYq+EGplVGmo0Bs/Mz7ZiwFVSvzNW0ChWyv
hrOXijW5biRIYM38N4Gkjb4leiyXQlY3TZBsgeTMZYhnFF+Zu4GfTJ5rFE/MvYURCUyPyexlidjn
n4wgh4vzpxRfqvsl2aSuNcA13mp4kHHbbSdJc4y3rqv9KCReRue4i+EdPJ79xJV3N50Ph68tSN2G
5RFZXlKyolZeKqQPVEPzyeAxJmxD//W8lx4OZO9bOHBgYVKTMgT+D6qVUvauQgYU0nRBwJoMcsQa
6PZzR3Uquxe8IFCpP7orfkQiCj7Y4/665R644Y7FjzRZjQHWyELTGfd9Y6kFh9JOL15O5FAQLx/c
tgXQ7WRhU37ZI9IKpFeEkE44ZVObuQ60Jz35uknu2jDzTP+CPaSroC9BUFrQwO1Tq/CRlpWE8tsW
AYuwkpL1+EPFBvL6YEz569mWazwwdoWZHZG3xoLdbBj2XcIY90ZQHLfnCn/g052TQuJnGWbHiNNh
60zBqHFqMgrK+VRWzuucR/3uCvNzrcfTAROciMTMynQEXBUDb0AWfLacIiQBejSid+4Fb2Lud5Ul
S7/BVU1a9PPVX9OPjwi0rZpyn94G/VOynpQNdzMHrxBmcxfmF4iU5JX4vVeZ/RT/4k5wH7obUbH/
whlECzDOHzK3wfBEk1M/K2RbPuii4eEp3qavOITaZ8hMAjHRkEb4HI9H28djPZC/tbBb+VPpkn/P
f6vUE27L5xOGXksyuJfDL12LCP9gfk/DhZVka1a5+gRymrjRbmRo5VDINt9AdWf5tdcbJLwGqo8c
/LdWN9mWp13/LvIrXdZRP+erS6itFXWCoPtcemr11D1mK7MAMRyuynasj4QeoearziaL3J+35PHv
MxlcLw7BXOciuPLNptfNj2xGluE6OAeTYjTgBzepFbrB/MGI6ljNE/gODe4ZVQX0xIMUZu1FX+KY
3feGVG1Cw8d1AUkMkeGqpAhmPZFBtIzHQYxFy7v1tAKJQAQMc+d2yMjOl06uZ2y5NYxxhLkSLNdy
dbVYgeoo+L7s+I6GBeTtdag8NcmfltW798OujUdOG2OgyF63xKVyzWBFwmjnvpX4CfgxcvgReYUz
BY6kvrWzZmzd0Sfx3phLoknWcGsJauTMY00YE+jyS9N/G97rT1T+f2cJnf8yEuzeuq2riWC/Kwq2
4kHM3ObildtpUIRSwWUqvhyaNaMBtwuO8EHeM0oOF7ksINpdSPNq6VqSJV49a6GcVDB+e5eCGTCk
NRve1eaw5fyl9OBu9DF58mzlnDOC3zMcH2qNufhTteStb4ZvHwTf/BH7yyAXLI1AYoZHFbhXyt/n
4RQ8m+kRVKB6IfHnhzynDexUgov5K4rA5u93M5t26B9Z/yw1aHR/muzxJKu39xWzdFM2+3zjCr/5
J1Y9MjAdOvg4WR6gzx8bWistMl030a2Rzwm0Yk0GnCi6m8V1U7NKR/dEyThD1hllNGi0ijtDfnN9
yNZ+YW7S8U3HqZ2pKhZU4dISW1W/nUO/FELsY+jZMNsnUc9fchx0vL+b7BFCTphXx1Xvf8Sy6PeQ
TL98NIdbMMu0qh7U1KGEwh+/XlK9W3TSVU5lSBmHrnqMjn8uPcARr+iNACTurRs1ehxQsHOdTUtb
MZ87ApNDVfedrPHp28Ilxxs+3AFGSqpLmY2yHNzvAuMIxjdNJzpSLA1yxbSuLLOWK+QTAwUuvynN
hKEHvqoukWmXL5oKzWpE5A6Hunde0mL8I32y/fuP5YkoxHLMKM5jM910AYmnISaQrUuFA9Mws/oF
iHTMFn7yeJP3w8dB9AS/RRjvWGmbzYIbS1YJljkJzzZBKdtQ6gKd1dS6HJU03cHySqNK5Hj+d7XL
ksw3Ia/+wgBLpEptWpMUD0AsltlBbEYzfHJGeDz1aZykdAQ9EpeaTzaD0Qvfy03cgEYqZHlVr6L8
sUU7wFBEc7dGt+pNcz2EBHxEHyhCGkhPT5cXSJwKpCeadXUEcN9hIrdsiHUSmxVKYH8N1z+JugsD
T8W7O0iYq7PLu4n6n6j1/5IYW3yEqA5hKzJrHRcSutYl7JPXYKi0eafRwBWDTKomK8S43Sjocgfv
LjIOn0PvxG8myuxMShm4gw3NFI9UZrZqqMDa2+MVpq4L65aWBl9TbZ8cYudLaAwwI2UD5zAwAY+u
e7xZCF2Qngv/G6ahm7hoeoiG8THSAu+lonSST1JIcJseTKNFXMQfqqyYiLGqZ11uVPvcKf08L+2u
hC2S9l3EmRe6fHIH6FAzJrZLh1y6IV7iLEh6MT9egA5XvdFRITVLlmOEbbaBdjJ1BTrFm7QYTL4w
VXNGBGfgUBJOWSKuvh7VcPrl8m1YtRtrVuR5oEbgVk7pP6X+tx+Y+2DvJKvYvnWaSOlMnyBxAXE4
lm3az/P/bBtmLiz4lJ7Xvv6cDu80QLtrAQnm3GGQCGrPu7GGi0OcqYfZIhJySTSJgIRgdRXF0E1U
8Fvb7oEAiKMBVOsinqW+FzY9UB/Xf7iz8y9aasQlDFcGla/sC87ZjWoUst3pZ5SsquO6wykrS8Pf
Fi0wvHeUFgrz8VUMj1ZMAijWzxfuq5uJQzwVaHJhww1eA7LL+HoxDxZttMgDlyWwhufEd1USv48N
OframyCC/WW2Y0gaWix4kb2As8SyjED4V4ZYwy8oySEiphm3UseG1xee4Zmx7p2QKITfJqzUq5L4
aO2icCfFD4RW3UajWpcmllCZ11c4jaYhrkZ85r9SsHNUMY0sMCQ8PFTEG/G0SMnPag0nXttVhZKx
UuIUck2T0Xq5QJnxywoidPNcl6tSz5iIkgUIMHJvQewEFIw/v9ZqlH6niHyrDuNx7gFGxbDMxMk9
iUAR6u/RUzL7tj6DPgBkgc0MaxrimM5t54xoGxCxZdzD5Rwzc0QSU/iHVrqR8M4CJXceBWGRO7EJ
vR1Rwkij5ORC48AS3uzi8/D3Z6lmM+yA/Ev3W3CkGdw9eAzNHSy6yZmKI7xy/DDoaQISEo19v2O9
I0Sre/e4a07hx4rcIxWittAHRmmWV0+bUqrjOLX96JYiWOoE02CLyfcLr9QkmGiZx0Or0iiDiH9g
IDQXg13C281+otMrfxSAK5r7oT4EAcUBcy0eu4ef2ziaxy8WkJmVP814qVNhXeeoifLrBxJ/WEPE
GQjz4UJ//DfGxLILwUSeCimcO3nIykxz0XpO5yeNvMYpT4C47qf/XASUZDx9DX49DpZhrCODq/BH
eT8RPOpgX6qlWTSWQJ3y7R0J47DhWxjd2Zof39sovrpn171S4uyTdk4IAz56GBZkYaWqEdiCFPIa
YHLJ90VHTDtcoy4YfiS3KZ0filF3ttne4GQT+C4hqfTPst5md+jmYPs+yPnKQALSrdKqCSWqfwQR
YX+1XeQub85lsukkdbcAnXHkS3UkqGaCr97UYdXPhTrHaLHeM4oeTb4sVSb5ZbgReTvZmORnBKBW
zew+62Y63IhgTHjVine4SDhaeJocto38lrcQ7+V+W9u2MkZFD0XrnKgW8aa0tPC/4n2C5YW/fZOE
EALL4HV3NAiaZTFD3MRIzgnW6/IsVYJso18C33lqXZtbnjn8GBjcPcqtjxCPi+XbKUq5mjiJFXXo
0ZhWGPSCUqca3rfJ6GGaiX37LVVQNFMR+j/tYKFJWASlN3cen384dAKtqJA56MgX9F7geaQwMuHx
HU3mIvVJK1F26pL//3fl7yDpYVyBVsbEL6kc8hrRehypSDPaNjnkHG+g1j/81M3DesLh1dystHSG
zfXN3wSh/QaP4jXSQTdbURl99F7rDPCN4zFYG83UItLXPeCTpVaW2t/u3PC7Hoqv71/4CvQruAob
mbvc4LFdRlKznoonldyWso6m7IpW85Dgl6Z4IZ5fU4Qp9xYdzlR+vzBAVdXYC9KZc/+fS4HY+tW6
KHwCg2GW3P0hbnISAdUytXQ5f9EAycr6ZoKvzdCm2JbyGTFbU5dbdAXvK6Wlajem2NFCUz8dgran
y8Q88Eq+HTN5wDU1hWSxUJ2VREdJSgpGpPM4nbqTDE0IN3mcoo+MgGrEOJl0I8ha+1h2pz5+1d7h
Vq9616F+97zpZbAJ+1fC4QHbi2lArhQN3z+2YDyzh68/oAf3gh4zHyNqNIKhwA74OYBFgvjfhf/s
9MppLZXySp2xWRiM4G7LVxR2LH+Dr3NUaR3KcKjBxWOOH3TGAOIkdIqW22ebI2f1ZjGXmU/rCu7b
hrct2FjkFw6gipg3g9Y+4VjLpQf3cniROcc0pSYEsxlkmRqmZAGjYpXzlUqdP0f/lRpyLZVc1TIa
r9sO6rSJBMCjwfPRY9YjEReM56Cj+YVzedHtwixDvoqDlPAVpH0DQd4v/nYP46qhQW4xATB/w+jC
mnQKbfG+8Y+wbPLDvqzfByc7FY3StLEipwotekIJ8isKyVl0sILa6TN+JuY6RYFRNOAwQVU5JIPo
7kBzVVBWrsUZJxyJycdyZ2aibygyLxHOGeqEspf4Jce8fkwW/9cADiBnLkVteQ0zncH9XvUSVr9S
OGYPamcO4FwrKrjtfUJVFti4y3uCQQpghPOKTo7r8PS8vUCzkkaltVegOry68EJvKs8ShD06DiVQ
ryLZUFH6SF0sL41KawVI6bP4Dzjs9T9CHAay9EG//JeqoF3EtiiuIXezPSGNWfhyWsxf4Ym74Oji
Xs9O3aKVq/g5r6gRusH4a1cm8bbuCaaQpTbut0A/lX0C9UjAaQXYbVmUKBBQqYXl7dgQpNRI7vxc
MZnXF4J0wIr2FqX9Md06KpgqH0be8f+ck/L+YxsCSoXRsMbYEu0BXUQDDSLo5eWMvocQ4W6B3pvx
ZvBAQWuKGIA7bupKocGKEum9CvklRLS2GnlQifFFNwd+JsPX6vrKdx21t5i9XeqPPR+TQWpaE/Rp
1jfH04/oflprXQP/PPcsJ4JpfZmObEnrvtCYzYNJfwpfjGJrqcvCvmxQ8iWTbQ4EPMqvnMMzIjdh
97bTaGz0KPuYcN3AmnGKYoSK7/xKkb1OLkbx0zQ74hUGM+lN8Kj/HkvdjMx8MO63X4hQxOYlhsGZ
ro2yeOZMwCFZj742NiH9sR/Z0n89c5v5ZNznKQh/HJFBAlsNJLgOcDc8iifMV9RHR2pNqsbJb+SX
tCAtAxideQlDlBo0He7+1hEHjSvkO8mxU/AlReP4Hu+/+G48Z4QPwhVy/gB6z3+bb1uVNrGJPXbL
KW/YQamfnbGgWOlLrZQd3Dv5DSrjGNadz+R1hI25BXhs4Tu/Hu/UiDlV1zD6KzskXCBQpLdUOuw9
XoeQ7AuRQmfSfYZ1FOFHYBkUvpJpUVmWHpPtCL6ajBke1EzwEElK/dI2htBWbVu6Lxu/NJu6J2Mk
GKewZSORs7B/lyyYUQhjooBi35CylskQoghWet7l5Bx2b5ZPkpGKPkT41bcIlaTUJQWXxSXERA7R
FUnOaL5WDuPOzTqyBZBNaTmPSQdjbC5XH9SNsc6eLzg0kAIwz7c8zZr4/eHhuBlJmtCrP97jEkz4
G1ArayPJBsyGqyriLvM+MMysmU3h9+1WWkIAqCN0ydH6hqSe4eC7oUsQXMH1aWlEjeQ3JGlgR0VP
DLazyRqL0TY9fJ8qrVXahQFCEr4Q+B33/0RAtOpUw1YO1SOwKFgWF6XYEWiv+PEakk3yf9gb5r4z
pdYiJindiAPqR6d5jE8LtlsEtEBpBIvoUTDLumGfftAGAxHzm5olTj6FA6+2QJbrKlBsG173vdMM
RtqIrc0m8tXsigOGOcPV2Zdd+Yb6IppjM2J7iYIMDoPVodTmkSUQYBq7zVGuCxJrsVLrfMcserE8
g/O2EWuOp7h56qGCDmAK1b6FXxd/ohYoP2g5N2SIWgrcddtQCKOZWzYYKmUeAhMLjyAo/iIvqn7r
DmwqhOcLZZg/bx4L8YRI43yABUugZbOpihpWJ3/whBK5x9faSgCzrShwVEImi+JhcrrQUykRfOFX
gF0nVoPT1E6EH8ppPK2MfdQFs3OZ1TiiUHWq5LaiW2JL/tIh/VIWF29bRHCIT5ASj5i/lPO9Ou0r
zePqnNtERdT/TT7YukyC3qIwiymGR8qQy2eQbqyycNUPCgV2xG36sVAjeE/QBgc+ktYgWupA6HA4
BSCS2P5KwEoLwGwUho8sRa1f1y+1rAxBfdOdYwLKpE346rpAz62qi/uBgNWRAC2DzbshzuskGsch
XFRpE5s2SBZz/0j+sc/vrpUdLVq2Q4dAMyH/ly1I6dT3n2660yCSKHdw9RMFNMrQGpPw6eDL1a1S
l5cmOfNn5NXMNAnUsgzmEOtq3CwMbms9de8c/4mpI5K3Y3X4wvXG2kdL2af69xvEcD324pSLzDi7
6ZABeatm+8eKKqOXxndU3ioPGcJl2LfABVq5zLMlPt5oESeQ1IzSYC2487I2lLyhpa8byE19nqLx
XGLe5KvWo+u0s4QUe3A7D63RlQmkUdU/+9Jsqg1QNcrHbaSNsTdnuOKEjolHlIMmO5Dnlzr8Nf1U
H9WI4HlfbL18qiUc2z5LShFw7QpRhqHgu4ORrCYd7BviVdvE6k28Nb3TT3Q4HSnGkewOuQpR9ObP
u+jL6BqJHIOHrdPXnW86KU37lKR4iKk9sGorZABMFA0ri+gnyoonA0M/YtzGneyQ0lXXEGE/mCHJ
3p9e3la5NfOpC+Hye0ijCg/mNJ5ae4Qha/pmDI/xnBJFhszIjNiPrTxTXkJ4+s1Tee7SDXm59IPk
HqBhkIWnTr/32jAVF/AiIERtW6DnlRdlA2/NU0j3g2prYoM1K3ogL7bgvXMbGEd1+k3sNlHp+M/j
WXqjJwpsWdNSGLNTqSsdRMBnOq1+sYKZxoGulYo2crttXuQg24pU6klCC8wcd1w8imNJWdlR0frS
/GH54M/LLIQpYQPB1I4UqEIbEGzFiSioG/aYT4XYF2+LjBp3tDNluLFKBhlsYmjY6nMiuG0YP8gM
al5gNhbo6p6fyejanR4HHaqDNE6EdDB5JCk2xao2z0uhF26v0m7bFu+Wgsmn+Pm0sRUoU0Gc3x7n
/viTNEwlFB1wExGMOjnVxqRRsrXBGDl0PwyQmUPUlVreD1oJ2CHdKczmvKxRqMROy5DgjtASVbt3
so0GSVOVvLpwIqTGzZWTvwqjJUQop6VRZgJjAsArYlS8/JnZ7UOJGi0ebusaldVl++JqupD1xse6
hAczlwrYoPNp5/nD8bewbgRjSnCFSaomn4SdybF0El+Pk9HQ4dLynIj0Z59msSs4qiwSuNbxYB1R
XR/kHSqx0h9JMEpLVKptKJl3L3XZPxj7q4vEap1UOBJ8eutySy930jCs9SCNRyufNZHzoCPTiHvf
YIBJJR5AzeU71f6sZbwrdIc0VYun+d8lLCRKdqaY4dZok+weHw3sO/rsVLq0rhIo0rslN8UfxPKS
PIhkDF8bs8lLaWfxLgW8LYGtI/ywe7NvFuo16PJSbFBJemz2HCsl+ymrrKb8iq/4dMpYK74aseoJ
ofErUHxkxvcQ5E17Ef7KjBH6TjLS7/SfIpCjDRtNumMvOK5D+Bouruu9/2F9XpO7nwdBjeG6z5WM
dustgjiYuUisnk1iX2JQTsRCiC6xSaYBZ1PASrz5dLBdSEj8a1lSJukjAyDAWekQdfCh1U1hpleI
a+qj+HIwv31Zc3bWEIYLs4hbi647hoFC9TqHv6xXJ3ckOIPSdQD4c74lbNAcDSNqMJm3U2AiRkKm
EEQVLWQ7Rmqh0RAueTqHIS7VncWRN311nY/tlUE70iMtFwF79pe8lJQ6dDjT25/2q3n5geV+7WGZ
e3uHGNZ+bl7iOuRpush7MR2nt+loCJN3nKLqEvVzvzwGSms5XG40/DAgqCR8gXmL7OoZ9bmx/CBi
mzo30Zp0oTXuG/h/TP2hSFkCYsF4ns8DaXuPw4pjocA+Gmof+SsBMZaJI5cHtr6AjiiocrEjFB82
M7PRW2YlaIucIKudICx7DDQsJjseRocX/p3CPs6TH/oOcT0O6cI4xyXFjT5n9WDL1QY5MY5rO8ez
78Yu+D6X/NU1wZ7L99I+5tbeTksAMbWaJia9nOYCDn9mMmMpfTrrXTXBdNWYCD100/jAGbtByyWA
hfUEdoo1dCNxo5Oa/DNAtNYGmJcPc10WmdiIW3pVFaihUIgJso4sQrJGV/po5USrVcyqR0lJ3KO5
cwJlNATO2zdUakc9YUYeDtA13m6BjubkZFW+A6NUqwUXtQe8iyYKVha9SDMPigZrUrucDiJC9xcO
+BONAKRX6O8jVPFL4Jb86maItuRyMi9VDJXykFzYYbNZ5yPZ7ej6GYciugckinLtnhI3dDcFMs+E
3/PCYt23B6L8k/1f48Nm4zomwF2aU3fa/MMJ0+9LIrourWzOiXRFFdC3pTGHynBEfg/Opx16qcba
QsJa3pGP5X94jvvxp26XxieQcNZhO2+rfQeJh0HnwuYwKYt6ZpMpDobWhLRyQPenOo3GJ1/Mc2Vc
aExlvZbnm9U8X/yCzhecU3e6Yflmbg7lluOpgacGnGRarUsNCMTUqkUOdSF5z285mvSvRwfWznhQ
jzAnm6nifwuteTsgw3FdU2GrpnbKshbumAaDbYXjYCGQvXNn1dfJFzvQq4KXHL3o9tmiSKZvRbOS
rrTSpkhHNAyj0MmAXM3KndbNFZDpz8pseO3HO/erWFE6BFkYxTWoz2E78yphSEHzy8IfgxUNoPVN
L/cg+85PGAvA4Gc4krvwhonow9VJP6XmBFdCFLlrtprCHedxdfbB8n6uRyqdlAfjpfEztRfcNKcG
VShcBCpO0L9M0QmGVWaGoEcGCnuqajgbiFefu4HqXBWOLSEHs8j0vXNTrSEnuKO02p4J0Y64RxbJ
6F5vgs0727Jn8bHvXXTYWnXnVhPlRirx1ZAlXhFFo/Vsism/7ATmLbBLLEOnW385bvUiC5SnERfL
t6NAe6AiqUz9EVBAOqP086oL0MkleJd160/dLWb9ve2EQXTBdebJinr+S4LqATqlAS8GKjjuhC3W
NPuVcaQ0G19dwH4+arJT/31szWcB/urJ4y872kiNKwdqhu5vVqpHUrpNEeE143KZdv+nU5Kr+g9G
6gnDrQyGnS8oztyU9O3vF+n067sM/16W+kfpXoN9dqz6l3BKoJXjH4BqWiM8pZnSrEFgXgPPCGtz
bt33jq/x4xSPfZ1Jj2m79y4/eB7J/mlBjqfs9HMUvj0+MtBydIr6Obk2pVOvp2mdm7k5rSHbSK2X
rMcVEHcPzedRX/JwVGPJNN7PWk3WcdY83/eTTy/T/er16IbSmCq+SafSV+orhMRlqR2tDxJcQCHm
IdWYZE04aTUCoqHGVe2O5EPMEO3EuR4hq9DFrtJF6KZt44AGhK0J48BFvrOCBvhXohREfeEcln47
wqhPfayTluagEzdRaIictGSeeZFyOOh9OQC+6f0Uko+W0WD8kIjrfUrkJjGgPTr5Icz230nPXPxC
UySfKO693vlu5+6yzbsoHVCcRsH9/gnxF1+q/d1xwDUaycLAGbXNG7FdwoRnISCw5rXwwJvzY7v4
sbb0NjBEGNO+nXZoLyishLMWCSRsVaCtsJrDAinK1xc8cUjtvyocBzh34x/HyvvjxUgCbxjj1NLg
grX9q/2bzX4egPv61/lAjlPhOxaxbVkgBj1JipnUKGpjFnW0hxz9JLFZ6vDDljxQOx5Q48ImfvOA
Cq1OlX6GOVX5xCD5dVBu4xZ+QI8QEsU3i2ZG+EQ1qnnQOOSVqTE8Eil/kmEU6EQBy3+UxA8yN8jZ
coJZWlmfjaAjTonar8ZHm3vroVEhP/MftbpfXoOZy0YmF44WyEkR60wW2caB9B1itKACtlzqnEeV
ifiDnQYgFuuFSeu14+ypKQWLXJqdZHjfC5YIhCYF3dggsr7WTY+Eftkeu2ScduKK0uMqSotwltC/
/LhuZZQrSHFIRt5GZ8oG/1lmG680VQkaSheRi1wnwh87kBUnX2lQoWIaO48DxCoa6+EyGjb07WUH
V3eItZ7f/74LjMrGwJ261vUOtToxqGNK1K0kJdM9NRJjBiJo+1N0lX8itXsj8FxQVTP+bLZ2ug3V
4cY9ysB+gh3orvr6vhN8zBjYSjwNKrdfjEmChYcM8P4lwUY0R/7mo4xldq6kELNgbppopCwydZ6n
8uFPqKZsSdx9OBXDsEbH2XiEN4Qd/abgeoXCZgDkeIcp5v+oGCtSbEYI12XN7CuHSE+Hu9q506En
lCqUkbGvpVFVzRjCVA6h5hvokRzUnqIkEuKvBsPNeksmsgbC5N5TzwdKUGn43MGVCmZ2yfbPdHcb
MsTvyZoKg6FewjUjw217i7FxkdGzacmhViijBzOW2BQF7T0UJJ66wuc5/SmUblBEABWMje0SyPsO
jqwK3jir/AcuV3NSyGC3VK1J+1SevJRRwxmF7AecGDY4uchZA95WuCdTPc+s2CGHVUyeetSs6NI3
80qkKH0wj8LNG9ZxsAonp1Vec69jHO/fPW+9ry5IIi7M/gIti+/ToiDfrVx4TDJEQ7zVUG8iQv1n
+FmlKGzxIGlI72jrYWeIZZBMicoaz+Mr53SXXyrM+1f5Hhn5qCx2kgbpiHY2XQMVolSwBKb4f75C
4i2OCGS5PHoR4k53rfB9ox/su3gUuGIy7gOTsArUUmH6QgTioKNhXXf5nNiU2YjuRlqAF4SLhQVS
UyJc2gaF0rZhsoVyShAB8vdSvXwaWL/g5SlZciOSIa6K/phwgk7flKGSo8+5Xcx/u6KH6kt4OpJi
wX4s/owqCUSxaJOv2urxoUxxmNiatYaH6WkEVik/ngK5Da6u6YDmYy5yXAC8XJeNNDQVa202yHS+
SOj0FW7wEX5MslYRlinu8ibKtelmOEEjeiGtuBBD2zoAl2kC4W52D1Srz2E9V52Np9th67gMqWdk
UyZccgJWBnpkkPYnXgLti7kz2wpU3xBWIZq4iXJo9+KP0FouEwyihJTspDVw+ym8TWEztiboM1+B
H0uPLeqRXbE4LZWr0B9wZQZFW+ZbONZSE2CydasLS7pIWrGvbVAIqb2uWlMDSrFl2kdNiY2wVnjE
K2s9LohNcosNasGCZnAUttrxWO135WfupA3gK/cZGsmV+DEo+AiTgu2ffSPHkaEi2v4X6qM201CE
YACq9RZF/KzhgD19ByvI0MyLl/ES09UVXKd9DbeDKBv7jpw7qCSW5FlJiyPEPTWhjC2fPpupH9Qd
c7/vgxxx2O3+XTLpVv9pL0P7O92I3vgJRTIosgRYmLqCChGlBYYIcY+F/bXYTCrwf3Od4LnN23LU
kD3VMqt+1Pf/mgA3aIfduSmr0H0v3AIg8OtUvM5wFmYXSfq+v+/YSiXm8cS5eOLpknt7Hj7YOPxW
6CwRIOAHDsz+rvTi87xpGRSt0gnIrF9IsO4zizGYteom3X4U/os+B/wp8gkPddFIqE+YNABLntFV
0MJu6VgM7dIZO9GkkntO9QWkHWflRppDid19ovAGF8D4hXUtkkKXHQ7jIV/Kwu+5xwAUvFwvTko/
stiblCW9m/vheP5aok4mwua6Fc8Ya/9gEhq+gd0azEhJJHBrfrQ/zftqthL6q+fnQ5xayemNYFMA
jRFMGfmjp6PLnLjrg5Ke8gES6hcPd9ohtnLd+NNhxUl3cNynHiDRRHhdP4hnsKyUE5qDOqR1ME++
YevnWQE8Ag+6PEI/pOqSBFJVRlns80W6PkcGCAYN4hDfgkflh8lO/lu/IMluWomJoUckmgc5KVAk
ltLmjbNZ5DBhXmP0A61idg+TsJ6iw5YtN1c8n4IYLnIw2MJSPF0N0PS5cw3VOz65WQhQ424ShaUx
9LY0LaPXoHmYaCywgvW83wlorHoQdIA5l7fza9JCknalhMnxWp74N7QO5UFcw4xUnQaHDe2Xr97z
w+NNsUXPGHd8WCz4jG74mhHrNEhq2XRrEnuTMS2WEKNtIiDGhHrebXcsiPI7x5A2j0Qqi0VlwdLa
I0MM44sxyALw0Tf23Ev1A6kvuecv3Vf7XtMLTeJtV3rXD2L+JAbLdq4O+7Ik77Ueq15TMkS9Bw++
rvmOLAlDcITcwshPZAR8Z+OJL4d4VFqyAvXAiTLUD72N5n509TmuSBGuwhRgla8oTNFqLR0XMZaI
3WOVEo9wzdvwA4SiLEj8U/YcUUPRhleutetLqH4jsDaYFdXAvJQqb/qoLUdPNk8hiO1UP70+/Z/P
EmXD/hb8hN2ifGHqAG/hbaxLP/VIWJ1EP7RMQ0ZyMupgei4O9+A8H1MPRY26+qIfmROA07iwoAe7
ncqLWbC2U2WMiTdTy+90fFC09siDMhsdgeheSfQOlhXLgudInoG7ehwHblIYwC14Y5K9yG3PNNOF
+eCpuTvGHqVkJcIh3I1zdhTvYSAWCchjxqr9/l7NMyOLkJrPzrRS5Sg+FKhhO2GPaaG40SZoCsLI
+H8wJaoN1e9gxTz82EBNJBM+nlhGNBKmg82XzHQwNHglUpYDpq8I/Px9FJ4TrJfIFJJVqnEkk6dn
l95Ai4kh4s2D8qChSmIZym+zQI8DwltXOFPtbUvKSeGLffD5Ce8XlZRuilTQsd4J3n5WLal0rGIy
vfrdZBA8PRFy8f9h4nQI/es8GVqsBEyH3Edgdx0/Ayu4qsA6lmHU3yJgK4Kx6HR5XZew9kzy4RS4
qn5TfYN8OXLYODe4oEtwNF3335E94Q00KOnfK4/CHcqKBe/pSczv+pO3VW7a6hqJ55S1FB9nH1/d
Cs8zhrEm1eJCxseylgZL+mnIx57fbgLGAf02AM5wMIXa4q91yJ4bdMYNAV/dupGfuJ7WxF10Yo39
ihWzu8ETdLo2YKkrKDDjWJHovhb0FPSyE17O1rLZfVYZLANdz8FLu2YdhZ9X9ZR7pieXNJeFsdMF
R28kRTP8p09vEcVrFlXbHI8/87liwrgpjWnC3TNXJvyR5hlSJtvjwXZuy4+6xa+w1bFYwnSDBkme
FvIK59spKEYjXxhZADOhMzbfoJQInvLoDBqudbi1tKlgQL+IE2U9pr5qMx86PdnS3q2vSF2UhCij
XspIca0AJosdz+sLYWcOufkRfjNJLALeFDnRc7jp37tMD1PZFm+AwNQZt63BS3TQqUpsR2aHdK8S
DUx46MV/4wfKxcKdP2ai/ShraVFvLhZe7tdL5aZLdEfufwi2MwP4icOBfy3P5tqmnwKfHzW6igSY
ss3c4iBY4Tv0drAkI2xy+CJm3SuZ6cQ+S7bNPMJSPNSkuwu6zKEbsno5MKF0k9AiNsEX5NQrQmyQ
XoNtF1SNA5/84lQOrxKkRDpK6KerttkuJfAYxsijXjgpD9gzrAnb9WnRbpfxNxpe2bzyxa5Po80l
2kqNdUolbnnT19izF1vfGVElqKerd21AjbNMOSP+nBzuEbZQefxjZfHwHB43j2GLY42OmeUYOyJp
Htyqc2zTZVRldQR9XD8JkFEaxCrQmny6iHm9Nw0QJ/oLpXdcuVtN2xjnm0bnPoL6MuLAPfyIWE4z
XHw3yrOe2I20kwQaud4iMWHrXIa6yRAfsHnvDJwInb63Vt4huBr2DLjGsYH95DSnqKWEPXPm4lev
uopIMekJq5qKlXfJgHenKjcj2jEijgiajMy+btrvRgx+Rpq9ew8QFltGhdfFD0EqiBTYIZGOBjvN
ezzQqgQOK3Hp2HroKxDiUKlZ9gJDxGWd+CyiuPWrlI8D2lOebCcOYoFEtK77WJMBGKuWWVvBWJCt
piZTmyHEUQMVTSiWmSeYOJA5e/mnA8d9lnDmFWYQ1/zFdmTrA7nHFdQ4MtitsudnmbD33NZsIOiH
9IqJ6V0ZMMxN8BjDqKPAT76rxo2tATUQr5ejMKf/HcTjgkJadsgi/O9LMWtqHhMIvY9y2Go2GWeY
4TPwP5WIkxSJ6I44v36qne0XMslsr2EqIVtVduos567aVHk3blR8HqhoRoeuGdSYCdc2EFzL1pl6
u5xov9Jux1w8D64wW/8RiZfDHVKmCXXz87UEPAMm7kLJK3RUl/QXhtgy59ot6sxcNrvS4wvyLujd
uZPtk1pAqwQ28Quptac/iASDsGyI5WkW3t/uncM0VEQ3wk2d4smRFSIVvxXZaxzwOIrCINcpt6GS
Uusw4XA3H6Pg793M6u18fJI22BjCJJjqmK9ZdeAdHHkk+CWIBSJf/syuNJcgLTlRTiffln3Aqv7L
h+ANZ96iUS8YSpec/ixj5VCSiJ+0x4bpcGXjBt0Lp2eZa9+unimFP/b8NcruGo5AK6psMOVNLKus
pU3oUJyBF/S+q25S32g1gtQviht4fJ8K37SgAOSXXRxGYLCEFRLqRIUWz1Bh5PdsFxyd4BoTQFXz
ERztkm+fd2pjvkv0bqPn0aultIUCWxj67X+oBcslC0tdfkLgF8chuEqfaMhrbwzPgn3UiHToD3mf
365iOXVoILlHS1gIMtcrix+F0SpiaXfjjFt67hLf0eAQt08bOcxvuONRYYgaHRwiB8xYcyNON5g/
Rfl+PMn1mH4Eo/3wzybaOJt/cqJVF7FU8QamVH+gz/mEjn4Wf1ZLkfM1iOkFQnOR2STQWAI78VBf
QCrYl7LA7giZDwHS/CJbCYg1TLeIBdQbL52mLPG39Yv4dv8/XJFZlS8ry/2w3AkI3Aqej0Nh288I
l/sip0OMqHVhCPovTjlqHCAi5TB3f/wNIwC0MJqHL6YMx/KBXIZ2q5UyPGJLVA96MoeMVPPq7Js0
E9Vh0pu23e60mj/XFcilYi9Kr8UQA3ucDqUdcY4li03ki+HAy2Dz6ukNujTfJC3RfO9D+gZNr7/G
3bXefdipzWNfCcMtay7u7g3x2sj+PIy73C+uaIgV4j8L7frU6II9dQDi9mxIx/BM3nhrP9TuzrVR
PPr6kKy5h7CFz3VtYkYJ+T4wKT92d9p8DWRLjW0o+t+3LCCOZXPp+MKXaFFG507GTB/JpDiNG2Iy
2YtLM8iFneHeu5LFFc93W7Tms8MJ2cJeqgt0ri9ZZrjfaGe2eDjwgfntY6qRVjrVzi7P3qPZ+iQE
uoKlKCTaqZ6CSUlTflFViIrgsiwfZj7v4w6maAmEPDNoj3Y9qSK++awfgxxy+/XkePpSLDO/dZ6V
/JVULtXMiM+HoWG8QYo+iZUv6gjJ0rLEzd3keO08J/5Na2AJlJlVrtwWLa8Ad/RnkvcQkqfSmRq/
Hv3HEYkfI6aJqvJaLrZwukeVIc0Z5PJyW8I0ULscJY1n4agIg9NwmGI/bY27zOr3sKdi2F7W7uPu
mDrPyXsvxx7BCszjJOb75FYN4a9tB3CtQ41uKl7iZOdqFUPaaKCwIBfnX2oSvd7RJ9XHm0ZTA9ym
XJtjmnzg9h8upa1+jxlHZBDf5RL1b3aQA9Zlx2QPoSQFSYsT4z0Jq6JLdMGKRNnEnYG+QVNOnQiG
mBz2qeSzVFJhezQfU/oHHPE7gvFAkStcYNbOJ+3PHDReFOYG1NoLh5qSmK7B2RUup2drkjBJWV+3
UeYMoB2dbp/SqeURGuITDtfL/6CSmmMBcYKd40N9ye3SdH/hbzryvYljuWJCua19w/CzftTWRm2C
6WUH9FFoRgQUaDAiqvfiKg3i8Qa/hTzzQT4OU6LgF4VIqUIHA/v2DpLUYXMLvru2zXnsD9mlk9iZ
8BSHw9SeEZgZIkTOINKsxODS9aEchroYF4438y320lwESzK1tvqRLvRZ3z7FajuAvNTf7tT2YWgW
MQqecHh7X4Lsa8pcrfvjzqEHqK52/mwkVyLJpt+SXODu4+N5AGwzwNmHnKQO1buVUHcduv1c6y3v
vjzxWPQG8gVD5aUsdl/WMF7kGQ2wmXzs1/F/sCeETuBSUP1XSPcUu+R5i7UkDAKDwM2O435igAcu
PpbzqJ9GstrvNTxJVeacCv8+Bcxa4riaSarrttSDeacvWLrVV+pVbc9VeSKs2SgyyPl6v8tAcS8B
Tr3GE5oNb76+ZkVZuPm/xF2I6NP0M6fj3TyRMDS1hwHTPCCkRbkfiWHwZbrR2dW1hlSYe+EwL7P/
CBXvgBz8xJC84xv056WSXlNlACF6jS3dn9rPEIQQwrr3+Uw2vlWk9/1A4t4DbSvHAQa/rMnK+x1H
cnfQujg7RVe26EMD+anDup8Poopl1iCyvk7Zdt+nXFnrsBFQXPwOqeSr9txtA3g/tjrgmdcYB6rX
G7cQzVOQ2bozfYghc1yIVnYOodaOpYGNA9ZmbRJueRKxtgFw5NEgi13nQGUnidOg7LFq5RiQNsKR
OEk0tW6q4l9VpZg0DVKxF8dQSl+EDrtVaF+KjcaXcu+6YgTx25LddrPuibHJjdd3mHZdgOEVp7DJ
zmKF7jljRR3NaBJWc2MW+iBr2rFq7AcW9Y42WUnq+e1bIKVkpgv+Hg/BNeuRa0u218ObmWtZav5y
G952xLNvKg9TCie8Nw3abIJ2O/vf1VbJRoVmD0rHj2UiM5CN/4nRdWnWGAnU2k1BDv9ugknM6W8a
MOOGC5H96ngYxWBhPlCOO6KImBYcfE8nzO5yJr1wONaXVJJGkOuqF+HFrJeNkFXj1yJRyzbjyLTo
blXZ3y5LciDpq8jkqJx2Wy0uv2lty9+JKBZHZfU32BQopxTwwIYjlXGYRSLM6CB80Q8Srt1OF4Mo
pYyaZQweljk5wUf87tYYzDnnN41G84rq2hzSrHzhyLRuFBQpoIW8ipX2ZS3ZHaPdNn6P7GVTwxWN
ItMQi6eJ/Y5berjHlJUqJmueZW5Q2H8erMYR40HNM1dN/cobNjKALeAfglS55WZ/1MhFG21s2b90
KJWnq/BT1bKOuhWvzNqDrTx5s179+8F/T9QsOJnn5mrb1ZwPbtfLeXIgseWALH3ZpuMYhM6mOf1A
bq4YesO1L6C4CTMg+lO32ydDm82/0czJHqWtjgJa9QHczFY1kMdT3axmmXhvYJSHwir9sGVivfWr
u16i521s5WHyHsliJVHGXpF4t0cZzMPS0YsPuVV2CfwwFyDsHdLKBXAXOPmAGsQdkU0aZfhTJ+kF
cQFSommp2QaWsYYG6cGf4SAzn+OJsZUC+3R+0ILxlrl4AQ/G9W8zosmu4vG/SHhVIyRoq1CiiSp6
9ugfFwOBc1Bnd/3NwnjasZIKB6g+qxLKwdOonSYar/nRBhHWcjeiKoafachH9qrDBMSa5MbKGTE3
7PPc+N8JV7xP3C+lUj9lOageaZ3TF568m02jHZdGwlxQFwMASVwJnijhV9Cn9qXhNMbHtl8nA94J
nlWs7dn6gVwAACvLPQisdE6PKsdQMtIGbje/I2NIQA/mA6CC7DdDWCQ2+4GDy450UdROC+OrpwSW
yH4KwwxlVGud1xm+DMJYhjWxCREu3tL1ZilTDdlhCOL4V7Y7X+u52UcytmC3HcN3+rNSjlE49KDc
AeCqYu/W88lue190BOX3jdACDo28OeXH7dhZugkIYp6ld+oWOwO8ddIIn8tnC9M1QnR6w9br8IlP
4iDCotvgVsR3ddmvVGwKS1Th7+nwDv9xjDln3ugPe4aHw+Bzc9HcEUwampMPoYjzf6YlTDt80T2u
v19cTdFCxzlmuZMGC0GRxL4ww9QLbTd/qFaFSwdnU4k37cV4RRAHv3prb4yVUSSjgMDgbBZdO8to
NsQ7ArW/haO3Q3oc2MY3LiOMnB8s0hl0nvWdX72kQFn4EFrfa9+sbIw8vLGj3s2f5hqp3U5jrpji
xl6SLU/K39x7zperj/IwvnfihIvnE2A8/dE9bnEAINcPvRNDC63ReuPo6YlZV9WxViWRl/VZA6Pp
0NM7Li/fpyOy5X2x3deSBaj+ILg9t6DrQwn/r5KNJsNRc+SJffDRpEpUu8YyMWFfpEvez6GG6ojx
rM2OBq7JSrPpJcCQdBM15iCCkfQqOA+27IpUOsu3zEVhbq0mmHRJa3HbWLWj8/GNe/VHAMLO0gTG
FhO7cqJr/jH6alwyaxz9Z76KKxZK/oLZo1NDqFkE1/+el9BFix3tXY4FPlNCl6n9MQ4pvYmueqVn
ECyngwfpzmou9IlPSd4zHowFqzh3nJhMXTHKZSXSYEHMkm0yvEiHRiWnPAZI9Mk/IAEMJ6oXgwwd
DecK07Mn9AKtYFFJ8F0lccdvdpbWhcpkgffpI8A5NzdSpOzkPPyQEV/5Bb68fuE+UNKvRTsXwtYe
3JeD4swgUXnGI61jrNumOKgcZ8aDMlqmeChFdJ1oOrrN4SnEdLiCoo2Wo+Mohz6RLOhsAsssrtUd
OdtvWYs2Sr6/QCgwpayHE2eX/z42tENfuqp7541LHZol3BqNcxllv2w7w+avyer6dLxEAjgbJGKC
R7quwEAv9IaylkURC65iyDsSL2fndpZrgQBl82D1e0/N97pNAXDJGCH3fUpKsDI46IyxlRbqYTua
y8T+eqGkm6cMBcblMM0b6WzKpmOOzObibQqBU02UXNOpIZxUgcN759sOo0fGa/R5lLDgmwmDTm7I
BUHOgjlRB4sN+HCwLmSiVDipe1kBkSKTHrU9oighGd0ZXWD84srfUE6l93Wj95NP9gtOznH35I8t
6Dd5nwWoVld6t7vqRZEIy/FF5f7YNq9g0+BKBGMRxrQaQr53pSpAUXOffu6TAAOie6UXeqSg3U8i
FvULtjeL2dTE/jKfHw18y+SFUu8hTpgaeYctVrKYUM8Z1avvm0OjKVt0ypzbTK15UmXHhbMz6beb
00HBzf4p9ERYccHBwSF1V9BX7K76xHlKOCGAzVc5XFk8XWy8rxmSsvGAU0Rboj6TCg32g52UncS7
F6Rf7fdKb+dQk8cmho6IdgTpHwHlzSvsa3RQNvcz35GVL8piHXcj1Wnc0ACzRnC+tRC2wpXACuu/
XRy8tQ5mRgIvgji5NJjT7KBO+jcYkbaj4UjrdqW3TPtfkBhdyoplNSNtm9pzr/PBpAA4cZS4O/nC
Q/OrlbCweOMPoj3GVdG/DzL4O18z5pzRHnS2kpPqF5Jk9kjTvmdJY3NL4q7Mq4F8L2Y1cV/PqQf4
ERTwAS5yLYUB86gf9saWU+PFXbE0ItYxr/vGHXYli5g83pw0AjUMFys5DePNZ6cgmTYaI+Kc45p3
SpJkMi5oAFDGxyF9QE2elNg0OxkFi4gwzYpiS0obkBMdwhu6stEMXqFeVU+Uh8ToytBhnAowGjiZ
OAqs2BAWpxzGTlShrhFF28hxomwLyTsp+In+vtsn/kS9SjHzeWeRbV0Vm9lGz3cDTrcCZN/ur/qK
7fme1+2wD86F+VFJJG4X5bXYYHA9+2bvcse/UJ0G/eX14yDVi4C0MrfQhJ+iDoG/P0YjhFnucveW
6sjTTVigtzoEq+ZIiuRagoWTpuoTypvAq5iijT2hKyutyApBEi+YE5Du6xGEnXvlABu08IFUI+2S
O9LOXmUM/405KAk64o5OIENljt6/rX9TWPgJSYP996o3168mwGcy0/xYlAHDoNBDNgXdyaZBF/QQ
jJBSaQoZS+isr0RCLqzP01AGpfLOyZ1F3z7V/+fDeD1W3YLoLb6XcJBaaulo/qN17mlewGbPxTK1
tmS5AebHHQIdBCuTz1C7o/gdi7LEolyddWmngDDThxfCC+RAVv0tNZU0taaSYjCF5Bl5vBJeLRq6
0wYzg9jFixKXQe1pxcV8ti8pJg/H8vyrT527V4FSaTRjbRmoAhV6YIdBBnW+JuHxGPZxdyv/kNyA
clQ2b1BipQePMPq+TuqXFNmN8ofk8Jr4Sn46CLMJhOO+OuXPkxyB9jwleM8m8Y9mTcGSYYWeAQWG
v3fnViPGi3hGWcL1MdfwvFBvvELo94FRCX0VsRGHHg16Ix8qUFpclzqCeKCt9yzJ0kJASZBN4kPv
ri/o/Rg0yDpsTf6lIKbZ2cK4VrN39AXCYH4IJXMFl96IOPua0CUvqhSmVm6E0k1kFIU52AYLmkn3
hf//NhBCQAuTZBM81ryR89V1cBwi6K+qua8y9NB1IEjFpZRPUeUYjU+JsRixR3PknJaxJwg5MFeT
IMkN+byrTG5DACOjh67AhhMq9uEeDMMpVvA7ey24j+1e+vQFNDehLndFJDn1hXCvNhJlGqMxIbbk
zluk+M1Y/dqhhEL/V3I8rIBPpsFM/5c1UDP/MeXuetn2Z0nZfLplQRIKOz2EcJiEEuqbqYYQ/BjZ
SI5lYlmPDz/zg/JVnp2xlf4/dJDGbAyGJAk5+NGQK+EgjE3Hj743asyK16dmrNA6tNXXTBjIDmGG
QAEKxkGDjoDAwcDEESUGhBnRpitSbMcb6yTr5JP5VGl711k3Z8EMRwKbOK0+SBiuEStIBmDQU67y
VNJ8rthspT51hEXBPXOerViVJlm/Tcqu5tdsXhIpBr3KQmWb6ylV2v2+7xNvvNCFyCeHCDx+PWhY
WcexpIQFY41g5Vs81LwvPU99EK8QlChpGtwhQq7f2oMX+Z8alJTFqR8HiPTLuLkd/A6AqFPqMeGS
Tt2AAutY5tSK/gsoEkNFoKGe6u3mGIL5MirwyRwPSN8Ffr0mXhs2sqoq+yeiF9YCr8++p9XDjK+L
iNSZ40dWB6y4XOgZeS/wgaVWOyA/nq49oxv3ouAj8qEPjbZO5eJSobZowJwLSUvcky+d4NPrcH1Y
4Al4SAQ5Ly9T8Ne33muIg9leJ5Y9WtC+c7zn+J78d/oVry3zUanRIV8V2MCqcpuWBA6lL/vAw8cn
9T1Z+uVzRHheqgRHE/gaaK/9pvKKO7HnvPcjcrT1iQqcBV/4hxMB0ivdqtrLYUdilVSBdZoNMh/d
aIeh+Sh9f4dvqmrfA17BOLugiaoGWwVAlX3/BSQ37JIdVusCPEN6pHi6t4NOU1BsQFcR5AMZIvbS
fcxtBoxdk+88V8+M92E74XkGCmXZi9FXwj19SSkiJahLPy6E1WTGnSlko1Ay34xhRspxxQ4tebU8
lmjPFxbIBsvHSlP4cQ5cAL2Akrwmjw1TIKjG4q5vMZVTtbVdWsCQ9kVbpbLWBO9r97F01b6SIo8O
fzU5+xWi9djG7dE7vYxHLwHZijvqTmtCbXhWUuMRVL3zsJFE58LkKV8cHBU+ETYZB01VBbSHyUDK
oUCoLK8W/yf+58UPhAUMqTOxrXIiruZeK6po45s0BTH/X66uUEDtqB949PZy1YvKx+H7QmWTRehb
dtL/Z2BYKa2mGH3ci59ev98hFOFoO0fmiz7QDNWjxp0safYK3yBB0AB0qKl/eEaPZLO58JSMlNf4
MN6k/tnsWZ5Kqv1vPX7m8lO5cJJnqmXsF8FGt0pKRmbIBgd18yuQG/GH7txqrVGIzVFxVbJM4wN4
0NPI0O/vvfFfP06yhVJTKHMAFv0UV+3B6+Q8mktLA8n/NDt6XZMGvuZV3LD18978AGgzFl4PTYOl
VQDTt6FZpc/QZvlMhOW6yqxke14KcOcywKvTcOmXQKeKS1UdY12TlGNFKMvNPE/XD8laq9nulQF3
lxjv66k8mCK8S5wvwtor5/JfhW+1nRmur1xvSS+YeT84lO1OfkyzeQ41fIZcu83zBZ5BV7zWQCW0
WQF87t9AWCiFELZc6QVuDEVZujbZ9g9rOUGwsCavfE2JDYjENj63AlHd6tPdd6HDVv+WjK/MuroW
F4oNCv1Qiz9WwD9O0SRbEG3BV+WlMAdz0zC1bepgmcrSj7xlY8H/yuOSuNPQzsUWd2+r499xhNPi
IsMdvznMhUtaHVdmt8T6r706Kmhct/CJTxwyiMa9GeqBiWFqtL92jmT1qQZNdpfqo/llR3IokTH7
1abjdYL+2v93jaUWGkCc6NMZm6U1AuDMT2+zCppY49FNFxcGEJmI4WY0BvV7TjCz21aHunzQ5w3U
GuLNWlINy8Ek3NzeYi7BqWadNi3LYPEHf6MobLdm/vciLGQDUotHDxXT+LtnABsO6wRoi2w4+h/q
Uwo3HGQx0GxnfGENlpLqcaVLSKrEnsG56LngyOcFsRuOtHLksjE9a8CtJnaJrXaJyUDtXOhrkv/c
toRkV7xu5mXHdnqKgNVaqADvPtjgQmUKJEecLb+SmSgb1cuEVK1CZIYxxjIMT3SY+QDg3487xWyK
33MJ+DVxbT1ib2exBpAGnji3ypQ2ZPwrGXfI1UNddFPPe5FXnVMPnBI323FZq6FuMeED7EUmIROw
zFhr+enWqhf+SRR29EU6LHl9RwIMVlUpc8EIe8tpi5K6FJMP/47bgymxOGV5s05/6XMZFVeTrthe
j4uqT9PFg6TGAc2uGr8Cn1vLS0d7JcWAQggY6n90/hUhggMlcWJ5AdGNdbg4o4mxdm4/kw+TAfu8
qg/RH1SZrr0Ip/paswtqUZ+ygefWFN3jKdHPZOe/oZkOXW0EJGaZC8lWsUbWNH4RJ4OiJL+d2ieX
Kt7saF/ankpHy+FoYCQC4fqforGSeoQDe0PYf0id+TxrqTsD2+ORcsN3yzDDEwR2UEWWuutmx8RW
Ix4kjA3gpYMJenJagD2zv/fEqcjzZqqKV5IPa8IJhVz9TG0R941vCWygL67DtoaG3zeUvU+qb2R1
rTOthdySDQWPRcO7WZt4Z2kPDfArKWHsm69U0oaL2KG/j+S8SfiCTzxLX0t37Ol9GXzkimVoE4k6
maTFSk9fDJbOC8rs+NY1UHi/XIDpWFvcnRDimHS4QqHO4sDhOllWrkv3nVeVIygWMI/YTOmtKArC
7RsJC/Ljq/QwUQcbpm9QahVG9rnXew+ITLySAjkAb1YZPYpIEosOk6IIK3dYlWyDk/grSw3k+OpK
DNQzISzmfz2MOa2zieADpYHn42zh23xwLxkkUkI8tPbYky0/2h3YBuKj5dN0AGIgPQUxOUWtAI3S
gp5VCXls4/H/TzWYtS0ezPZUeO7kBDCjjxyanbHPvATesXJ2HA4yYA8xTN/1pDvcXyJuszPTtIwK
/9HKsQxmKegwKsLWyvOnHySALdkW0SjTWQEL+wkfZMlV1AXioWA5Tle0ciM0x5VzEKE1m+Kqb9eR
1g5ZyhKFvRS4dIH+9aNRgzFSuIgubb9M4/XAwIFSnt7/U7aRvWSc2oSKIoZcsH2VcoNl54sMsAed
JnDALxdTWpuyi8F9Bzp4FJ4O0SRnjlxk0jnJQinAJcFguLzTdPlMBkQm1SDnaa6LEdJZE/bkQR+X
ir56tatfUS/4P+b++ox2djnxmw51U22LHM3cKZD1r0VbNHySRgirQzWx/3aAimOH6yt91Fn7781N
LrRgUrZAB+NudR3QhC4qReJQtOktQGDj0Jwep5Og/Pq0pYJGJ8d+uOOhdzTFHOYJ0CN03CxAM61K
FwRd/qByU1q9kWDBjt4D31GBxUvvqcWskWCctlNYbnU0cIwXuwB3cZNuxQROTt9SddlesMhY6oU1
6Dggv88r2o9SH0+eh1cT53KURwOdS6BOkRsOsdwTXDtwxu8wAt3lWTrjArB1viLuN53fW9pO8CXu
iB5bqNZ/PnDCz3VN/sQWH+doYDEIVw7ke0K3hXzUBhZhg1FzmF0hlkRPf2/1OYM2xs4qN/MUoC2j
b6CqACbSlLw7Lv+OTj22A89fVcYFVB5qjeSdwKii3bzgbQmihi+kMfjGrq3BIJTYoJ5KOxU9yynu
ba4H5ScWNsZnsL7KX64pW/iAdRqGNtfgzLDf0zRuMzdSad3a2SP4hBlyYt6ga6yKdnb8naTSK93U
FJ3XvSqs4Ym4TcxgMyQLJoWKpbh6XJAucFfJhzeAliPvZ11roIecnQZXXBEnxwoe9ol1UEESZ5+U
iqNGd+3NLzRJ64HByDy/9u98/fVMFZuDtEMgYuY9rKPi7rG145+hGmOyA/kwQCO6FWFnDLdlKe+f
rchDR0INHWGPuKHuL8CI+qTsvl78ztfCRM/k6+gFk69TdFDyhD/IK4MwL0ftdGruWHvtAjPwvTeP
STgAQppbE7ZuHyEE62QJ0QrXyBaZJiU5z02i5HzHVE5a7Y6RedRoqJu7iw0+Wk6zvK/2UYtDQems
NHEfpB88cbO89OhvdVmtBwBmUfqHslkTJELLYGSvelv3yy90obgdDqwUkn4Psk0P55fD7aFbfkJt
zvkVwHxp6eeCf7U1BUlfNfZoIKshiHSfJz2/ScWrFdUmSMqZLprY57rRzBSJT5EYFUFud3LkKrXl
N1EgOa4arpL/I5/Yu3KOlAwZh9zVL/GVI3xzvL9364tkqlxDZWicV22eo2r12G3ejhaQ/ue7f0Yo
UtOUKmkYf0Bffyj5dlI3V6mndVU8xzNdF08gP8At8WtKv0mciZwOvshp8OMNIjTRMzTmzw3NaLbt
N2/tSdb8ClE168UkXVWCev8d1smCx84hWANSznJ33ZvZaQLsCpbDp1+wFlRfir+TeDp8eBnreFLk
cFwqpA3aLyjaIpzjvz+K0uRSxisuoOAj2jvZT3r6gHjSO3c+/jHghVlAHc54cvxR0oSMyQO2qobC
SPrp3HHqKaUjaCNSbkLvRLR+3AHZKuZO7HIX3kyNketgoS6IGFHRkNnscoUJtDeGMYCyWqUemlYh
o81gWPDF79/cWNP1cat26pspaF/ngQlmxwYdz5O1rh1UBY9+ioQzb6Z9tbVx25V8gS3wBanqRZpa
ozZOSj3cXn+eDs43Sxr3LXI9YWP3BqJYlAPZGDCAXR5eYGK6j+BU4QohkIhWtO6fz+M6gLgGSjZC
loTrRnROMmm93KBEnha7bvSARn0oU7Y/uHf2a9FkJRwdwTr4sXANpbeWzuch8RSoAoE5Ar4ltR/I
LOLBFgW52vkzGtuNWbNN0wLTTT+Licg4N/CMObAxl2SYAAjzpiI/Qa3pv4f4ZQ+IaKjvQ30UtW/p
hyw0dkz4OW01+J527pJPQT1lXvMqzfhEL1lyevxxWK+F5Axr8UqEGAOPJYKGxPQlhPgsFW5Fn6cX
O+zATfWQd+ZyG0WCmkZzn3jGlG7B2Q5bS300n+wkHHdinUfyG4UbvqfwbAUQx631oMbO6CIz3exL
CmTh1ynFIM16GsVvdaUq1YeityZYVPqN9F//eZgx2tRFwlFMMMyHBYYvVpBcZ+zxM32U0fja5axz
p1/IEVl3iMwrTb5DPt68NFQqy4asQFt5UnOlV8tquc7YyadKy/LM0MqqNzEjbEqlcjqipYiOBvxJ
OgA3h+sPtvluerTy0sjyttugfpzoAv3UruhI9eGcTp2aRZ1yRVPXORauebjrjTssghjQHS8trDa6
dnC0Kc0QuMAb0lsjpt6B/Jhc+JUn+T2bXljLMM80ZDHWykU2yIBgwQYQyhI3l9QN5IieOz7rN3We
TNIQJ6VKhC7Z/8SHaVAYYVKLl0U2+ugBB+p5QxT6I7m4YRQyAlwzU7FewejL7nPIGYOG7W+HdoZx
cZTIQmeUzzBjxKeS7A1lePpQKbp9ynjnWPucWBLjhrKV+6b645T7uWTZ6bh00UOJP6r7JAWBG92p
kKul7hyh69Ccugea0Vo6l2Sz/pA+86R2EPHSAQkD5pCvHPN7Ft0giSE/Su1eIPYbKuZHXXRCu7vO
bg0O0UXZOQ3/pqjoXJ7RzTXffbsg58BcUADKHhIvZtfcBtzDfYeIfEBAybgzw558XR3Qj/fUUFQJ
Yv4H9Gv1C+gbiTFIGEnyG6ol8IcN7CtbhEOdAviVCepe5f/yT3Wh2zcomhanA+xMQ/5AW38SroPE
QVugWWo78BAzmgfpsYCqzIwiOcVWFyVgV2rLhFbX7NyxwaDdSSSU2xHTI3iQuORvUNVL6glToXoW
12ENHCOQbviHWUQ2iR9k+Pfqz3IVLGHlQpPLxeY8xzO5NA8fk8fP4En8Ubi9MPTJM3LsYN5cRLSH
iH/qYuipmfLXI7NTeri53w0TUqxqCSkGMGrcpg385YFq1+0VDyO4FeJsjPPDJU/PZm0OKzlYK3CY
vrEhVGNanCElHcVW3LQED9KxR2oVLc8PD8V67mJ7PkSHhYYOSuYtMRfCUYUWcL6scboumH3c7gyT
yno07LYIPhM/+kQI8A9CYl3vubskKSJ1eNekcZ74e+TdvF1JtxJuKvA85nYNxqSw1GjXlUFPhjQ3
0hn2XHFGUgeN1vvjBEjOaB+3cuJMTcESEOZ8lf0sj9pYjdE2S/WaZtJcattHFyJ795y7Zw4izi3b
GAVQa3+NtvOnbICuawJE2/5rCJad02eJzRlfayGt4yQlpoNxyJCDYCoEmXVHxjKahvVvt/ZwFXuD
re2/OQ4NV6SCdGrxaPWui+79SpTKzjkn0y0vX0eGaUOBV5jvCeVNL0RMjtwD6ElrC+7nFvaJGbYq
iDGeHNaWgH3V4OwXpbFfkULKFgYiowCNGtrT5OWIvmgH/vaGtL2f+8T2VI5pL2A92H8CJhk/TZLV
GzYAiD/K0jRvbgK+RU1QGk72ZVRFj7qStTMgyr+3l5w1aXRIm3a3blAEWJS1aHdO99IfNuqGBsN9
vZj4oNtudX21FlRmDKqahC+aH3QgEWTGpyrAOLwA1Jz06NOgl2TXiCK1FFfvzPcQlVgk51ICXDg9
hn22IxOOkNzmdTeJrD+9epTDL8fd985nqKO2SH8ITkvZ5yiDCO4qJm+WeExXQRZmm5Ex7OsA4Rqb
3G+Us9F6q86DeU99XTaT92FfjRPzb+3uoqRvayu7TwSmQndy3SAwQWTPc7o0AyMeaKogimvavf5S
GUjCLoRwHHqj4qjeVdMfE5PcDKnVobNRD9bRvx7+58JE34r9niZ1hNrUSBrUKefxhPTUaS1KLvLb
nO79WMeNz5YS3cj1J7AOCBJCwQVlEj1hhVn15iMC/9P1JP5UYjgAASYwao6jaQjo6/l+SGRa1USL
guLJq1in72nJjH6eJBlUTLMWG8AZiSQNjkxEGQJNJTyxObKeBPue/2fof/we4q6zIHjLWeaDC9xh
0Bzu71vmkDgnfxIG1xBlibmnyn9EHgtzo7sTRMEAz0bspB5vCz5hVuda+68gd3f2Rs/AU2K2BL+c
mabE8YZ7vFvjd5DKpmoLGXGNJ8HZin/BvQV3douJOQ1UbqOXyLNEwDjdWwc296Mv6I6QYgCdkJGm
ChfJ6/vqyflROc/tFoz1OgHMm7WNYKl4Q734+4r+Q682o5e1nzIbsOBLqK38Zn52iZP0CC+7J67M
xrBIImijyjzQKN1JtPkJLAkB8D1Lto5jRnlD10pf+49ErDoNEbCo4mxiAFtH0xCBhgp1N8ON38jW
P8c9NabzR95iSiADHesRWpEWttXdsk1Teb4KuCKpnRVu5jqMadOYBO1fhXCCv9y65SSlrrTRCslW
paDimgHxsWP+402j6G9OAOcevEHW0bgdwveQ+vlwSpBshg7EqszHBevNJkZ2wFAffUDt2QLsc06e
jJQXWMTOC+FfUm+S36qK2S2FM7+2zGNSTGYhfhGxnkiQRKI4gFZ1s1p04irdrLGO3IJyND2LYuZg
6cvz+CYcyzo1KPhZRf5m9tapQKPP0FkHA7KYhBle4W+PW6/NbYHmqa3vISGKNe2rRD2167M1RRYU
Pe02QyLlknfpj7jDQQhykj2uUy13RxnYObY3o0k61mcZj8j8cINiC+Rr99LR4joQjmZFxwDVIfrb
R8DwDUTIhO8Jqjzl9GmVnpNODCJxmOFphgMn5yho//hCW2fIgNq/mO3h9bYjqdybJvU+VrONjy1Q
RGVoQGzPM7EYGuSTb/Ck4BQhapjZIfYgrvvN2CiMbAZNj9uJ2/774gjKYKwxxlhLPMRAQVwNtRe0
QQRKvJM4EAG2md+/vcHZb8ip2TRBD/fpWpwFYmRl8dj6rXLFWcC5au6XJk6vI72A9PSut/hClz82
L0CzZQVUmzAilLMmibWgaLxUAi+hq8/xi/oT3xdFBbHSMftwoVxQIIR5E160gIUdrn/gBo4zqVTA
DA1+xVN/91grriXZd3hloUjsFLGiOiDiw8Lv5h5NB3SvcTiY2lFg38//1Vko5+kvtzSYadwXj6JM
K07wLmmp6AoVMO6CE8PAOd53CMPYRdXOyMjF+BDthkRtc2dzNmZTch0nGKIkFz3h4oHWA7N4lDlQ
UakExZ9rvy22sRzBHv/eY58t1vC/6LUnEY6rDNbHbJxj00Ya8Gf/Tx8IZXfvVDPco+dkYgE76Pf+
VfDuNb5PsKREfxHaA7hKCNGe61HLHaZ3TJI+jWSQ1pFAC46A8u8iQOCz+ICZ38E3No5kOw/6PRfW
T2GccC45rq1vGVwb/bsdPGbMWAYPWMBiVfTljR+k7p7xaERibJ/hZxIfJeZZWwR7tdC+IsMEe7V0
8QEEX24PyYxNE/qD0kG283yzfaZoNwib1ESPv40v1Aj6cCzYSofF2XekUYC3gRQk1ncnQeCa7i1S
PL2kYkKyJ8Eo5CggFg65GunVQ8FczwqjQKgUrAL/vDYZBq91Je3U68DOAPZZYzRqEoHGVlgmzzJm
lMPTXPN8Hff7iSfbcArkTHHLDK080vtpwOQuiwGaalgQz7+jWYoWShYbeXcUza3vMxWXK8dTpkRN
QxL7pES3bw/uYasoItXco4lOvd3VsS+XId4KE3J0Jb6cPjvMLD8Lo7ZR0hxg0dYqu1e6koL5E351
15nBSxWPgBQXbM8250+8npGWHnE8VgDUMPJ42O5YIxO7eOVEF+9XEv2CjMbIVTE5igavN16WbtqO
SFWy0jOt93OoJsR3bUXff9FvfUjWQ+fpHeI1DLgFuPrn4G5MhWg0MDvndcAbQSNpwhPwvfgvZT4h
T+u8dtDP9kDvmRJwOJTkPycPvloPCvdAzVnXyXsZQHKmigEGm+bvKiCxcb8/c2HzBVBZEy7x3FYO
3hLDDku2GAHQ5Uqq2lKrKEdqtkEFP2XA8THq8C+2/r2m38LhC9nxp1+buwkdB9plefKKEhXMjgOs
30CBEmCed3ZGhacRCtVzlViwKvqE16m/5zdApjxs6WiFkYUt8l0fkVlD3mVN/MgVffettdxaTTKP
4hlwms6dA6KBGze9VOajWhyjkraBxUIEpzB0QzEHL9su/NgQ2yMMbAFH0RCT8V1yFQdf+IUmkgef
GGCA+7NI8fcSgqQ/tMrGdwH7fD11wOXdtQgfWPLv/4OjwNw/jmG+r8v55Ch3xp1fzLJ1HoHdkfrA
/qcFB9hfi7mkgzEz2pHhBB6D8nNV5SZNG5yURSXLfK7lqEU+PzqL00m5ajQ9l9Bb3L+XojI/E4cL
A0Sd12lH0vKFFb5aKR102gCUlIKvXIp069ujoatJhB+wzUKWvShSSQuaVBmD28whXQWB/wyxgRI2
0qUVGVco9N6xnp1+NBLrz0Ytxep0cZJ1atMyFEI7DyDzIaqnLsZPsbHjUfqAFZA9N6lYM7Myb6DS
rdJJa5avJ1T1O/8NeQlE1DNft5JBmrgOwNgB6fBG7qDcJmB71aA+2bgVlfms0CdHgu+AxKUyDrcV
hYYLQIR11luKLjzksKV+dYVt5enCNKV7BQ59acCu1jWJEUz4D4+4hJvWuapKu3E9K7AOkqf6k252
nR7nn5ek2PSxkWCTXy3ikYj5J0XDIJ3wtmnl/f4flKtB4WYcv3gdjrGlPSBNfQM5XsC0HKzlyZsQ
4hLpj+sqBaFYzBfcKF731+E4gu23LaEhUyQNfAgvgy2whpu3IdsHJFJXp/NXmoAkB05y9qP+8GEF
3OSZabmsypvPC/UgnaHsOQ1QBNkLqql2vLThQrkVeYOmUR0gsHOYqhvhUJuK8YUXCmoL4BnKv2Yz
StRMQjJ0/M1R4LDmdxNRAy7vHt0PLbz6VEJdJc0vpq/qYnOsywnKRc2g1FBuk+bhV5v/jRGUfYeX
Mj1llwRfxawHw4pR3CuGbw1HPEfwLZMPNRQsq1Etcw5bB7phrwWBidKNS8IxYzMbwHotbd8M6fBm
fITBePHh66tWh8tTS2a6/E7tPHcq7oX5dulJ5GjDpqAtmdxD14lvqPJx/bhTAE6b/Avrw3Q2KCKw
ZpMs+8bqyLUc+9VaENOJtXA9eMXmM1PuBndL9ZjW2AmySHggOfuX9TcnPk9e9zk5sjidtFcI2J+r
zK6u+c8J03mgIsKv/lrmPFvxRhZBBTtBLdUijXlveCyH/ZxdbVo2T+1SmfVhW2KF5TvTyctSJ+rr
ZIUmG2d/MPI4KDvoOV+wOZBY9LIWgjvnismgFzqiCmm28yUL0j4NRfGqFVa12FrBzm7j8lHZrbb6
yAPoP2AjUlPd8V6IMq/R/KofCA3uLndqloY9qfkUlI8lDu7pHnHJjPaKgiIx1B3ClUQBQUNIgNKu
GTTYBdZeF9/M6ahSTFLKfuXle/EjX6ZK9R+UzqpxeNpQaolkrHtRMCiqK1Kjkhgy8OJzhZiRNNqn
0jI1ZWZl90IActJYmHECV99Mi4zM8ciMdUPOctlhI4gvy0oGs76QL+TIrH5llQhY+AYvthCdYygA
C20Xw4sIeFdBzVmMxWw8Q+EifXfFq+acsMG0GEmhSG4JCA7ngPKFqUyXz3Tf/MkgQRE5b1ddEs+x
tv/BPL3E4fP0QVYQ8DNp7y7dFYFHzDnplBN33bXx+IX4YdknKPLT5qqNwUUVdyZMmHtEIkv+utVh
c7tmrQ+M5EsAnVYoZ3MEQTcqrEwv/zEdWMTKXHEnq9lhh8utLZbVAdn4q1Qy0D55wkEA142n2zSC
yraKEYbvSyb7ASom9s0eeD+ya7+Pv4SzkMN4eeKjhu6WQ5VMjlRAOLfdqg5VJGMpSI0/s/1tUDO0
1K7oRN1iyILyjbn8j6+us9Fsr6YGQ2J81BO3U5fihaCtSFZVnhZ/b89fMrcYi3tYvRKMjDwWiEln
zOsbyRFKAjM6Gu7NeNrtKeSCvZb86PihgHKMLZPuoGb/S6WwWmarXSW9+Qi2BEoszTUyZm3mqW7J
aSBy8rU87vVj20E8Swhxq9F/7rMiKilDSz/JZ8Q9a40lNBUGwMvhVe1KEsNDsISiiCF/V76mn9qi
PfQIVw6hb5i9SejaN4SbBZ2A7q3EqVg6gse4Y8njZd4e/ZwyeQVbFbxplZP32ckcIPp0KkhdKrRP
gxZbEkgmJMjbNDA1f0ffjqk5faKCZU0hGaJZiRaQzFvDMr7TZmDH0F6kElS4NrGlHIp1anQHwZif
TMquk4lxoeht4Q/O7Xa8KbyI9HFGLpId5x2cDV3WOoKJ+px2KyLKTgsiJeq+8++Sk/Ysp9F1qO6B
b4SOT5DoIbBicqeOnw1V1iZofnQ++lT51xkg1zZ+gsVEYNK0fPFjMRDy9SD+tEzLurdsaPr7WTOs
eSd6//8d4yYHtCIfH+XOeQWnD4lKAod6uRvGm/iIThiQ8+cXzREj+Vw/Ag6SYpBW6DL8ROhieUyk
yRbb3A2t6sSUdQ/PjUtaHPv0daspl64YSwAA5kOJpk1NQmtiPfy1RJYV6vVNc0oQWqHxQxO6nGrO
GBTxon8Zx/kssrQEFyBoyoCEYxwPO/S8Tau/u2BuPZ0Yp8I+5z2iRwl1y6oAj1emgdNThzuf2rL2
fD0FVELvEFs5uITZZhojRjksum3CTW9jn1pnKaTE9KV0bcpIuwxHwwcGEEb24uM7CY4MVShTSLnH
Mo1Vml7KEzv33vTmrWqTUB+x4IHLz29bMnEy36WR486Yv9AS4nwWYsqvB6t4l6sViha7P9cdH52z
+JkBfxaEjG6/t9SeQWVMIKreH6H4eFGpUhgac5s4ny7dm0jfh6NRVzohchjOIVvsq1++OGT2a9wb
jXa4oxGGJVKOZWrX4lzLwNpqtvhKC5CMNjeyo3MY+sI2dNbb2NfdkofGScqP4LvadVtbb3OwJ8PA
YLf2nA8d1hxvpoyGCTe5UZ5qgP8gDWBvqrYjoLK1OCI6S/pBgdrYpzYdmzNVE68xb+5PJ7EQWPKl
SNJKyFDJ7bEEGBb/BvRtOIB+R3YlH16R682j+j/ftRzR26uw4D9SI+JgHZEwjxuQQXvKJW4sDiL3
2FQWj5xzPOsCsUmZZSIp8uJqoJUgYdy8dMcTJPy4udABMnk+GxWLMzOq3hfbRBBWSei6psxQBDOl
/BE/ifxvxV1JZgsTpqMY3LPgKRrZGbhuW/s1vNP0T/sw0l35qRX+1UGHmBX0ezoh6MuIN7tTbQZi
Bd63i3zuiD+ihMt2CViJIsoqUPEtLAl2jnH8jyUWQSMsApWJ2ayQvKjxI4DvuQM+nfHfrTvz/IZL
EmFalExvMPSc6BSCHnuTlID+islI28AO9jgdUiHrKrL00wXc4THYFCaTOLfYgotXL2ieoXcUq5Si
PAyyZdh09eIquQUQpradIKvUwW1b6tiYV8Sh1CN7kwEBDtwOMyrG2OtDCbLPOUQOY+9q5EpnKcGI
1JTmf2/Z6FXbQ3JgvPEfDDuJHETY5fzZkwP1dTKWvMMGAPZy77j65mxfsScCOy9p0E0/rdHJl/aI
qlSKFRWUs558eoRpUfyWl5aux/Tmo5DoHi7ibf7bsxGelJcgWi+nQBEpWBsvJ2HQmzkyHD6Hb4Hi
JWV0LUszr02ki1KvruuEVTosqwFqTsF50ym++uvMREknS9fZPjFFpTrNkaBpEmbM1BGqlxuO8ZpL
nx7vnNrUhne8oD4JxIlJk+nVWyKeTgTai3DfSMKsKC5qBD/BKZG2pXMU+MBYhbMjeNTA6900cehI
FPmMrASk2f4UJnvkZ5qK54Gg/gYJuDf5bwq8r6DIhqbX7zooGf3R+Q99bFuRsoD8MRieAlmGLSzL
LTvFV5zqTi69Z94vTtKizIJHDsqZwehqxobfRZBNVLB622KzitaFGf2GGQh6jGvSrzVmOwJOgeq3
GmdTNzy+1Ul9G88YdKSloal4S763lBrZHyl7ujifekYtfy1rKmlj3rwAB0yHJCwNN0JhrC/Zr63J
C5Sho4TgJLWN0qjMP3lNAkiOIkJf7pxsq0REPRdjzRt8v8b5vXT0Obnt6/YRKf44VLoj+TGrmWX7
cBNaUfVmDBy5RRJYsGIiaGa/I8+CIfzoFVxqof605cgrPjZ3G+OIRUZwdrF6Z2NdvxxW24e42FSE
Og4cL0jZVRaTY6lsjxSIm9LimilZYrvoBPvHklE+2lX1ugHG+7Mdj0HH3WyvYziEK0ETsGEnVQIW
UJwjsl+NbmmMEEWDjMaAMnCtlswx7sTv9pbRPJ65c0z2QRdpoCrMtYE1s9QhsmjkNCK/4+80lQ2Z
j0mpbrjncYiuhfGfKFhbFlwnxn4B9UmFwPjTqBnZhspS7VEx0w5qQtQMf4T9+W3or1RL8++XmL8I
FeR7klc4BF0AxzA8V4YAv8/hbYCGCdCEh+FhcESbq78uXsQRVlRdblefMkX98KVeZfn/CWikKBkO
7Xjt84ok24G0PBJXkxeNoNer3bCQASQtPSRHDABqqQUQ3/OCi3KcB3cU/iF2mHhbfS26ZKr/PzOI
3+anNf6Bj7qyx+oLum5LFRXTtdYYk3EZLWllNT6v+Hi2ntUoDs5o0l5d+tH+Iwo7TGLf+NLz4VNl
r7w/x8XmnK5xd7LwZ28JeTiaw1XxpglpnQzvNRa4MC6f8nw/1XT1VsM8WgTzoqtQiO178vzIMyzH
GaguqZOn2coJVm7rjC5VJEDgURAEX/3Ksq5ms0wnmWqXeey27REUQmC81Xq0OpcQbdDqS5JRdVfu
gxlGdB8zpGgGVSVpnVJWhHrz9VQxBI0ebJDY1HZ+aZNgz01nqrOLRjfrh6j8nvN7WlY6NeP/yJa9
/sEK+fwtLWeQ6cUsyyCBUo4OEk8u9NnYNi7TE/+pxikXOIqCkbAt+bPNZVVAlBYC6hsa261Mma73
XCCA+PFS3v+ekxYlNyo+ycEQV3XjHei7ELU4NRPUfi1XrHdnJlQ5mW/rMQDJmJtlyaZr8YtJMdv5
DAPoahxbR42p0RQ7JitiiYnQfbjgVX9mvBgUg6/c9Jc0Str5f+hD9wSiSoiYWoHgc/wP9EwSB+Vj
hbXXQrbPAnDhM9eR27nQZyOwbW4dCSuLPffIs378iQeJw3m3HpSIwFMhRik9rv+N6OWjWuMttSZU
cPEyXJzgcQsV9Lq+qOT4nohIQur7FgP/Ll2I3RHJNBb7hGkjN1e1iTDZX2Wn9QIq/tQoVfBTI2Da
wuesx79ivWyXdrCiUSVhfPf3vBu9dBa2DPnuqk2k+fxXTmT3/pvGDGW/T7AQ9O+ZwFFg1BMkjHfq
B1TNvvotvyb1rPs4wbN44EVSA47ldrzj0wdHIr/8b74ZrI6ieTsi+qkoudieMUUEczCbOvMveIKY
x/2epcajsjglrIWkHonUpqKVVyv6kSwMV//DMQiOSHsnOGjUYeevJUvzRTzgSfXQ4cINqX1PJXVi
DCMkksMY2qfzF9lM2PtwMT9Jrb34NUu2PjuHvz2mMi/gltunTmUzM9Yj1PL5QvHd8Oo/csdRSgCF
uZlYdUq2/it/tvX9jgYr4orIkT6jTkjnU3Tf2Pj2tdpGMpw1HFpemFOV1E/darPEpCntfJ4DRQkm
POFkZAyDxC/jtxnu3Z1NaroVgXQQtIk0eeUrr6gKNTfs40Trl8zr9cUon+KZ1rip35yXbIn5sxyS
Gi0AQKdKSizY1SNl2YEyw2fGE1nzZkLkuvRIk+7ixsBDDnJxtNoflUCekB32IWAMF6MrULbsjXtK
bz8+tP0IFyk5KcOPNISMGFQZY61ZEw5mB+ZBYrfOU5U9ioz7XtukgSINs0mdF2oemgXOm0JIeIfw
kYbERJ4dgiVq8HA1l3N40ylQF8h584CfMgT1BxcvCq8Dw4wwOERpmp28kixEQexYEDNL8Iqvrrp0
BYeOzV//hnqFmCOIbxiRR2hinlHe8FsruCEOjJwUdv2HMDYpnVTIkA4DEmTV6mF5M+pN3qv6XbfG
KZ8iZL93NLz2V+T044Z1g68NEKw+D4/iKY59ABjtggrTxBcv/WqKaTt3PfSFp6pvvnqQfkeCKF1d
w1mBF8lC+Kb5ENXcTPe3dIZ/m1GVRUFy72BE5sXsaRiWL3ah7EiUOVrupGrSpRKKA2DTGKn0oT2M
Kcw7OzPMu7b5Pz84B0diGE+xJyfW2B0ruyyJ4P04YoDmaMRvF0VKahYcxHl2PvmulbXaCMQXwFir
iJNO3gtN/+tj52/mRpJ/NVsrxLuCo5+IPtxhoY6jQF1xlTdoizbRxY2/waGlyfTTrMVwcfN3CGF+
68TDcTkmpOcdsjlaCTgkh6TnWIy8vwjkErx9QIN9JTz5yYlhCHgHAGrFfFiLRc+t8ISKxOiU9Tdr
2qj2l5CWr3Gdp0FIZylKtOiw9SUoeAa1rAG34+2BNgjABRup2oOKTTrUZnAdICUtQACJCWJZhK7e
Mrjl3CE6WApNzy4rfjLkoUlyGaitIoNFdxkOFlJXUpT3j/aXJwVCOZBEEYgRlNayyUTQdndd0cJi
JO65WFEN2JMMZdppx9b1D3wdIe6soarruUtYlC/r4Lt5viCPokMk8P9zQQPyD27YZDiTgSYcr6Sw
zyScLTPJns+WaMyvp3jHhmnW2tvxl05BgxKwROiy1WcXPxUSveeTpK7qA2avNRW+W3xpPK7B+36W
qudeCrCiu88nNVTOaI5AOgpVRvNoahzgLP512i9aMaY8flOE3LgLZu5zKgxbVwEAxF5iKGUnPBHX
W1XJDoKNFOBafIVodtxPG+K5sKe1FKbjxY/qedru9cDis0yBL3W/ZtkTpDzpOB8SbZmva46p9AHa
4WUm1OWUp8Oz5pKljrzNrjHyInMOV90Qc/kBEV6G/G34AZRGQXfw5ZidDZqdETmYjpwBrHl50T0b
TBDSPordvNU/OKfIbwWA7DDzcdZQFMGRHJmoq0wKPhhM9neZ97vBjF6FUXtsy/tuGCJs2Fodpmes
D7TJEukgFYk4vx71AvjM2DUfrOv7LeudVKYiLZTrCLCkRi7/fBDLLLu/Sk42gs/UQ5bP3ulvX12u
Mr4CF0XWQ38mAmtlXROPfn4EERgZeiPJRZIhAuSwBc8PCIPPEkKcGBwasUsAL0bJ85ncIoWvE5aU
xCbRFaIH9UU3SN+y1YI6rf4Gt8QjzhSiFi9DzslzqDaUt8z16dsdUCDQmLE3iqYk5/3j3klybPG6
rR4NNe/xRJm1TvTPN3k0EZiGqmklGvoQVB4EUP2vbVDE236nSCa+qrb8geU8iaWzPf8XCVvfm+b4
Hh2pORAywLNSmUcZ88z3LpI9UFXblaYPhHcE5+VfqbrbgdK1EyCYtHjOXsbzh9/FelWuYTjCgvde
VtIFCCRZMv82VJa1rFnMlK3xMKwc1Ca4LEbCLLb8e8jR6s5eSIGSE+/QhXU7o6w31nxzA+s2a0y4
oIFsJtlggUQWI6STyq5qkwaFF8c8hSqjnouIMfxCNeRd+KCFfixV3Sw/mU31O9rdz8dI0ArTzxdh
XBnDAlUHxs/gjTMfjyHVcKLp7+rfJWjBhW+iEdGmIbvBxqzubZBUCTdMsOQzRazjwqIh4vyo6S+R
dTxZ60pts1pP0zVs7v8iXX1nYNYLPrz4DtrHHczCKB+vQA4CKl67vhvprnoXD5I9JjYOqOEJiNq9
btUy1M9s8Jgr0F4B21nmoMcwMeufNt4lX4ghVrCHejq6sq2Y6wtWJxxfppjlVC9hrZlMju6U84B9
q7fkyk8vmy9JLp0PFBSFSz82AqGIX+B+UAvajk7GhZN2hVgcU0FVaC4psJJPmtz0fSVpFQsWVDR5
qHuJ7H/nWD0QwNBmI7ocyRUBra2xufScTt+V4/CPKda/g/VtNEo9fEi0wR832SLedMOXqlXs4OLo
R/wnUgHPl34vdhLu8QGx1U6EMMEIzUsxKKlU0VP3oW0VWuNCaHvUOn0sV9vju52Ef7yLVH941xaE
pe7R43GO5CEHXJqhJcXEinbZvV7yskTcMdhWQI6p/xBC7Kf3CzPtgT45vQZ+/Z9Uim/z2ndPC3Vb
UX9LdAmoDRRKe7mY8sgNtaCQ2CGLUI6POnnJ9e70Rc0Lu7noSIfDfNsCvImzxExhnbCv2MU0plMk
c3lyj64ZBFSqCJepkbdDwo6kH+Y/dhquvYLPc4gnBmJRUaXwXcAzbiMNuWO97pVQ8lH5f2SJDHg9
fm4h7ILseo9PUcIBQ8zWdCWPT4E5LWHbeMOqwvmAZyFeHmZHC9KBZbZhjJr0i5hi5WOS3xnDPuHz
5FPQvuupmMb2S4jEdryypnjCDN4xLX2BJtj7uk6C0q6K7QzvmdYdJtxU3ITZdrEwdS5l3V21sXl1
TihjjrjVdxhCHWj+Zi4+Jl6iQLF6+mDY8cRqhvHWgaVESOgGMkh/bL/SwhpEIGPyAXpSWQc02NaP
wZlvCDr4vkEcpRHcoPfcG5yxdYfdiBxr8sOwjWQe5zH1pBc1fnFGuuPxpfdR7SS3NICJWRigL8jS
Dq9HuoDCaYlxqKolFiNhZJhbHoA2X9dawTAhvSXomd8aT/6nSCVzZw67VjLNaJTvP2DQzczKGnUb
Rz+UKbAXCi0GPY0pw6ct4yjocFWGAmMWP6PkuhZMaaStCHNkZL2nH8iemkcYU6hviDvo+TFQQHBA
p1N4Raq0H86g7JmM7apFhC24RLRIHOag9B4A237uAxLSNfhvOUdIwz4JRDT8JiL9bxjk3urkYKmF
YwApnhvmZ3AjKqLSyI+OG9ypKqQrzm2frMpOKZ/FO1UeqrU/mhICPbGfFXrFoyY47nV+fM3gCdcQ
1RrABFwP8mX2mwX9YTZttuRXgLJNFD0XSAwNFguHc1eHbZryrSyo7H6ehW6H/T/f8dpU6OMOIyf1
l8w6fvs4C7HCpvrPeMClRXT0iL09KYDbSx6c2nvS70QWNkUvs4QxEUad/ORv9yPRbvGI8rRxLyRQ
/Jgg6IEyAI+zWUd44GYSHZo0jWWsCkklh75uir76PhQ6oN+xwyr+OXcbGRgY1HWIBrwBrZyvI5zj
HtRCZ00AO3Ate+zYTMp+J4+o1OXieUiricP21hDB0GRqW+GAUpLx70FhX7ZXRwTMcuiXZS1uZwUT
iE61LXarvdRzJLDVWPx9b/pzE+nGsdnu93ZutwbZqY5EXFcWqy2HTee3f5lSwD9lQXwSYq6BDnEI
by96/Aw6bNJkXv7ugQ3TQPS/VxkJ176d5Kfe0JVAeSS5yoRjhDpFgvzc0sEApGZFrkzAkdjwFZmN
GMTcI/b+O1jaIhZs1Rw1LwXQJ2+P4yz1Wwndhug4dUWMcIutQ0LWn0eHaBjXv8OO57QyO56GMwlA
wZV3ZQnb4RmPicX+TuVhNrk4t+9Et7N3TcITVgBQe2vB2vy3EI1zG9MyyQdCc35ZIGj3nXex3kSM
74S6KaNEGhVC+bSR7wf9JNE0O3dKe1t9vlWdYXBzh9SxKwuWP9RFIylzM+eZbO36tYJox69PzEJJ
NUaQRcRo0ITHIUR9b3szQDWjhue6N+RiZXKi6/H/ItF0JJn2Oq9eY0my2O/1YTXxD+h7b5qrr4XS
+pLpzkwnYa74WszSsTl72Vpp3doLWbDM4Ax/Dy8yMHTF6hMKk+hPxmZn2Yteb+FQXbopG/YHUrzk
D7Q5Mht+CHZ91bY6KHp96AX1ukYACGt2D/5RAKPXcNeiKe0tj8CVGJVpbunKRH7V/GmkEqEu6928
/pQUEXfVS08yaNmfG3x8huitWIb9WhPDinQ5JTSOCr8zdSyepNl/Eyqxx4FafGNBNCeybAAyzyGm
/PRLt0CzxAwhWAY1oGkyCXDe39UIRI5ceLntSQ2vm2YyCIOJ2uOBhEn0aoBB7SG9/qP8d4tEYRgz
FHYAD7/yj5URo6bobuxBqQD8wKEQaLxy8zH1ubLG7MnaDClGDoywL6RAF4sKoNQTNTj0cWhO1JFH
LJkzOsW+8PClXiqJzS0esiv7X/R8n6jLwH7XZ2WRO8Qz5XJ3I2d7Ahf5QFEJeXYNlpr8LADI/3IU
RwTs7R7KxRSU6Q/3mKAGxr8PYuC8+zRCYdgoO6IQq5DBRiV38A6vvHddbYcATDocv80QLPpz0jYU
smWHKX+QpBum6bEEgsdaj2MuVprKwm1lpHUmkFsFu6NlM4X0QuN+HhpfOrgRbLXsh6Fj8NSC8iEU
gTc5K3t+xLjrGHXPAHwHwIiFQ2Qr5yAwqt62V25AiylVBqEsigC2uclzzT6a0c2qm/7PNAHVnPuO
MYxuJPFaQSeizttq4xnsEejMR8SxlFkDYnxraItVDTjHU2B3WnPC+TGZQnM9SQqer1XbLFUS4D63
qJCoC5Y6GgItrEQq1VyDraWznuGxGEgXs1ES01wdLpFoT1PyvXDrGeUMfyskzQysFb91M31mNpvp
KZ0KYwQK1tk2wbGBlFvw0HuV/KjrtzKi85EftwIdUzRQit4lc7AMscT0KOwsCIgnxqA2wrJjgipZ
fHcLgyKlM0hm7Fe3v9iC3Ul1+AvgqzgwYt5vxvEX6SXZhAVw4IyycPeMs/cU9n42EGYbYynysXQj
RcyJe+ds6sf456tdV7oscOWeLlv3BFeaPun7Dg/Hdl09idc862OzjSMmAK1WHJU0ffT1/VUgVt6M
5cw9L+jn8E+DZSZ2ocCfzYWnCoNw0TzfAbH+8lG84sEAN5+GEnNmVYmx30NC1QhyHZPcdEi8NkuE
KOjjJ84SHEz2w+tptGtv+k4pDEgzc2KaVJK8oZWd6mjrH6A10FjpgtI8Qd8ftpT7HVe+84hrJzq5
HryAf7XfxXT8Y8xHdoh/8oB0C4ZybD0KsSdm2eQmradfB08pWv2oYp6SXxreOxK0SpobRl1KIXKQ
ScrxYAadF1x9Ymy1V6/X6vmq8MvqIUUh4MxsVRdneqi1dA8wafMo6IPAji7GxT1NCOGAMP1Yxchy
aEm+fj2NjeePH7hzlHMBzCo3QWWsPgtarKh40vXBjQt0LBApjaR+urrpgPlH/PkGLR6Ghop1raGA
joQJtsYfYAADSq3MLxfzANx93iFcSDjJ7pJHHFoyyclSKmX7srulu74w/auLFc1Eb+FDK+aAbOo5
PeOnoHBmyy1i3D/3P0WEpl6LKhb8AMq+Cy0FYpO8jNb1zzbbuzo1bRCz/+flWpFIpTGWL/IdA0f2
00bMm5T/Ev1gx19DDgm/eKGUaVz9EBfN8ASU1P3qQj3oU/mYsOoHgGLEiYgG0NUfDYUilkD/9bs5
IhTLhhzDzcFqP8VYikZdaZoL9vqhiuruOlMQVboGEJrTs5TpQL4xSF5J8nk94KFwWveVPiUGIoRP
P8blDg4U0nddW4kQYttCwV631+YJzF+k7sgkCnIWnuiiwj0WBu3ugJGrnaaKkrROPH4uZeZ0VczV
An/wjn+Y8/k9PsU2Tasq64ozNqhvns3TD/dSHVdbJ1tvKQu6PcKxf98nVj4NV6dHmSt9+5gKRUjW
drsAo8xULEYEG/8uITSQ1SpK+3B4xsnH+YbJRs3QlajFEkPGGcNv23I8PmbUwM3hiN67dnc4e7ND
RO9zNQ8jM1xamefTLwRl/AoQ3aVbTYSaAHPENq1HANFREqEl4hD6rvS2/ccCsS9g1mPORtyUhIcz
hqV45Xz+YEwFaFl0a/u4G7oUV8VW2ZBHrZS24p6Aqu+W12bLpT4sbsPf5HWRdvNrwxRZmHC/m+O+
ukVoSHIGVzpX7lZ5plqi/TDYMQFWYWcTJqQHojNrEUCWivtLKOAIAaEz7eLUdSzqfoRRK4QehpPR
qA/J2bhIiLdkHkI5T7TOyuOZlv1G5mXVRNED8ec3SFzdDwvGynYWeIiaAAXqsUaGR2l0bvgtNv4x
SkMvHEgXayhnqP8HLG6ioENx2PRWTr9QA5YBqKXSkX0366LA7zqSz+OGO3gSPsFgbxxq+uhhTqDm
33X2UQHZa4TpDv1D0Bs+dH289JHcDoUZG1Cysw/q5JUjLLXiCIMPYd+BEj6e+bKViai54JSxjno7
d51J2vwshLRWhz2cmZUQemvoMAA9oZywwhCvsFuuCrDU7V+88b+Nmc3pWcjBKCS+PMS9AdEMt1RP
dVB9gBct1qhtcekvxcP7SJUt+kKKDWGISxPp4VOb4VHHraR870I+3WJlkjvYuS6SWCxfyhR3jZ2l
6UI0YeOoIB8yqstL3NHIeq1gyVOHe+af/LLapqrbFZW9u3aI+Vlg0+yq2RYr1zV5YHc6fmkyx3YT
5LSatH2wDBdzetTUIikM9WNxW7Npc/5oWvqEHzGT+FJW8n+wB9LTiz6pbhvvAN2Er5ufZUW7OXDH
pysTrh85YwzSptnc+bPNwCQoPoxYy3vbQrskiWotMEfTtl9Gm3rw+k+8i9oC+45tt5yjYaeQ1XGP
FxpfPm5Gv+ENcqDdNi3pN2K3vjqONEKMCcCO5uMGvrvj6ZPB2yqGMIbtE3j2OwQp+M2xeexLJ7zq
wn3c9V4vEy5llDiE2QwmkzLBXQ4tvVVQHhjJe56HBDIAfaeTnst3ZnOq/dm2c6yWPOKse16O4IOD
UIGRqVOpcX9bM1updYJeRwIFNJVH2IvoRxYGCCFGykLD6m+ijdTvkcdnvjyRLXiB/N0ZiR1oDsOf
nEc8Aav3S+X1TkwPILUtQIY2+cUOfx7BEAFW6L5L9kAiGSFw2BZH3uJhj5GDCMmPBwPNJ9n2OqVg
Y8qzkU+XQTWN75fVClfFdjGXTA0je9QLpaFKu1w4rcEqD4G6gNMIjX34olw4p7sInEZ/LhOnb6FI
FL7AK69u8nXoJzFzFmIluFYLiew2LkzklZcVLEKFpsGrO3r44gBg+W/OWwvXYYqUPswV0Q8S5I4n
lTzirJQrN7yi1pKHr2Ge9kciqp5HFJpr2irVMCHl7Y341iUJoO5Hiyuy52p/DABYJgQt7GU0Wk89
pChvx+4orG/+9AsfxjYZ9wSrVb7FZTe9El/eSTM3GAa0oC3tSendLvjivLSQzB8JCKdcXRsb6luM
xPJQvZQlEK4TB9s5LX2bjc6JUam8Qeb7PjPUvd4KL6rSDjkFutHO3/lBa4xWuwD2WjUx8hrlVDyi
TxqS2vwVgP12VcNIXrgzhXhIgE3cZCuDOFsnB1nzNQQEUk0ohUyL27OI4KSUgqhglT+QqM1PCgCw
THtkvGHMTJBu+QU2C3L/ZHxMC+wFTAzj3koWmvSUfWF19oXE36y2jg4QBQ0k0QmruNZFMUDO5Uv5
x0s9yyYI+YaODtxmHAgypTEN6JQxMxJY/nYca3JN45cGOmlp8D+9zvw6LsUse5cD+dqsvQE3V8Sq
agw1Kg70nXPNxqlVW3lGYcNAAT4uYJW56as+EUcONuXTxn1HSwBYRkTz/bcK6KJ4vicSNgz3S2OZ
906nAWqn+JL3rgPDh++LccrBdySz4o3wUt+O/CCR9THx0HzOVO5zCHHO7s3s91kVd8CsWh78UgfP
C7hlv+Ui63eE3sxIXGefq9/oHK2GsYhVFgFYTAOGdOzHf+HHx77QrZ9xFjtJm6GLKzCN6ZY2gm9f
lp/0MvGlBzmnGsapIJc60AgD1reRYMpU59WUnkfEANllhDhOcXlTpUQ/5+vnxEXScxjEVMvMIi+0
ojn9XZTgSHf1xt/b5zV6dkemBUDmESg9ZQyn+ZR7xlV58UDkRBWKGWZcft7eb7jYDnegZ0u+dNWm
BWv7n25kTlmWn0ugS4FHCOetgZi2WVpvrjrRIt8LiQsyEDHlutPsyIgyAEl2gDtF0SK/mLhjBHGG
zNn3dqci5ef+TlayE0h73rB9CByg99J3KtCdTybhqEvTp4NU6H16MLEI2EXXgvUs6FNUf+EGX+nb
9CtMmdCKct7pGOUpf5j8VTIMVKHce4NiiIvE5Olhm9vTXD1bUsrCzTxhxyFxBFNof6nmdrXBBOJ9
uO7XHfqrcD4vPbV9SpH9apjdyFmfeG+cszIXk81x4UMH3Y2/vgGXaj8KVDvxhj/zkKoeM+7eeTp0
ibQFv6LuxHzyfyMBOHEXAFMwmIiR2gL8RxPSCgZRzqZt+e6A5dhXTbTrp0GJER4TgYxqhlPezM+6
nJXw+YqZ6dk988ItsvLZWqHHfPRy6L1t1n3Nw8NBu/ZflEDIJkQoRL/I3/8v+PudXMCcwBgbsnbl
caeVWo66yvGrQt3vsQY2J5+NliwLVEW+OxZPfcj1noXPQhsaN2puGeHY9AkgwVSz3m787SN+emcn
dzrGiY55FfdEdClPnQDxzRVUolpt60TIJsUaWYTYWMCScC2uKMAfkR3RX6AF7dKjiGwwis1k/wPO
+XkW9CilbEUO+Oo0e7t+fZam99oYbEmM5/u609EYrIoMziiS8tBDH2tspgy/0PEZ9FRFS8iaJmiW
70T2tTSFTbM4gOHOmOwbwxC1hfRBQ0+sCvl3Qvl/yq2JFPoBjKlbHgo317ijrOAIi2vqJoB3nImO
TTLwk4+Lxzz2JVgIA2J5lnb/g7y8MqdOcyC6HLg19yI+7zEh5DIzGE1f7v3OEnz4zdD0nLEkPkfZ
4TctJxuTHfj57gxv2iUlsN0hEzRvAuAzfK/T4o+nAAgHqquc+ixsIzHjwYdnMKiRUfQt6678lZRb
ADHs/GdiGHwiuWXcv4z94U31s4kv7BXeprhh4JyTDLs9yC3NxSEdIAulI2CgunMLPrPZFN1I3ZX4
AFi6kfayB0LTETOJ1X7tdj2Ton+oE70nSJBCiQF+5UX/IXtQoGa0b43aaSFADugLhwZZksepWmlv
84KjB/80g4G3F4RiJWGqHeAH50tYD9RxQFSrN18514cdrS9VzePyrmTUe70pYgXNF5ogWZprCDgy
us0PxLa7Mw023AWXAUvSssuCNf7M6C0fyQ2B/iCANPB7UHAt0MCgfhH43wuK0GXdlqFxFqWwE3rV
Pr4FtYZDbopN5x5Ub+havmoxoc3Yfow6XVvskUywh6ETK19sY9iOw+rlgapPk3qvF6z8X3EXJr21
ju/YqU5hWwcsyUMzuMphLwSFhwevim/Ly4opp3oP7Pb9Cxg09lUwf5VAESOP7h1y1W8TFw4ItOOF
k7bUMnpExn6liMKOHT48XaVmuXkRLLsEADJ1u+0hdNZ8sLbVN1LM06mjGVnNHtt2hyvO9jBPH8k2
IghcSg3pKrJeuV9tEYtrmpRkMnJTyuHNwxhTDR//h4WREFyYjZEBMAjZl34DabMm43UdwdcMWXFX
ttrY0Z4Pm3bkNEL4V9U6K/UMeIPFLFrFYY/xhawVLTFEc+S9IetcPrb8JT2GMHHVVA3cPUkRUbEb
3J+yHERoM6L7KDEDKu+FEZualIDv0TPjQXZ6gQ34j8KIMjJ7nnslvfEneBcPILXtl0QDhidTv9bB
vfF0s3WPK2VOhdq4IaXSlzGvh99JAejVFXxAbXkMUbq56uMyVfZhqIgGeOQ+D6GpcG3n3r9WPsRa
oRLnE80n6gTQWQqjBeG+d4/U1w/9/vESpOvrJOjWCVhkY0+brzj28kra3U3eXP4pLbHrPtAiI5FC
4vKKQEnNlX19S47wkKsFWWI2jU5XZq4fSHQMfOC/4gxlgBMkWXf4GCiJcs8j6IKadXhANM5w655L
DmTo8lz0Kfcr03AqTNLIu8Z+Vxpg/Pze0Tw7DmQYRfN1BZ+Nkozgn3gba1/av4hU6LZ14di1GwUy
zKKEbF5jJ0tgKbh34ptWgGYgynIJ5WA7567lcFgdscEBsrS69jCHbRhmiSNSVfwkt7/FaiD/Uon8
yIzZPIjF1adyUVsswXJsROGY5vU6k+PD0/S5Mmsue5EtYH9iY5eGtMJnhuBZkYNbQcuOq8+L++QA
0clzzBAJOIpcYoEIj5l2/aWkg/3hmyJnosvQm6tqOjbld+XA5YgqGvPqcqnc0d/L9bxMOQa1/IYf
zEVPuf60ija+1gV8Qb9Y2cC1/dm86kJSEy0wFz7F0rn+iDKjHgF0BUjQZEJa4LWmf/QpkHHLowGP
hHaANu22E64sg6eSMjipAp3ZKAP8rbHWKWJoIkfZy7+bNnpnkLYL5eu4dAGq//ffohSKb/QMbOld
Mpv2hRn31IpNInEQy7/RiDLFQMELx8v+lLJ2g7G3BDtnxQw7nDrnGcHHr+Nub/0PnIKfA3+RKGZ2
inCCeztNb3KBBMOCJVQ3nVw7qKrlzCruPjy/DzNBpkmkxwdZGpHdZdLNShKXAy0GghZguBkiy7hB
driYy/8CjW6tS8cvEsjhTdByOXesjHsr9XtABpmmc9J1kU/wjciNVih0l+AazZZILMuDDlou1LyL
MvIwXdGrSCv3jWMk/nRBXsSSw078ncTyrHrUXV0KRx6BQdkBds4v/+1avdH5Y6hc1zxiKJTcfTjI
s6C63L/gK2X2wTjgLfQYAW1Sxp3bRA3zeozfwZduvoeH2kZ8KTLpvW/sAAM8URqX/dtEpb22aWKT
TRdS3vLgABtjImP7Fwed3JiGmJIeDQYE9e30oAjADNhWkoqeTGp6p/tIdznw/g9aMKLIAFu353b7
c6b0rhKFohptqjIpHMep3n0P5TvfWEDT9jTEVNb/ePRVhYXjqrswTn8zkmxPEpLDrpAsa8GEwn8B
AsrtFFEuBoU3fkhFVXUknogKOSTS9FGXD/4cIyculWghsiVkISoDChwio3VZhRepwpWqj4Tie+d3
yVPLVnpzyU0hDCZp+ERga0cv6wq/sO2BMdmRe4O6+IfOGMplbW4x6IAac8YLSjbAf91a8/eaJ+2S
JdKJpYlie5e2Y+6noDcB8K5rSSn3Jf6GLxBDEV6tD1JgvHx0Nq98xO2EGCoqqO3TvsFhvzUvBXOu
ZKT+WpmFQtc7NNUEGffIZE+YBTUc4+LINQRl0AOBmyB7491aJ8zk2sz0RaMUKYjkTGfyLhicsJkl
NYa9p3gbvYHGolV+jwvDBZfsrSQfwWFaXuP3FvzYMrSCzNzoRF4rIX6ljANnYkYjt0VBBtoVioBF
M4KhtRzBQvw0mQmbBQ1fqrSbMsjb11qS1yxFXEl5PNvxb23xIjcsyweoGBzHGjqrCFfePmZNxY23
a8wGZaMuKvooV6DcUmp7KXOERV36ubO8A+cpPFkclR9kYRAm3gKnpwDJMqjbTbSjRNPB0xEzA9zJ
IBmpYHRsQMHXTx3ixfqxCXrJefCjQYUr0UoHCmjpUACPh54M/s/t9QjjmglV9US2lkbX4rZN7qcU
ksNJpAHlL+DUu2pzvM7oRo61jnnbLHOusd3NFmQ3H/xmCdlS5R12OnYWl3DDqrr1bEDfXN+k4dW8
FCzizhNQCQ50aLg4obBsvH/YWmHmpX4S32U02jzHexLvuurO+7qvi6puMXE7X3S2lixV8FyX9XKH
iQDWf8cZa+eBrjHD+hKcfagXdV87qNjcGgnVA8hsYTgAaVtycwJBPHJmWiI5fZ7r20d2Q0jtPWWk
TiRder68sQx9DerD443MGcY1TWrBsRpoSPt8D1jkqImy0kB+Q2k0yGwTKG9v1Pj7RiGsOOl+ylMP
sMVzN1CobX3DBwTNtNzbDqojV+nm3u9bK34uQt+OxazlYFvxbyj5lDCkZ+QebRkve5ULbFNCoSwp
/z+nmGoBf1yAWmk4nrs5RgW9uvrzUScx/V0qvkp5vf+V1JAw/JLMP1QMZaSH1aGzlSGdsYC2v8Ob
1lYOmm3b3q6mXSznbo5kOShWhdBMQ2RpiZTBcHwxcVazQm5wW8bjlG8tk4nyBkU0BGCG9o+wpXxr
XjoLLTSlo/HwG+UD0S4mttS7pim9KkoFnRbIB1Lsk7WgxhuB1iZPsVHjec+ZtxZ8GHXc38k9t3lQ
Tm99CS0A99/BnjG5trh5RuHGngz6mCs0yldBiVja6jzMmCA9f9jrWAufYVHDKs4K7LkaFIUmcZRr
7Izf9+ijIOrP9nzbIKiWGSyQPJ8JUh8ubgPrtJw2du8/B23u5qcATw0Xe92oGzQZPd9V0+HId1sU
k8q9zFjGTISrBC+sMTMF8NQCjuhanuP8ke2n9xeuR3uhqc0PGU/dYK2KEQd0aA6HJctfpxBBTYxC
ihMGSw2bfusTBIpxnKQOLyqfHc59R57bBVESgH2oxch/dsbm2scRftprYUDIatX+XzpnIEsnI516
fsYVa6G/9aTzmYUq1NtQ0XUQ+P+dsu0rAuzs5dGQOQ+TXODBwp59cILkLfAk/vSregqr42oo9xUg
bQsB6htvzs3Dw7XwJ8rt1Ph67AW3OBV84L3iMlAolddHtmvD05JR2OZZnmm6AiDsdru00oEbbjAI
g7RIpaCP+M5uhQB8Jdz/g/X3RacBQ12BrUGfZhRV9xfA9wKBWgaebHIb1N/xCOudv6hM+4xKuO7f
meacWD/04JzJrUTBy2xoIBWkEsjXouAXmP+5PKMaDx4SiQEuLHXVF7FbnbD9m/g5uiTr4CtHiqch
TVJYHG6nFBmWk/0lBxNzs2AITzUUB2tEBuOuDZOsKVyflCCztpv67DWPPaDTh4Z9NIlX2rN6s0GT
SIlZDK5vqaTnUaqOS8cHlegRn0paVzEZqTK/IgM8Lh5N2Z/HnduVt9T58AnX2fdgzDz0uGSHpBji
WcuP0kbMf5ZHwpa4ttoCE2om2L3BjaaTh+Y2yo+a9PApcmhhhX0qtz2zpOXKpugvvT6TbAK6WvUn
gIvQDrCEuRdE/LHtHCMfAxd+dd7Tz5xRcwH3+Nm01AREeHCX1CD2nrIRiGPaDy04FjXgaGHjabCJ
Ic8pJHqnEDk03EpnQnM9se/DjmiJ6dhcd45qnJ6xm3jEeOzJHYaynIYuUlDC/41qVJGIXAUqjOup
Wd+l42Lgy1ZWkH2+1/MpSIR0WxJArxJj7/Wwx1WDiHjJQiejJCylI+3NQoH4exRuS76MLUKCJVGX
ocwjJa+Tg98qE7UD+uRuK1cZ5sJAxFtqD/AZMIuIrotY/pwE2Rr/Bo53sct+yOnPAMJiVa25r8JG
ODn6bFAq/TvechYroPFzXV2Ih2v0NV7anBNe9+NxyJzCkeJ9sGg3DqJQZJ18xkJCqtTKYG0XUMhl
No5ubk0RxEXxmI+7/VPMljiouBmxALrSn+tI+gXmrxUnfD7QjVsMb26nohM8JuQOFsTUReWPMXBQ
wbK2SwfAQuD2trZ25HfjHdtxFw7hP3yt3r+EA7BF1OprwzB68NkAQdwYRiypCAmTWchHtWg6aISP
2c4Y00xo5c5ZtMDNnPorKm6NwrH503vF05nGNS6cJ7jfkhilA3NvRMNYIf7+s+ctIDGp9c1PdUNa
cwG47MkmNQovKZ0e8kzqxnjQOyU+fERqx923wuwKAmeO7vDRmeCMRZKwUP5gh6JLBQIHT8WcoxhB
dJEVoDcyjj1Hj1zqv39NGIvphBpKkDmU7V/2+I0An2mXUhPL8UAC9qwCi7G+m0GfWS9FTbfB7PRq
w6ge/yoDAg8u76jVfL8y811wPVHAMgR9k1rs+9vLedXbuZR8iQ/WRqpi0j/6MdnIUy1ZpHjsT9b4
OQmTuu/ycbmzDs8L2EEeQGcvxcoRuNapmlZB1S3cKJyNgJLYSC0Khn+TM6WmfJANuBKkJoBYOflg
cbkVvPFiY/OOicwcgQHrXxvzf0nkAb0dbstMJgavDl5aOGVvre2OIR8sxmvwCvWI+nMt7wnVWdmc
I4CSMzKij7JJQiyMvSImoARN+LvY/de1AIPRgGtLrUGEr0FIDMXGlasjSoNyEAKqSfhbuY9lKQqK
zcbay4uP7ulEcheXLOHYCeV+JT48TU9QtaRrtH6ODJm27NsRBos5J0Ag+EOcX7XkvMXQrjeAF0CU
ZbLFWJ3mezQtYzPKI6wBk05t5H0JoyqTDFOYzOS5fsBYbmyAa+NMx+tKf3tIMkWQK3j00OtVY+H/
PpBXP1C9cMadmxHJiG8n80t5mYIa4maFzVehtCauqo+HM07ZcBvueEm5gS22KqGtgebIi54YjrKH
2Bbqz+08ge5ZwRNuSh3wKTMYWAZMaVlSyIfqduTE4es75jfRvbAV//M24TAtOEBEhi1utK4gpjoP
cSh1xVNOwfBAj2xBuLwZIrU96OCMZoaoPcJONoJtykYEn3Y17nS+YE2CM9r+xT9+DAXtZdvRktwB
/qosDuGTCP0l0/DaxwkbMiHBkkl9dhq7DhmckiQrmRr+rwZzyVUc9d9NElnaAmg0ga3Ye5jzP6RA
e5PKAGLzlhLMFVOW0LsipUvKyM7ia4NJGCiSEykUKNwFk6tceFyCSWcVH5Fk0mcBBEAHo6T+exPL
IOzTWHucxJx5e0HIAtcY+LyZCznhQEnrL+4ICz7oov61cbVxR4Z2aeSpo/dKCzGgG0e2PlX5TTcV
Q2Z3oaR9AZTcqYIc5BN8uMZZdmkhRfahjCdRSSVYPif6F+VMWIxFY7vnoM1xnxYwFNcKCXrxpR/l
Y1catyNJIf+2BvrJaGDCsuQJCsvrxlY+MVy/YpyabybXVibD16XmsOrl0S0MzbczIYvzB/h5gkZY
xiqScDXS0Nx0aKnx+RKkNqovB0+lmZbQ+E/LDoi9T5g9LacfyQmWD7Pdb2VW21FY9O0ReBDD0kTc
s6EuvGloOGG0pzzz8Ou38JaVXFJ9LZy+D400KSAVEtfhNv1MI2bqz37cH3+TOz2Z+9z5C8GkPXkl
Rot5P1ON3h6BMSkAmNlD0UX/UsqZ9LNOqxbKSXVSsGBKUzBw3I3205JOyIGm7Esq1FtQOPpXHaKv
h5WGbIuITJ0zlu8oloHktUkfiN6e8choxcFz12gHDinkzO1Mr/rNEcBZDJR9XPvXT5NfVu4Uxuzl
9YmIcKMhHE+t53rW90byEz2N8jXIB790huAFJHFzuOfaxkSUJaAR76WqtKskPhYlz55MoHOjYcCF
gEq6EN01A5hjvO0eoefaqpQE/akZxd4/KH4Pk+JCQUXFCBE0xsy7un0wVp3c3NlcKDWiXH68w5Af
j1JVE9dbITxoavhjNQTGlAUORhhN2bqi6ld1ZrsXs0aotOKoi3fXbvAythpVZ2Gsz1FncIjsm9bc
Sn+J8YTBEdabpjW475YkCQA2V2+Qk5WrqIf0D35xpVoFARdrQ4MzOZa4dOj1ljtF7sq/02QA77gv
dbDsYeRncqDiFt5MQGbgcJMsCnbL4+M7PHPFHT7Mz/D7gCLzfKE7x1i6F14cK2D50jxwP01jPytV
IZ5DIjn+pNYPVncc+ABclRrTBlkXLXlqkrDd6VJADXWDFhtdTOHEmz8lsA00+4IEowi0uIUmJGtY
IGwb1hJA2iCzNXyddMOh429dKt51TXJbrUcOe8jFedOvxHKQUrEGgEmkffkn9977O3hRm+bbmIag
0BIe1SX3pQRacy5DLQZhvQRugfQXJMRqjju93py29nEywLLVd0XH5bRIERp5DaSal33yIbAMoYgD
mMMrod+ikXg4wObF2zIRT3lDAUI3/4AWKrEDsDstmRg9JIlqE62LyfuGZl4i8ScNnfKgOYxvrGHq
+Q186XcxZxaKPSScWk4bSBcVCJj3+uCp6hqV5REM3CJca+jBDWykYSUjOEi4fUVv7Jp7GeHPx8xO
boO0afXEtcnItJgeytd5Wa4BAHoOQbSex+RZhMCWuH+YOR2REWlTZCCerCQjmhLMyuLllNKlXRTa
1WUZWO5l/AcEOi8qPFfd3DExe81txucK7nEW11ZWvPRl/cFgmHkigC/NuJhUl+IhigGxxERo6qh3
NNCPTUKKk/fsfS2iPV9f27sAN91m34qQ4xwhowiyYI4PyDGm8x5DD4FzxKwznRh6TkY/uVWWRTqU
GvSKyx0FmbslkP3FosT010wIKF6NPpoaL6RE/nxYAyl53Kippwmg2gtmTZ24EOkbG62f9Vg0oGHB
4FXIa2/BMTKZRXvAjxkp+TaNJqbQ0r7yaJNQ/Uzsx8qk+wP3iiWVSD64DOW5LR2Zui0LyRmbwacM
H6j8Q5w5yJpqhvsrBsh3ywHZnz8TnCoYbWSd+RmbGJjlyoxHhMZRYAoTqZEw62QqYYmRJqg/IzW5
wsJbsD5FIh2VzwPzkqU1dRyD2RW+ikT8i4KuBuvcmr/c+BtZVepH4K8EBpnIsU5YtoyLSJs5sBl4
i/Eo6khJPaoyVHOLox5K/f6p4LhD91K0mAK0FRBt48bB+evQ3q177+VxYl8YOrZI+Mi4IXgou/Ft
Tw93N36YUoPvv904pDtz5FPjlI/0OBJCBD0Ww49Bdz6ztD1FYWbbqnltqxHAhI1m0SSf02o/yw3J
THVyMdWsi/UHn6dDtZpoUbp42JGt9M2HS2ziQawM6pZZ1ahXei7iR3EEiUPcau7Pa6UI60scNEvi
We8/KxlSN0Ss5bmgRrMkG3Tio+z5g8pAe8/w+TAP3cfU21jQLAukNAoudaVpwff4h0s7g4+T3xDK
UhycHBLaaV6zN5/4Fw7TFL2tUe0px2zlX04AqW+I1fZN/QIPI+cjRcbjDvrB/Kd/L90h/wjHwIFm
GEqILMmn9+Zm4q7Jefq6pirTzuWYbDw6XlNMdxlD9Bs17c71Asz1i2il1NcC4oS3gP82YpxxUBnL
r7kWxM8EBivCu6Sn7q9/LrPxxAuHpPxKqQel82S87b6il4c+oltkFMWuR2k0S/mxGdCUvnev5NYS
+xvXSgxxBnMbKTdQX2PIV3OX5NoYIqynfWJHJsrTL/2HNOjq7RyDbkGv8dxXN5HBGGw1IHUBAAW1
3Ynm9fbvZFT1PcI78qEC0YXtaHfaTN90tU/8R2Sjwjq6LcuyXJ2cRZFjHU/ydEOOt5jrfHMwnTWp
QTDCrWk7yn8CMRehs35mwVv3t6kJ3gZ76rt71KNky8+Y97GNjIpUCMk+00Xzzkjv+ZEJU2rVSpt/
XJDAFzoSWEiIXqLnem4qZsN7xaG0Ux3BgHrSnQOFi688ppXfOCkSbgYsCLD9jCZA6ZebVBVoIma6
Na9ppGAOV4rSICx48GC80AGeZMYN4fYEERAisG95frSb/DmM0EiDb11nItD/0pDrrVGtsAHr6bL6
ub1asO6IbzFMcoqYCnoueh4Xx7VXpvQE874/8xEfP7EIzS6UR9hJyiEohD/sHp66G9iteTYR1H+2
KJusDejDWKZCRSfZzmGok4/p6rVaGqM2PxI5znVSNM9P56Vvv6mbTWP9h9rOUWl0WKgu1UNZyNdU
mStMjE4BWhYx/E2ZOJ8S8bUEk0jxk5QQ/5of9O3tJLh3Rnv56f6qOXcYYbcyQb6SPiMPXl60H1b2
3kgozIF5ymEMQMQTEiQNoqiqk78Vz8L22Tti81kUqxhURBn0G7LKSQ4XMD40beIsCuac/ut+ryXS
lE8cjmhyTO66c4PFEnqq4X4iqcexN/XU5PMRNCHeGWBu6lN39LG5HB4hpUY3sqQuIRICjZb6qX8Y
zriycIYFx+N9NbhxlhOY0KHmmNK7EBFohuK9lCQJZv9T1bRiMKOJiSh/IzXYYgcbOhbalYWrd8XD
2CF0SSsOa4/zpiHMcu7IRtIusfRZTz94vwnsOGD+NjIJPiEc74bUu2/KDpuGv+z2f4aU79ervF96
JHX1JOw7W+x0PfTPRqh2O/SPkQKRyY6JYezn2B4or0QNQ6BmMCTkMV7oYSRNYtqWOLw4QUXDYSD4
wqVeSD+mddu2E0bfl18/iN6uxAR0DKKEjpUxpG8QxwpxdPwdET57N7b7HNeCbgM5xr0fl+3GPMmK
qDgHCCNbcBgsFbavN6ebI/mxs/dPEXNq6X1/qrJ4aPsiaky55lVdxtFsY/cvcz0ePp8czP92nXj3
Ti86xmxYZaDPqTehqXDATNzsEnGv9KneAg3h1sThSmHSs6r7If7NRx27VxzeRCZCM6cu5hd7OWFQ
LP50Man0LXKEvrDPSYe3gVv3xtdOhdpkK2aTx/nQUyTBZxAn2l6VEE47VAfzmHmQSoSMOh91xaBX
wOxGe8/fUsic8FWSE2XEx4lxBErbjS7LFt+VL+69gm493kmZKi5hfQPComjaBzHhferCOE/6hLcg
M2aYZ6n7NVcnj/REjn90z/ZoY4c4qwcBy3/yoaaOBpwuIVb6Ok/nWHHx0tHkyXAnTGlVnF4rbIc1
iZ/FCNl7UfOGQ0rEJDQGj14zOQ3xBJJ3AArJUvp8YQ9XzdaLrplUIfr5W4q0q6nE856U6srjtb52
Pok0vtK2wLjFWZNTDvqzWFXBrTw6jmnu5zg7Ei5PHgnv4F0/hPxdXkdOim5XyLLDzAJstgAAP0rq
a4K4A3jVKkOhD+fj8NNAPFMYT6pDzkkOh3xeB88lbd+r33RVM6fviFXwPu58srxGI6ugKHl69rFX
nVQrXWwNrONoGE4Vn1u94D5zyl/exqLYC/tQsY7zYmjLhhSt6tOHxmdrORMSMBOzHY8F54oRqLP5
bLSYD6aeAJmGU5AdqGMmMlprxxCJy82c0HJg0xoXRiKehhhvoMdnfFHoRVqNnoXLsUj/3ZV5K7vS
bo4Osl1YZKLYm/eJgCJoNXh6bqz+96KmFBwJDI4xNKARNLNZyPj6ETsXfmXEG4gpJ30QzqEMEMwx
ALRSe3irlxtHmfqHLLC/VmzWf7bhj8lyH+a391zIDIx5b1RaQ+0HPLNU6bNDsFkgLqv6Da9shlo6
Id1byx4sIOjB5fV5GZgrzdi8AR3tWWvnFNsBT/J58nbyuM2/nb6QVlnD8sZkMDRuhzh73Vq8Km2N
nhKzMrYiWtfPvxABNtjzuaVZPQZASZUjKA1XozsyqgIGPusVNC3hWifqnFGfBDafM8x/QJ2tO+Dg
sDEGneXRD1R/6NEbRyRTvy2Kiv/4AWx1MjB9JuZ+I7OnNvrNdEyGHcLfV8meGl9NY00VyaOdWXLN
TPhDC58Yg1XsLFsQ2AS+BLqul6Ojau/IBd7lzq7BzBtZ5YnkCOZoN26PPhN+RGXIVzTawalxpJw1
72Bcsut0aC15wjSmF8DA5z8Vh7eOXII4onML62clqq6VSqfwfmpK9Rv6tXy5j8whnoT5Z6tFHykx
jZvksSaKM1VtGF94lwJfu4S1zrxQLwmN/VEEY+aL5y2YRjWDHNV1CgjFtjz8gcSabDL7AnKTN46L
jU1uN4jT3/THXYeSMTdTqB5C6pTyPQiPRZJUQfw4uA7KgxHoQVsCIZS66GDknCoOeYVv1Nv4onXg
u0Do5/f8kGRMQTwXr/TXNxzTfxTGYUcogz/+R+AwXmuqCgPXmyGw8SraAqQzq3LkgQA5EFC5Ee2i
DEF7TCn77kPvhjg+j970OiOZS4IjZKZYfx67a4YNvYCPRdveVkmJdh93XXFMJVbgN9vGuli0Q6lU
y6uYnFF9Stu2XugEn/wjjDyRJ/zHAstMuzZsD0W4327ELRaIrDjGTHsQYwUKqQOtTCVkYTXAfUfJ
lrdMxWtbe9zZvXA9lKGRF5JxezyqjfpAV6oE7mhNkxrXLs+HRyhkmKFzVH2oMmY+qe2ohwfQ9NtG
iRTol8nfsqP2VwpFWPJZP4iqW8Gqww0nKspi4DPFDtFOdz3AlzeUvelpM/8KyWZd3HbGhVSdLPtr
LgU4d4emWOr93cS/Prg6C0cQ+P5UBrxY74g5wSCWcXrfa3NSA/yuTP7qK44nTPt9uDtLR7sRxm5a
LGIyniAkzh4IRA0yN9rUuHZsxqHfIaw09DJAuU4H28ofNfcTJE5XxwLJGXURrSh5tNIB1GJvF8Jp
vGvBFmCn6ipXuBWGajGKidL2R9qE65pdpS5okmUjInzWsZHXH1SLJwgUnu6gvIFQ6tVeYHKdBvZm
0FWTrKgmYswHCiG+MdYl6ucclqwpbVLlpAfiqRcYUnRPUiYyf9rOYVByQoEz7D4IjjAX6Zu//hKd
+uOzzHbN0TBivxRZKMgimZ4qx53hgD8FY0frw+fxqQMUAkcu8CxC8aEMJzt6QO+FpDizBK9gtqr6
yGi+SE6Loz31zQsqcO+jt/uvB5pTT4z+eQ8WL1IbCT2lOKbKgiFIHkTM97gYA+QcMLCwLiataUxi
G9PYBKSmMR59TAxNGbuITJ1V1GjtQA59q6WCi+bYy7DtKH9NWw6EfMJ3HEB5EyJ4llxtnAc166UN
YTz/dtdqXIV3H3G2WhLrnTFNlb66t9A23C1Av554N9/08t+e1+LkOuxcelOIO4XGwHom8hNK+1ix
409BGbFOfpf7VJDIaZ6+vIVzvvbr36LwIKxZhVesSS8QlAh4apcfX17FVSAFCjR94aMw7RHggsZ7
I7Xazg0X6ep2m4Q91R6GDwBCw1CPvH414j7of184URrWhagTy09MFqqmYJcNBruHWUAjut/oGNar
QDvQb9b1dM81RUPPSgHdljaTjKC/lWpGjv5bqBkCxPOKKJZw6dZqBJiH4mur7dik7RSFd+3Dl/9V
vZ4uiJYkyd5GGf/m69dijYLbdEOqzLWPScuMQ9ctJzDV/8x9Uzis/Q9wA53rbhli32GHHxO7o/HZ
R0l33WRrRi6Bf2UaSzb2Bi7PuUFFDwkGW3ehQEyIQmZ82c0eMbqjFv5q4thWj7TbCECQ5AxsgF0W
wjAV6IazkVfoKuGBG/HiWk7MV+BS9cq0UcsXeDRFlYxwp1ydya/v2KQYeqxSRV3YbkUc1Fuqlpl3
g0U6LpUjiPB29K809gyudQfhxXbOy0wcoxzSkbwfDfHqKJxk4QjEeySOT7/4SIiQRWBnsSMEMUFj
IrVK3VIDMdxKPmH7twGxfVC+sGy6QNwpW10JMXasbHKdhj9m1Mh8lXLVJtYF4y7tWfelxRDLlmxB
QLlSCcD1LigsoKs+Cu9ceyy8LxyEjoYChQHvsZyv1x0yY/47VZ2ExLkwbv2ZTjwzW86IKKOABJ8l
1FUDYQMJOWZpwZkPdcw/ifBVkNSaJ1An/plhYDzr0AoI7EbOiPOavEyhLHYhpu9x2zUmcE9jSy6N
tWjL6LMgtL6UZ9pez79phnseL+JxrYg/RInaoJYJRs7+Ujt8kz78dLLmobAaO6t9Tlk9IOJBijOb
EweswD9xIiiG84GOZctghYJXmF31IFEJ80ch3uQwPOmLqgVxW9TeNU9jQfkK5lr/VPUAoGieicUX
Njmd6wdLwdjyYa6C88e49/AcOrF3Nq1qfrj1jMyMO1rlsAeDMeEpsBcZ4crLOfnJr6awEBWIFaKO
uUd87ZRZRcCYkZUcTqsBrORCd/NWbLw6wHjWE50nGv23A/gOy2BH4ZiKNtDEFGFy7SEzKgK47jOg
jqVcpOEHhI7LxeKOVRD9gCw2lkfVp8IpKnLmiZijQ/2605v4kvtrFslyVbu6JcvTVrHBJYkH5rqM
yLlURtGf4njvsD1pM6INx5Cl2UCH9NBzWvu2iPPCEfaaYK6SUuKlM9CV6R6G6Bh0dzH/dXeyEpaf
u4GEst5/AvaoRj+XYASEg9LSmulWl/eecQ98jCaTcEVhTkgJ7BXls9g+mtKHK/MAlL2IdahCyqjh
Lxv16S9p5vgLXfcd1HbldcLU7vOUH01gU1rISpub01H+eGlet4vSh8KsP+1A7N15v/IF/5zKlQsy
r+vja/tCBfiYX1BlzswqrU5UL6bVkYpjtFZXBpHRtrqooxLYs+ko5lrk7fnWuMhbjb+QK2QhM/Z/
mPPEYmiazHN42xN/PlMwBIvszV+jEQ5FrMMp0O7MQmRwSYL4N3DUnh2W8lNJkbgz18ymhUsePTGk
1CKDlkoj0iyqizdAv9/MMv5K5JTRVoUaAPW6i6HoOvPu/CWsDIYVKVdlPb2nFG2HKe4F7idIgP1E
JuvljLTiU/p+pOTa7ONh9xfi3TzVzYEFNYtx4dOOSKIj4G9fd6vb+HvuKMSuNrk7Q6N1vOoo94r0
vF0EDoWoJtl/qzohDNFZrqOrYwSm9YJVbSPOncI4IXzItOKA4GzdUpv3XGl5qtK8nLd0bclQyPDg
GRRtr5XYZhoPpCQ1LbJrHD+DcCE3ZqYZvILYGfLaOcamKKrrCdN8VlxnZHY8JGbP4sMeGFKIqUgp
4gVnEzZh9UzDftmQn/FXDgH+yFggltcGvdttHVlj9FLrcD5BaF7QL4jRaJ9NRLiUWvtl9XMaI5W/
AfvcAW10qYSHNgGGMMxSYTqCtpUrqYNScPEo5a+VFSE+ENDo8v0/Swc79qOTn3qu0EuhHfZtL8vC
/C5qkzWs2UC26Y44Dk8fI9WMqOr3U+RTiC0KQsw9NA4Pe9dH7jcOgdTQQfU3BCGftDNNx64IrE2x
+MR4oviMw0fk3YSOqlvVXDx0Z2GDcqG56XHBFywk3bMbNuGiA8/jI2hrXKChFeoyVTqHUWtfjLR8
Bi45HQanlp0CfWAoWgBXlhTtZTZD5F0Tg3zrKaeayEBisrxdxGkGM+HVoEKh0ii///0RUdMYdnJ1
4lqnufM9g3K1QwbR0JTBp181/qqYk4hdqopw5iTm2uOGy4iQhfKGvCtOwLBEQUOJ4Mtrw/fFC8pt
VoveSotsaXb5Y//vQOVW5058ipG2e4wvrfNi4BkEX61iooh/AqSjRm3/5Px8NMtreV3UuJV62I+F
jCwWKfbNHGcOkgVRpFbMyU7uRKkENSfi7PBaJt6CM5zd4fPbnvcbQoIUWTmiVU3WAfG3OLhP2ehv
JpoKukHhZJSy0MTBuaOFPZhE4t2HAaX+ymKe6p1NKk9hl7n/c82dHQAjwEcM25YOfFx7MERVNjoM
7rnyiK2vzTCEDSLL80Bb36GqV4bPIGDQznhvIWcblNafadqQF3Yar+UBtXfsUqpDQK8/1IHhcrf1
BrXPRnomCWs+N6yam2HDU5vnFJbjqY2kCHqYy0zNSbhHIZ7iKKp2S/d0S/gi0Mw54pDvcObZqEo+
fLI4XGTpz/1xqGIrf3sI++A6DWedIvOhbL92zgF1YIjB4pP2V6lulaMXRznJmnImaY1QfdXSjaIW
R68Mwql3q1dh4fIuofJDJ+A0klCvDwvg27eljq4GvrfWUZdosK+lYQrNnJVdv8YMEGhnwyVOi1NB
tWX4uhTddD5IzC1uF0k685HdoSK2i5WYOZlonmnXxwc4p1VQO9c6yzzHpFLxoL8E+kPEwHBlshBG
8LmHwYVa1icU5bkw5Mn6TtSK0HPODnvtoqMduygug9UyuT81QkLHijrfblGb8qXaV+ElgkZ2QNzd
c8k294nNT7bPYFaiJLAkLqC1YoCAlMakOeY3jlEmxcZkomW3w2x2qX187JotLhebA8IrcosAYNPc
ere7GcIxjCdVe8zGcyDbJHM8vhOn+ab0QEO7kKk3gpTp5s0DKJgp1eUO/cmnNlvVmQ6KxdcdbMXs
Dpc6h8ITRlCFyy1YRIE3X4wcngCl/+p9lFV/u9ERC8hOGDCy54gpKqxFZpw3BzIFGfIJoMVEWoYm
NUcT2Bw70ilc0m/lleeITuWJUjPYRgO5Z7zNGu5IJI4e+jVWiRMc3BtoU+zwtvDNO089oRPAj8N7
F3rWAZ0pLaTmEtkLba4V5E8ziXBxWuH4Oy6Cuv83AWMN6OVBfe3hewpHhqIq3S3XRJlBLZoR/KZD
3jPun65mpuifGbFbjHVj4RDHuG2pTGYLAnbZFoel7IVcbQD2nkM6ZVjk/qRNQt+2uQMAX5UhuERy
wEWoaZ7/Qp1mE4ENDv4ouE3BVfEFHKQN2OTs0dtkBWR+A8CI12n0+kvxbx3WQpTuHNieihnXkpTC
kYRwhw9QdS/v60Ack5I2P0t1JB5JTg2ciDM9+O6zgqQhpvftXuLsI4HYPja5a0E8kn8OMShm1mln
UPdqglSIVPfHm0gBPmQgWpyaBV3RBIdwJwGJAt90pp6cOU9cwRcqpD7ERpw8dtwWK4GDAFOZ3J9q
TFtBZdigID/1ZK1w0Gwu2lP8W+xd4nN//LK6TsB7mgz2XlADTuvvGvPmRvY9VkELBJnAsaPy3TYk
8UOSkycqB584vWf/S3UXzm7W742scyZPDdIT+HutN3cFnoU2WsbHaHP/3Cq29tZQm/WrY6isVI3g
K13M8N3m6mXay1A+J7FhwpJtcBu27gHMBDlk4xtZsklzAoaR5f1Buf5LcgX1C8o+ibfy4PGHU/Tg
QRnOSj0hooRro7By6Bxz1O1IV738dGnIlq3BOJJOZt+ETX+mMXIOCPNq+r1Mz/rM6j0KvjDYZpKU
St9PVUW9XNhcr8dBOzMGvdYY3lxKSq8cHEcHumwvkRc73OOABUxSqCMPAgvk2b3PCMhDJFkkrJRn
oZ0leetAhK0PDJztDGnrIGTkc61Hy0oIwWI1ilb3vkrYk8QP3OG977nMEvuQgIzunBPJa4zosnLA
wXJQ1E/UNCz7+vVdZ/T6PrD1TsiqKvnf51GNWBYz9L2faigDKAOI7SWSkKgcxHzwPNkMUi3c0OH1
7lGEcmQtSQrCCwr55TmUeYq6P/++81/jrzYQ8f9eWniwxTQo49wOezmZcw388gTMmq7yZYU43xP3
WzJn5gaT6mPqBH4B/qXgY08Wx15VirFe29+XKyeGeujWHdSVRonHrKJOls4etp3lR6ffammiRYfV
mXK4RzF0L4PPeeEoYUxHWsGceKp3Iyaoq0MevVoZlQptz2axMcQ81tkWtCsa3P8qMG19QpZmAnbv
NrC7Fl5qAVFbFUAfQNZV8MWUbofyAC8VjNH3eCUbjf2vPqWU7YFW7Ew+SII4KdPNPVyHb1SG1ktB
Oao6XqASbbt9+gYBCVMABU7JSEns9F5MX2Sq9i8JKc91Bkm6OVO4OhDrqfxmKfNgNL6DvEfLhy4d
AvnlW0SstV57iCqm98tZMHHpjj9JzUOS6vhQrBP7tOLcW3Dw77F2LjR+P7qIJY7KeAA+w5o2N3tN
UGQpbDNsIUwH5kPKQD4NHBrcS6e2lvIdVzFiwh5INYw9+f3BEXOsUuGE9XHfaWesIGAfjmh3QPfc
OAEoXgOExloeaDY5eLqReg90fawuk3mkCYjPeUz4/5/yXzXAzDnKhQWzMGAnrY6lbvC/044C2k3+
gWd5tLSivCQ9ubTcQK1XchKWOSrBNwMpI1hhwQOweat56jpo4uE+1tQfIu39ez4Zj9EaPwPvdhuL
aNq9gvcxQEinBZd5EqBY8wU7FdLf15ObLpVpuwlrvBp4xoeoFYqXwk8oEiAUDWANypd1XeGjzSHR
V/fEJwOjclNFUYPgUrax8Ygiwm2ITiGW50T4euQlMge4sNZ5qxXkRwGTX3q/5QIGT7Wz7GTe8yYl
ZTdM1mLXQvMAxZDFdK8HylXyeEg63NQeEJEn5ZchhFTfNNgpoNt8htoLXL2Gk6M12j1WaL6luv5c
ZsbSBVuOoYWWTc5cX05P07xR6hrO1UER3STnRu1ZR4uzudKpwtEyWNt9XjUcPNf7uMb61FSo0V7n
Dv6BBB/KTEYrzzNQGy0G3kEx0DRERqtHjgqos7MQEnEyPTp+xHhPcvdsakdBx+PrUvwAY8fpxJlB
MPsYN1k6H7Yweu2MxbL5BCSe/fc8Xxbaxl5l7ESSR5OAkx/ZEYgP5xu3ZYl/AZyTbCCL8yIUXDsW
84i2/q0moLfiNY6U21AXU1Yudp3T4O7fd8FUlN/QB2lWqJJarrlw+oJBCKXplzJqegJjSlS0xgW3
BfbJc8+g5SCxfx4XJPtxaIZuPpavoPIoCV2j1PX5HFyD8THoDw0eLvt2bAJvsNYf1/6BG/Tfy/Yz
XPcNNldCf0ugG8MmUaBeVb5NCz8BwazBOvtJ4ove19PO0uKvKxxv017pK5rBdlq9e90LtI4FTufT
fUwS+FFyJJkc3D7cww66IccNgezfZX0fxvKmNbKUuYTGGidBwBhQ99tXlHwqqBt/E7D+wY8Tgyz3
k47NIBVswrNfKXlLOwudv1xFm/BlH/E6ZHkVmm0+pHbwq0d0QAJTHksOfjKa/rAfwSslisppAik1
hnk3Ux13JQVmLI3cF6F2sHa8nAEt9plobuDMlfMyVzdvYxQcj0qZ7o2Z2zghR1Wh8At0EBa/T41g
VmPcGmZrNQ6thLN0M81bN9s8GmnGbUk6HEqUunq7P15UtPxt6DXa6y3447poui/X8Tpp1JnRB5bM
C99zLSCRQC6A4ZfqKPdhHG2qBwUFzODegtvv9OiU5MFVhTv/oYHCWEiNn8+ecKky/Sz0qN10VI/E
yoYeGZ/S3pJF4vtYP+F87ciqT2gJAhcHyJH4f0Ubi2RVzcq/tOK6nnUsJgqV5Yq8W4d9u563oDhS
is5d+sJscl/gJYw7GOguojcH0gZ3ErEvgSHTwGLwzuSaSFtdOIH3/fDuvY969JLSX4G8MGERC6LY
1fudQzw0bCJy+SReG/vbXNc86wp1ZxPpYqnSWVhpvoJqfkbF/J+zD1aeD3OjRz7vTc9kMPrwndgw
w0QJ/Uf+c41oUUPvXTyQQcdJ2T3f6kfyTMF4961VTgaFLKEzynMgdDOOXHyg8AelA2YLRbnni6q2
8Y+vneYKnPuj3hE4qZtdas/NsGiYgQTXRqwvj+Su6CbHm45rceTwKtFWKcdRoAxWhQke4l5id2hQ
DyCwL7GxjkfRJqQzd4Yl4r7B262hsLqgpZ8kdGu4OYjlJJJbSpG/CDxQfYFSjPNn32ZDdkxcWnE5
xUX4juABr5Sb3EA2GFoWVXPJoMRxIH3WkG62mSLsJ20ud1zWcbKohNNAbeRaHnUoicRlWw/0X+Y5
R6QYOhZh0UUdeeRGEsp0SP8eDAwzm55t4XRXN+g5EPAujE3nVSOZG2GrjBG7DKYe5jvwKs0PLshV
NzTGcg4m3Um4n06j30i+K7cg+qworFYCtK7UOKW27s/SZ+pT7nqj+7xBLQyGOCFTX0L7VvYnsAi/
TNq3EBLMSyMbBAoUnp4gEaE2SD4pSxj8zdECe9sj0wwStqinpsYAi3U9EwUmhbZdhHgWEHP8YWRp
3YgoC4FbqOyGxKbwEYG7dvDv1SgY7YTuBJUJ8YnKEX2iLJqczIv0jh0ml+oOM3pgc2JbGN5IhboU
9Y8ENHJUKwM+ovVEwnYO1QiHedPC2xyDO6vRGjmdgQ5b6uHC19xVcDa4IQLUQQNYx+siYhNZXhFH
XozPkY/Kug6v0ndvnOHEv3JFzpmlEhe3fYe4KDftVjrrsx9hC+06VzOg7xFcaOdzWSCIv31xdPMW
ZTUB6wGULTopf7jQ6HUIRQzNhSaPE2tZxowp1lJLU3GAYR1WU2L6pnQOJ88TiTeOLCO/yUDczmhb
o0ahJ1tTa1LsVL4osIx1l8OjK1H3DMH+ZqO+kddPowjyRfdi6CmJqp9YUGx6QVcvHzzaWznYuicZ
bFVP2QF1Ley+UCz5Pmb54csZWc1CXSyVlbr+oU8Y9odH5C0gK/YBw34wgwJVJijSN51rN6iCpyiP
nIIVDsqvWbfELOGrxrTZ8xMh2h7zONg4Kc+WTbmRtI8+SADSfHv7trpaCdkiNrdP6vhP2RXD7O5H
fw/SLMs0ZDde8IPqW4+N3AXMBmENZFjNSFR+DZmi3UAzSjDMxdum4DViuPbFRCO499WV1Fxiy3zB
X+Ib1d55Fh1g0FNi0PnQ+ycObUGwyfu5Nd2e55rGArJePa0Q4OKDhFpGTycwJcRF57wVTYjTZbGX
+MJVJKp5umO0vmmgCGk8lCGWo4nYCWodJ81hcVq7lmEz1x1OWX8Z4+w9dIFQpOf3tYdrM3vlupWF
v4KR1q9LEzxRIKI5wggkesb75FkeKv54yUI71DaA+TAy61x6DA+J4pG2JhJ1dftCvCLIs7AJJvyw
rse6rMAYk8J9GUEMtE+jChb0LOwaQZEVcyaxzGctYSKSU3Urww8mm4xfcjny6vPurq2E5L6BB7fU
KeHxQdIm/f9tvKCdOuZpg3DNI6fSQxGajhi0n1cpuOADxC8xitLwTr8bN6CuKp1koPaQjdl68WZY
hOg3ZcWYK5/w9p6cTfvM3JAPaqUbt99RZgHZNWmZfYMcM4tn0VZxU4Ggf5vKeCBDjAE5b2KvL732
CUK7EllWWau+omJQ0helN4GXzywYL9/sQE+6Ai1RXJCrc3QI/RPqrN6yX8Kd3k16XoEGDlNPPZzj
zQkdSY+CxjAApSxx1zhMKHWfcH66TBkoJKjEwZT7WvCb3GDeOtm25aQ6o2TpOOsIdA4dxy73nDRB
KJsn0zH9/o7cKsUa36e2TkitQl5HK5OpOb5DjsXEBqCJhvJnfbzJ2HSpUcsyaxm8OCeRF9KNTZim
ppSgpzWrWsVKTrLjJNWOcun25vz1jbAJcxSwL5Acq1JXGpKwdFhDvO3bDi9av6u8S1nTKyW/rNk1
zqVLQP3OxLAF7cal3W50EPZT+/hQYPLyPijaJ/+MALtmx9soKuwsr3GuvCENpGIrSZAjfsCJesxc
HpmPfALphWInFh493ZCptMr1kXs+lebJa4X+/gBMiX32HTttugLroZu2FVKSEwCprBfq6TX7V00n
jj795QpgConC1erHsVvlewQ4oFPB5zbAOCkSggNSLV2Wr+FMULQv1GdOxF+Z4+XnLDnmHI6blkno
8ynZll6b18EvPLK7Jib8AXBU8cNm2HaJV4V6BG7SaUqJPCzKBcFgBV2RcAQtTvAmrPgBHowY4M0b
wd4KVU1QM7r48X1B4rl4SKPEkN6dQ6Yjy1KUPfbzBitwkM2SkcuEVapeC/cDKkv6xpeZ+H3dONfC
pQbvEy0BOpl1+8/6gqmSqEAUmfH387XKAk6VQUNcbTU7/dP0f8wbeWpEfRDOnJPUFY62ZsKptwHP
0yPChoL0woa9iRVqWQasRM2b/iYgd6YenZD141CTmA8oioANVmEMRqpGat7ZBOQ7FWg78HwkAPq9
LvF4H0E1qWlONwORVcsJGHvmTFTXmgkI6Q9I3ShrXspnBFAaPWgq3rFMiKSqYzoVeFFEtRDPZfwA
O00Fx8zZv1WHRlKUQJKhHk3iYNbkit5ub2q1TgHFvQQQ0kGbfCcJh4TGxtijtLfWS4meOxs4fD9X
tGne9q/lbz/hoy3HlNfDvfSWgtcXuXRTvdIlDzonc3DHijHMAj09KwGI0DGLzzF+HuUnD9p71dPx
4ENC7pU68Nexd2UlLVXGwVbVC8zPT5bBJ5Zwm0hQ0ZPp3Vaoy80GEpTFIVK3uLo/QdSBwxhFhwuy
64IaVOW8F/nOsEOJ7XqvOpWclZJEhXij5kYgFWEWOG4ZXc09HroX0FuYvVrxGtLlC/+JQWquXxEI
CO7kjVsZuwnQNB/awaHhXQOK185K362Zi13qMSl0F9eOlyrIS3wb0BDLuPisNa3wXfsbB3kYAXn/
ZCNnMe1kygVUGjxtatQvJ3uF9EyD/AxZMujp+OBiDi8xJ92OuVs28BTqzTRhDNv7EsgXvvn3wRTs
aWZoBv3JCZ69CLRgNECl/ASM3U9SgltBHVZuT3mLwcZ4+8Q6KJMTjM5jrxPlQDMqNu2uYHye487W
WhFQ2+KSn4zu+v5oIXDLwb371xFh91FhJA1EQ2d5BjApCm+ieoRB1Xl3kxQeNZSshX/3xxvx1Oif
QzeeRY2E4ElJL3yf5x3gDeWrCfyuUgHIVccKyxozwF+rnACPGAEORU4qk/viVDSFWmWjxfDLbxS3
kF8uEX3bZzZQCU18hcbtCQJ1iIzL9+v26YtNFliF+lgXxdd21h8EEh4Y6S4KrV5LOy6NEsBRMyby
ehg/mwyIbV3mReMXwxyjA4zS80ZVPZ8SVV+7esMsVZucc7Rnc0LrjUOWEWERNWL7DUGJcuA1n45X
UcrySFt45rqdcayyQxeDE+QZ/DEAv+ljCy2pCcU34y38SPS66m3X6rnAYq9Ve1BE17gt160Fala8
b9eUWcqH681k48gn5LRiAcO7N2jBqiV/vvp41c0mU5a5YLBmiKjW1vQuKfn+5YB08VdAEcFUJCD9
0JS8bG++djI0gxx7iIUQ/XG/9gPA0lrBpvpF5qiMiPGq5K0MURhPHWqAC0SBhZzk+QHxWhoN/zMk
qXVFMpbx0yKBHYwUwDVswPFEHJIW01Zx683cBElKDB2ER75fQi/TuoqR0C4Dl/chYG/XGEG4oFMz
P75LvxA+ZDBXmH0xlFa8I2tu3kY+iqecoC5yVI09jYJ8Z3trC+UYnUF8jysQP0ZjWxTDza1l1tbj
VwG8iAVST6bo3Vet6d0Vxa12YFHf8r5LN0oc3G9vl4PxUNhphWxhgC/zQf3Pvlwe0u4RrE0+KxL0
olFgHiBX8q1fEwAXdZnU2q542qBkSHmq5tkGhQ0izbpFHcUdfbdXmuxNcYoiZHnBezS8GG2MtpVj
6xsXfvcfhbslTZQnbse0AX7/tyuDnNuiTUQDsOSR2tRVEjICQvroBPGAvJBmsNHD8ztY8qUhoKVh
AB/BgT4qLUGvGyAhL7i2lhKQzy6dn58Ybl6Tr8z10TLCeAxPw31SsXBFgImvibUplhkDE3ZsPf4o
ReTRNst2Et+TFUg6uThEVo7z/b8QC+EJf0f7G/zlEIQgyWqDjlaAVIv3vAeqenvJgMv5ZJQAIhY5
+2Sgd9rL4KmylxmjjwEdvwtjWz0wm9yZUUf1EETgEt2lU9E1f3W3uP9gvQR1XXVBhGoK9i/0Tk3c
aRILaArwp2798pbdsi0DDqsHhNWAfzwln5eNeRz3DSkAhQ0FseYI+hHytPYjd+Zwkc+K+z65oSFn
3mu91vceQWFO1vZ4PojL3Ye7tWVGhKvE1ysrRcw+KqLgo/pE8c/HdeYw3fZ389s1rhnobmwOSNG8
aTy8jpWr8/F69yAV3L0wk8FwtNmpK2KpWFv0MMbD7VfwsIH0L1x5vuDpYZ9CM8Kw63+apFl3eL2c
9skfBzaJwc85M8TDGtAgu34f46d6lRMT46KeLvCAKP//0F3mGhtOZYagkZ5ZeB5oVTzLdud1iXAg
U7Ce+gchbvXci5x/XKuwQ6sVhJYlzpG9EileXSWEeuHhbEgCXTxR2OGvrZkufwqw81AuvhUvyy0t
nBRdq8EXqFS4JUC4qAbA7TfQkTWryGq+JCj/VV9SjT/dQyxGip3BAY9JNIpcTiN+HSWjLbMyW9JE
0aJL8gCH7itJJzTJOXS86tBRvcnOotMK8cFi6fTVJtUu44AUZ68mkSrKagZrBCy3ko4Z2TUOiFX+
9WJf2gpA8jJIyHT1RLEOBnbbv9fZMmpdRIPLRrtS3LDz/jWdM/voU9p0KaTeOrlGh/Bf9MsreYYm
62Du2cLJisQAO0biiNEjw2V4HMHqpwubUPx186rNq55GSJuP519S1r85BRWBh043j4Uw+nKTeeoU
vjaMcFPrSiN9Pytn2xKbbtcKM0vwDKEOgALKUHPgwvnMIYqdtrW1Unwqfhm8EBxm8eCQxoJIgmwi
b9T/xvuWBj0+iSwVQZ1D+kXFE/ixOcOMAW558n4dsMH2UNLCHytZvzu7bev/mQrZAXpibb4/9sK/
P7pESnuDIBZnvORjuuhjAEO2rnABeIXUxqoO6lmagU+N8/+tXrLNJlBRZ9hCw1OXpJgSNqyeNZXq
ot7V5h4BPH8qPcwrYyDyy2/eLBToozuDzNlAHfzQtM1v/u7Lnt0Kerjt5Ui14BsZZHJQoWrkhmA/
aLnhX9MSUj2WT0xj2aLjDiPdBWp2kmg7x8ZlN2OmBwBAglZ8TBZSLzWp0wbZC5cPy4g2EtwXGroF
vlzx0FSE+IbciqwvzrhPD0V6emBiFvHWRdnpE0xZ7KMp3fQUPeWGh5n0+eYSY8NDweGo6Gik0rwV
biWlGMAnFXN7rPVc+qIuXjD42SeZsZ2ZfZmVS/JK6r5AaOXWq6Bvqgjo75tdUx8lmJdB+cl3Ew92
0fHdWSEkcwaWKgLG+vrNjj0pTp6o9vkVnndIiZwe3Ns6XK6DMHBr/xsvKah0Vi+KturUKpp6GKjy
MmLygxAfIqoq/rdVrij/iOSYxKEkF0Cokvp39jjlNnlx0504RgD/h5P1aSf8XOmC6CKIeL5mrc8E
nwdqX+vIgW4EZkIq/JQHcfvR+EsOAC4U1t1F4uPNoXEyft3sHlNr3wZEIFwunqsRakiXfFgI1VHm
mgSTyNqfPruwOpkKGLN2XbuiuZa8ujUw3X4T8+R25/MonVFkJGahwI/Ci0syGq/O70hQI7wOrDJ6
J6z9LOvIE1bFrSE1or5CIotxCiqSyAtJkjFZeCycc+3OW+Kjzj5qwsyGU7AVTcxxIYTHMFGacvIG
MU9Cl5cyhBJyhSAN7dqZXN/GTouw7B7/PfXFQgIbjNQnYxaV2FNn20GXbLkWsH6Q2rBQpexMBKK9
KvxGMlPMhwo/4M7K84vMkMNqzklu/P+cGjqCG5yyBgyyJXSaeYNtxfVVjxSRmnaXnn6ggvqTcf/M
QZDt2tViHosu6ovp57QKsUQHefIMHLO0juGzIyCO0ejnSONqPiXFMwjKFyHJeN/i7FTJUoD2Kizs
Rpl6yCuGrqc9iZILb/o3V7xHfW2N7+/URFUlM5obRrOi/L06s04VstJknbSWCeswYoB0woIEnlxf
1A1iK+hZ3H5QfOd0gZe4YKA/qyceeSEk79ygRD5nctKQjUwOilzRb7G2/sq8ek6EezdvjN+G8SnO
mnwXvBj5S73VUj0Wgj4q+NEhfomV1BJDnpHyOArz/VVkFs4aJmQDhin7xzu3E/GsLw4/KankvnGB
+HDReMYXMdCE1adYKfBSPmGfWcog0yULc8lV0ocdRwjegqWV8hZrAmaN/5Z+dZ0HJfl7KQPerEJ1
U0V2RGX2hfhLCRKs0qH6MQiwVsWJpbhLcYlgIx+22sQIJSNUcpF4zmzUbq9mgCox58Yr9sTwXLTP
thpQMjorsYS5SDChAwtyXTVeqMG//Md7kxMqnYN5dg/y6OSfpZC+BJw7AvdchR9zcAkZ1LDHiyPG
EtRvOEZWts8vo3FON1b4oZrhLiKVJMomJpmg4ZvUhBws4vRBmZxYcVepgjsoUrMHRe2OgcaGQW8d
kl6ycUNFHvFFZfR9L/lk0iuh7FKNz1WgsOcEVM9KWX3Z1kANWEmp48MGsC/JhjwIq7XNieZ8VY5A
ZUMHcCPh47w76oS2Q2kk+rW0fQ0FXEsw2HkHO9DWkoeaY6l+x4YOl4e8vvKxedqfYzabJ5yQ36zs
sLs2cWMHNSozPh3HrwWM+3T1J0/7eFQfxLMvYPaSbMJlDrlGlX4AP1ziI7cVAvfxG4HbCMsaSXgd
6KYi/qVdnMazOvC9u8A0UpjkRHpYOHWRmf0UvThv4pd4oQaojBxaB8ocZuUn634K8kSmAvgTNCyU
jJ6DQDKx5tdmhJ1kw8uyWthsdvTRXN8/oJHDlT3ML9/UWk1mre8ZZgPY8fxCwhtwmFsrF06BBa46
MVXNUasYZkOvxfFlKdApEMjVTKmPeWPSfHoQ9M4ZGr29E6lJyGNhP3Zq+2uoMChhU0AevmLTUk9D
R8nHJgIYH05rvRU67BE8JqY2liFYZ8aPME4w7XmyfkgsGLkRD5fFE+NvvrkVDEIHw1shOUn93Ihv
D5vtt0cWA14cP0FddkEWhkTGGtJplsd5q5dXxPzByA6FOrOfMPzjHm27ZfaE87VYz75+EIFQNdou
YTd1pJAUGh9TrN2EYKlVbrqGvm/4qEChx3OULwUrwhRXZ7VPFjZzwbIAjt9yscdvB0L//Q/NamUG
9K+kYLOLnLgQE6r0Km710dWXuNp6AupT6MfEaJgAgjiamXpmg4hs1/bVrjgAGr2jaOnLuQoUXaU7
M9glFbUlEGgqj8Rmta/8p9kGvKWSH7vm5t1Nmh26q4A+RIV1Fvllco5dWok2KgiAlthM2sVh0gYj
wKoMZzdM9KhCOl+rmyhpOA5qpCwGE+rCHpVYdLZueqSqV1++fR1Fmi6IQzpZ66MIjV3l9c1xhzPA
FUYHvQUFzJpyAo5ebOAvTBMgIat5U5BB+68UI4o/NtVVXu7ln6OGP7Fxyqu1BK169ZskJcGu8iTS
QSYeinasVASpuYJdVElxYxlrm0R4GEtuunf68+eJ+fxzIpCxHLAOxqvJt14Mq73TQpT5Cxwh90+6
bXyqG+Sze78g5lHTaUD2B5B6FJt4yIPajZRHN4UX9yGB2jQzbMeNn1fC4zxPUbSphs6nswfak5fF
VgSMvlnONCcz7EGrkeAR4w1tDrftZYHwMJ5tma9IKku7o/+GiAJfof23R6dOXqjoYnT4WQBULQQE
vVWt2WMrQmwnN/nYk2zoDeAKi0IF+SLbRHufznDP4ZzYRiEO6pepP+35DjXl57kdkPhWsRYq3QYs
juLcqTdLeVakMaXcSJYLY83qA1KKUr2YTEbCDAIXGI7VFdhGn+ROhT2tDgQUbD2BYA98lxv9f12K
SihM3tSHjBBQg+kFLsZz05Gal5QGThA4wMJ/7ijZgZ/pD9kGdcb+OyRfZPuSdZMXX1s1FHbxPCTm
n2IOJqU2lKNKEG55C3VQ3N4Xrc7xYgSGEiIJvO8P0sW/8LGUTVZ95j5iddS/coAb/3fdSQGy9JEB
kwRMDCrXmY37EgTqI0gg43rHp6sJhyI3cPSkpJMX0yqDSyvWfGTyBNgxF7SvYNTCDDumaL9ghj0H
uwT0GnUs378BZOwvJ+eMNZ8J9naXI0lg3YHupigBwkERuGSQ92qNalEjRTP0MXkpc7rsb2zDXaqi
UhGQjOix8g4fRRCDUakVztvzczWLAqRFGXcY8gVod3WkEazDTCpr5ZCyqwRdfQwkgXIhX8osqefn
g/8SvWzoqlUf5XtL4VsRwNOJJSUgZGgCK98SjOS7YeDp6hNQ0kgogiXOySCIrCNFqA87bUHd0riH
L7Nyowf6iDiozB40mhmyGgktEy1lrZF+lzuqzPjksXLN0qyOsQ45VFK1VdT7lgQ6ewrsil4DGuZm
FfPQ9Da4Kt5qFXYUHzXSOZukDbrdcwSFUBBkrHlPxd7SRYUR/knHaqvG7k7IcQNHfK7swLyF7Blr
NrBEbbANGX4mqUotpTGs2EhM5WxR6G0jxUrWJnF1hJUa/UOmC3YlxumeTy6x23NZCmvzWdJegL6U
eWFeY30bg5gMcKUpiiso5SZvVQP1hz9gSdtZvUoeoM/TcpuHC06L/hCgdVMAARTLf7CSdx4LxOa8
XeMr8/gxjOZ5StgZ3XWdZKVBhztdkR2vLsG3AU0OTs8NcIChl7bFVthxhNVIDkYV2ajhwpVRHT24
8NikZMQyPEaQuNt/xSvTFlj9c7//ra/MjowQzL39tj6Bpr0npSFFjjv55qGoqgFYLsz8W2M4d1Qw
AtIXZAX2xPJNy6Jsuw4RP1kyVZa2Ru3/sApRQlScwfeEaZ2e2QIoSNvajBSsabCZ+OiwCIofdQf0
eB2zUL8A/L4b2r1C13GlSwyvaP1BjkuOSn+3GcydHUecnzEBlvPuah/XKWTopGSkU97xw3fOyllC
C7ZQtiAFBwNhRFizKj8bkm6h6butykhl+ZlggFmqFDrwSTcj0KAwqz+dWGc0m+5DXV+0r/QmLEBr
JDsD93Sz0vQDQANpb3nmskEX1/u8u7NycCg/b0OBShNjggbvygSoP6YN9RS6HcxGsRNn9dGc8wvi
HDIkK/OksIB7JahFPAGlyGPzrIzuzPzIChcPXlxhXCk9XjKKIAt1zgcedCZtCLP65rt2YPjyLr3a
jvqzEtdvCXjBC2ICtEdzCzilwziMxXVy8jS+SLyOfZSDAGY9s5wLyV+jhyZae4G2cTANOFDtw/aH
CWoyhQ6SJnNxx76Q9njl+DH9tyWr2gFfclW7LYzGAEjsKuIX+5y45csf0u/Ma3jLmcE2Nl7GFrEL
TOl2CoBb50v0IxcwP9li/CmUYng2/mh8RT5CAjxz73N0bFd7PIdrriXS0iso0WEKR4OLnKyVb7y/
vuj6h1uPdoqtmgGia3nPEthjiP0FebOJ98jgfcqmU1NqRgZMX7fKNjh9Ana47s46HW5Sf72Q8iDw
FzJHSZFGQzNEK7ZmmIdt5Gd8kuElfPyzhv4orQ1fyeEYnIJNg9cxSfn44D86AsBAkQdx8DTm1YXC
fSZkJUK1qF48AWPpxP2PegG3GrcEu0vu4r7feq7bnQhsul1jZwLlpopqcYqnQl1e17Q93ddhvKg6
9Jt1EcapZqV3plpbac0bvLtNexnaJC6axPWuBByM2NZ43/GkRNJg6Hve7Ptqy2OhgaTdO1Q8e27a
UxoeAOfyDkhq2rHE9JSyAihEWbm1xbbt8GXKfIfXFuhU4IgxXiDzUGwtLxSr/Wz8So/5sNjar1kk
y5Q02MZJL6zRgMQ2awXzDWfjbWsZpVAORGAJDb24D6xcG4SsgfMsCUcu9pGUzFz0xDxEP/pL+uuG
HoMGLMuZT5c0WlaqTfwx/z0MBTeCVnXcGUWO1M804EeUr2w6efzAxHA0LIw0/TC/xvTORx9P7Mpo
RABZY9JmZEc+b8/3mvSWNVS085Q0TMUArXI9u0fRP3k+6ZoOzW9wQkB/vOZ+WCxgStLAe8xFHK9c
Z0EDDcs0WT7oIT15ARIScFtGPTQMkV6OVAzvAmR1nYIq0SsxtECrgL+lY1RjVzERKh61hd7Fkpiq
9EHq8jF21MAX4SsMGEF5HG4bUQUOcX3o89rkhGq7ardq8swXKctYWnQkNYrHkgY0XWHLKKeyIarv
zqnd2zOoUEvJ34159WPPc6vED5r+AJFJkOnPcpZwI1ReyLYOx9+nXu52A/Ilp2du25ZTz8ZP56CS
4gBlGYx5kfduLjYrKOBrS+EFhE+fpEQFM8V9I6BdyHyJed5lUhouX0ra+CrB13cSfe+Kf2P02uCa
ZvXDEFGjQ8WnJcOJaDcZi21k/9QXnGDAkxj+xYU1a4+gGCKphCDK/jiq282jEoAasK+Bgy5et/L5
nlVbAU75+qwoDIyCiYONpiIo+RTE8T+mXeHTQ6KsVPjzNP8+ZM3eUzJVNA6U7kUFNbRWMEXa8Khq
cRdRdf6mkRbvTbGVeA17cXfnBGj7KGRxImDwfTmI/Xm4BPtYFIaI5Za909mZJ9gXtzMxCDANjV1j
G8eA8lYsEHc8UHIQfQOyY6POYq+HnZ4Fsvmt9s8B/PWxYt5JtjJAdo44GwD/nKmlz8HPDOeaeKOM
lcVjkSORHdpGQ9uQiYcBONbBGpTFxcrAB46tnV+DrEmyDWm+QURiAneK4KJlB3W4VZzZ1nLsoTDJ
+yTLCQ+wkQpPDV0WQeluJYZMRI79VeO+YUMNMaiUByIvQoX+rfAEQiiYWuT7y6Y5joKQVJsysTfx
o1k38+jpZKxeZaxaw1RPhzqlacOvZ8+whBnVLGQ10WIfVAQLzUBnGAd7y+pu8qC9Wgehrvlq3dAw
X2GsXycGEcBVSja4XOhNF5gpkNLjD/Ybu8XQ2qBU76LtATRL4uOk9+W4HX4gMMGo1vSAXb06Jr9R
QSfpBd7R71M2TNktVUchT6ZkNlRT5gnIwToXLG8wz+P2ABnpXnsSUmJhggNfIKXviQlufhYXjRov
wyrJco7ISa5fattXlitCDdvXhx6wwx/A5PNO8W1wL+CyciwPd0zOxL4vUSZ/yDnmCij2pMgjJ8m+
rinv42k7YKtNI3gkuhV5/6n+eIbK984nvYyy9eRTDWKQh6wqslwgEPCA+wwenZ/hxsLyYlgPtza+
RvnZcYZMBh90PLbmHgI+nLQGfgVza9iGV5ad2N/vOuFuPOoUe5/aMTZxwFBebMwTzui3jOnGQlVf
3QYs+AzYPidATp4npKFks3UawJ+RoHVosnIXHwmZmUlhFv4DYYfpuI/dt5bLOz2GhwEay5IPEDJa
Wi4Km+9DlJAFfZbRbb/PA7Ys23Dy2rrRNfIAM+XASi9yRLtpsQp/mYHYjcDvI++Xia5nuvGTW5tN
/vKwllsLA3osn7ZLiyIR62JRuYdmtROtZ69Cprx6xSrCKkyAcJOvJMvQdKRxpEHpMYhXEXqXtAOj
hSrhDwQ52BkLyIKX9rLR2jxNWwp2n1TFXtnJp5Caj2UMHkVCQTug4LNxlnND2HAsYkR1tmENJ+5t
hIlQEa6RLi399vyUtLCxBsn3zEm6trgB45dOqsnJCSoHR5wAn+JbszR+PvWHfiGmGStNZiLTnVM9
0YpR0mw0fAmONqEDGNFemYHzdIThMvHrksxuTdnL9aL9tG8BBsGUxACpkLpQX3XXj6eY/HDTfveR
1McFGby02J8KTTzEeR1K9xAwYC7LovaFBngJJTVHzv5b2m/jzGPBB0n40yp0J42eLvL4FFU8N36j
yygKs63qT+CGPVBH5RT8hYhm1z0Qd3J4RQK0JXUMxTs2voBNNjyvpw+9x9s/8eVlU6d4+sgqlK8Q
YuBYwxCeaPnOLThYUuyJpLSUTiQAUj3ZW68pNTrLygzhSJfKQssnYmJ2Gq/G4mP2LDBPyP9z6Q75
yqiF0LK1RPI1BdLOTX5EQ5NMKp6P7nwMmyf1m2hsquRTVzWIlx16SHr8Cg5//DmqFdTdvZZMo6DA
1NCsp3yGc+qjmUrTquHbSLwZbzxsey0m+1jxcZuUpMgj1nMI12obpFaCmntYbxKS9BGxmjk9xcLF
D4ZZJl6a8WeSXNm9VoG5nHOPuqj0Lp93Do2fjhHzXrqMxiLS8D078ERgJNkdSKPqc1PjNpznKOSu
tdXMhdZX+iSNJox1oAjRLH50meHx8u+gskbaNymndG/84vBZbQXVMbPMI7A+cwTraKt8/8mxjB/Y
HHqzKfnyz2sMZfHd+kM/e/OVtKLgr4PJ3FuCfHfR4Medv1PtlR4jVkefDLaKwmWmQ+yhZdFhsr/r
au13cgOYbZHdfe7u8d/ms6+EDVroF9yV2o2JR735NoKAYNMbqbnOJ7b2cCfwxp8iOLmEZFeQpLA8
XuamoellputQA0KYm8exxvZkHGUQnjwWt/AU0X7xc2h7JWlzzgpPKpi/9pAUA98Q8zRu/EFwynpT
x8XQbxtn1O2lDeZUcv0X9+wQ5z+TI3peiDO5t2ZhRiS3g2X5QngxrtzVTnc5K5w86BykY51+RR+f
w9XrGzosM1+q3rIL5xb5pS0Kj6LJKCJJaVpzBm1ZUUWn2xAFSpzhJwHS0KJ4r14JlgQPtZf/jU//
GsZ7uEpLB0g3OKt/3gnOYJtFgTS4926/RwfsbTAEJPTGUnfAx0pE6fPLuFkJy8jLWykYS7JV3B7t
CVXdIbwH/2hQfxAw9A8XJkJW43AdYaapXYWefioC+CgVVNUz9tahkGGlRpnWUUMuxUJtPt+a3u79
tlbWXy2avvIt2Q5c+lprCOvGd9Juc17GOcPw6zr5/y6OHEAasMKY+IBZoBddE9LZ1lq40bZZS9UO
ma0/qK1wR0M6LrjEwxHyTbGz4CEpK7FU9QqlkrSdNhvdaoL8DeIX1pmqW82bFiwltc9Q79Mb0yKg
xvQedyhGjAAakNBhIqHL3xGbADo5tF9wfhbRNYUFmv+ko9lq+m+z8tWbBaSod8DjkbnD2pABFu+S
Olpg/tuNRDd2YifxmFs1iqb6NxKZZkpsNwPagY9I8GCNvyIPzHUra85iItDpW+Q+OtTcbdgK/J5s
IHXqNi4TEMb1V3GxeQXgAGEokfy0WN/ExfSlA5UXgazWE7RdusSAjFbTMYZbwuTv6TMTRg1X5OT4
Hk40/tPogo5Z7Lkg4mBPeeILcJzWPhhV/n8dKtBJkbhCIkUhsZRXwXQPFbuY4NGT435wAtifrP/q
F/0Q8MSDuwUI06uNR6Zku+W/z0GXCr7BFuxeVwlm2V66mtgQ5Ve7gljmFNP9KUUYLrh201wGqBvm
mbDn6kcGI9V2WAae6uQenioV0a2KplodQ84dhNQ/j3OIKg4OfsqIWv6qwUiH7GCUsOsZtjJBQARp
oK3Cnsl2PZpgmjYiYKx0BTWAxexCr2HLEcuYf1JCbmRMxN3OFnIWtCnFuFZVbd2AwF2ToUDZmX5e
YbU6EPRAkPZQaszNP98O8Q5bJZ5oECU8nOKz8lQDX25gJ5Lun/jWpro/FcPEshdWMrpgoHPH+EAr
aMJsZBPBTCSA/M3LI1l8TljwXNarfixRS98s2d/odk+56RWufQq4xv03eKi4BaWoB/zSjvbpiZWI
+zNaaaLkDh8GG/CCCvwR3X/69A96szwNHxQq7/IYpsqIORh8tUXbL7R83Yi/xMCHLxKtSNfLRb2r
GW5CZFRkAYwmAkIoK3yjD1+jz7ePD2dqAAy3uRs3M5nPt7ZL/lhwla8xJufUt4E1q3gr9BlUPWLf
VQ5rT0IwcVE5ZHQM8rkfeY0Kkj1gdRLzhuBjQ8zWWPx8M0uWZhiJeGDyaUHmzAyg4R3JYuTDIoH6
btt3tOF3wY9JcbP23cDsCUTSYs4HzKs98DtqdPt5Zf5Qi+RZguEOAHc3W9OaMWeMphQpbwVnBq7Y
8pFpA/tYZ9pe9ILyd1PFVqycNUd1fFmLnPXYzCtJay5jxV6Y4WMI7hCueUc0MFRK7AuPTHVC1933
Sdco50uIq2zDl/5MVSb3yHOFEbAGYfmKs8iDLMpk2FzZcR9IeaLCHtxJWF5hQzjZEb70G42OrI5c
OicWwFTicDmup/DrkmuOQ3qEdThKFArFjXEvXuABSBb/hJaxhhqD7ZNUbq9VJ84UpVv6pzfDpJki
eN4ZSBQzn4Mwou/CQziEvQorEIeiKok+izIum6e+xfbyPOeuzPgxutHsJdoDaCsPomel4s1yaJvx
uydIEejPFNSPMDWFh9FG4JZS7m534Dtin1enjDgOPzCwWdf4X8sKyE1Pgktx/yxHkKLb1C1x2Jck
YW3jtfu4JxEal0OEOBLYL1eZKIy3MczUiWGFOinaIZIKTqtUdrnkhI8Y1KcwVaaBY0AC3bg8+yLZ
X8Zjt/6J2QB2l18NkDjG4qh/mBZk+VFbrdNbrpUmVYccRTRyElCAu1CI+3BOIhqLIUYy5nzEz4Bd
gvkBKZbnramz6meYQmTG+bFRTk+NCV8ps9SwF+Of0gBrOHJa2uSVlE9HpSRNQsGYbdRhsCpW1jAl
fo/JseQ3S4rYKqEAM3nMFM/0ZMaOIaV4vJH3K/DYTscrkjwkuxJEUIwu5haPxdTGFNOrZl7u/WIv
tDUjh25cnDqfKjTIq6MkusOiCmjSYr6JnTZYAk10KHZlwyuf9NSQe+TorAY0gQk2vrdLpuZdol70
mSbOAyuGHrBf5ab9e4h3pp8789mCpd1MCKNFZneVR6B2sBThPAEb0gUYka9IgqxFZFVvX2MYfhwm
+BosbMP71Vh25FmNY2RkTxb2F3yMf6eTEVnvIkL8NQhzkK9ihEWr+rutXmD330EZAzqOShGETiEh
uarrr91sr3WwThg0MbrCC1QielCkicTCoJ8XJyAG+uuYjvOFp4CJTDiLaE8SnIYbDkPVyehKFlgA
+YkeK6oDWaBKOEasa63x8h/03U6QfdL3SLq6sHn2hxPWjQj5hwFePifaxJUDfnmcrshidXgEe5kT
Wf9s0Y8LWPFD3T2lUAYALCiL6y1OTXOGb3DLxJ1XtfySl/NWpNjpulFZZN3/Rzdce75m+/3I1OVd
FGGR2zVO0E+jPD5DyXlv/GYVbUyyYi2uzFx8OmP5i+QFnWLonBLIHg7vzM2Js2e/t9YR71mmNlFP
Qd3xTYR0GyTFnUlDVRTVl8dnwXzPwa53CdOqbG6i1pjHHdsN+JcUYDSwdylb2SWM8j/T7zSAMPQT
5KBJ83ODhB93AalTiK7E1zjPuMAAXAKH8CGnGNaJL7zc+XYnPABYJiJ3YptF2jO8KxLxYA7o+YCi
MRL9FHaiZBytfJYapwEFYO0igAOfbFLWj/9ESGz/0cbVNrq0PRtFS0YOu7CNoq0OCfjSJhKUOAfN
r1QhGvboAi0F1Cu5tfYK9SHkOeO9uefsyg6okSR/jZgUFc8Qkok7+idnwrBeM+TUXN6JaJzg99aT
QAth6i6t21J/+FPhTKrQPTiv961tOMYKlIfD/myWGpmbS0JQHcWyxxv0w278cllDJ17dLR4vXs3W
rIxmRgrOK/jnsBR8FgK7h+vIZKHwDRnHWNPCtVqZa8srUEZDZjpX0ChsmJ0BODlzz83J2DlUyN1+
R8SvBbjj7YEmFKiXdhBxwKEHOo/Af5XwoyelpsyS1hz54yDRo5PV+F8ZCAk9oluijV9vb4d7/TLY
Hf3t6F1hf4U7baNWa1ktJeM/y+FB6icBO4ULpOaueAClDKRcM0bF2Qub/beGhdaqDhwDT2FI2bpg
DFromzShgPW0Ux2cKp1iMk6b7WRT8SwQD33lMQ5W6tHjpZo2XYy0uW+SafzEsDfy2atUe3L7Pc+i
4A1NSQOsyVqUx3idVyKp7uEx6sUWZFrJZoWiceK8T4kI0EwSyNjKtymuGB83bACBq6+4x1PRtTxM
xM1wz7UjAnCco4Ly414AlYZXadvRAFNCTw4RYrxNJv4jBrbzfEkUrNTAuldAJWl7NMsA6uZmaOPl
gMqIke7lY7d4p0ClNKzQWfBFvk67fx0WoZQ6i3zruG/hC4b78zRbSPjIQlR5psyyzgtOXNMQ29rj
CUBUAp1tOqC9pvTSU+iaZDI8sctTbQxmmGoZLJb9SboAbw8Hgk1WHj9I4osnLjjyWp+zE/qVXEvf
Kbe2yNltJEmshjDC4cLmd+pbGvChIaggUM4qTit9GUhBPkIOVARoQNc/jlBu+KM3ys8VhCQBKPOq
d2BN5DFKG7o4oAkQaUVbPqZI5Ccdvhx9IRqQ9A+5bAX1eZiygbKDZWxgHiZbXfrq3pIAXC8CC097
AUEuW2huIDDjjWpMiP9kTPChRjAqzsMRZkzuqO0vb0tzPBpmycoM6hv1hX73hBUUOjjtCQ+S9t+f
Bo/s0OG1vXNZzfglWhdkX7FS7XoqNMtYUEXC682aIGZEF+NuXNWgBbkrPGZwA7MDlVgnYWx4Qkxd
21V7MB9L87uIHgtK/Nw0AB3xDWgr0awFDv0pvjzrhJxnuJZax1sSjd7dmMCz8XxOUIJmZDTby0qJ
3jAxCuUK1gagggEeheZ8MJYxPkU4/bUbX5SwZo0RgqodzISZo69qiSVvR13MVKehRNWJCxi2bWn4
vg/LeFMNi3Sh/JPY1slEb/vc2lfYIIZQeEJuzX2kSSmO5yZDoQ+EA0IKnorEeFzLp1LtfPMsC+p1
EMxpamGJB3GSPmLrV8EyI+R18RTbl/NziyWB8a3ijyFskwQ1o+OejMSx4sg70LCxj9oocDkkE1yZ
t/THVOuUh3MmZjc0P0exSMlTVq8S0txOEZWjmYW90YpdQRk0YFlp+7Z+tATaYj86gvJRtXEx0Pwe
FzRP+1mqBWh1dZaimztXLulS5mV234tFanDkobn5lAPEJb4Tm1VXQpMiA7GlC1blpF5X6gAc7N0T
4kuwbHUCyhP/dEvsBEwaDMppNuqapDqnKifmBM3pCKFltIXcfXmR9sERhMrH3V5dS908ubiQa64Q
13ymQ0t80dHeh8buKEXPA439Zn4plq7n+jP0Vp49ywti6eRcDkoQ5cjLzU2c4U35pfrMF13n04QQ
aQG0iti/LzVGWRcgoyPlSaLI74GyLitPpG4/WN9c+KZtnj86LMUj3Vmdk7fGXh2ICuZdpN10V1iQ
SR8TPznjbzhUJT6vu5aBZVzYicLoENtDAF470o+Gci9s7+nPeZJSCpFWnUf2zObHlAbLY0VBBEEr
AVL6ZVT3KGSyIRpBokG7ZDU7Q+CQzKwn4TyTfBAnElcdA11qxKKvRW77sVbxvBDjTBADhCUouUg9
Gt5fdGlumWnebFFNl8FzPu7FqjHsfk2O5P7YphP4n0Q1sjU57Az2n6muFkKtjY/pjRb2qzNEEoNe
j+Q8IUxC7H7DSvLB5Y3jbqWUYUcf3nYkV6Anf7w7tG71X0/w67oF9Z6f5dlcdJlr0UcH9dAvbaO4
ewFDaSvI1/Go3UoO49ld5ZVkgxxplF//4EH+rQ/SSXx8YsLILZUrT9feS46Ly1xkUhJVJS9JUBzP
KdFvXhYuB5STGKYmxOxTrJpEpr/mVX50gqzZ1i15O78JBUUcLhGnHWSTdlrTUOuifZsJbxEIQZXc
4vLm8uZuTTVIhzNU0DP0+NS/wSA8oDGWWLmlLxpsz5fU9HdFenJdyj4jhdTQkA+dk/2cZmYS5xcj
3kS+pdtk0VWgk+ueGKQg+OKfYGXEUghCkqIFc0i5JZ/i/W0OLPyOqf3NnlgkjuptUecPkhypUG3P
j/3dg9GSl4dDLSEVx7WkLR4xKlnvdLDReHbrXRDQPsVspWh08Tywa+WUbQY40jUXIAu0gNbZQOJR
fQorl/FchtlAMqt2QAKCXZV6nyHmuBdebmakGbCAFkKEsv5Rl5JhLACZWK9D16J5NV4I713Sv1Ry
JUCfTt12iqWL0qBboEt/743PFO0h/8PGiLipbvT/pB2UmCAui5bsnN/4zBP2+KLdrHxvsd7vStSo
A/7i1WrGPYWt0y0Ht3sWH3bIQXs7HEWlpeH3FLz9ea4K55SsyAqAfva5D6zuKFXiLDk+aaP3G0Kr
M2z5vzqrvNqC4zFnwE+mJ22iotAPj+vMo6VC3DV5yYKUh0BN/yEDzAVZCj0ix7ugo9fzPS1RGuZ3
a7fhyyGYrtJ8k2oYL9fiGF19TJIXm9rwUzPdDhrQviiRAQ8mQ5On9BnjYNmmZD0nUDQu3uVyX7Eq
0Hh4duC8eOw4dBOX4r42rXYVG76hJyr4QPv2PUfuYTXQeo2a3a7dpUiNBWgW5raHX7whPJ1heJ0U
85NTefHT7agsbjVttCgwyPF1BtIQGsHcsI9rhE5codXWExs+T9W3gNpQYyaJPvHAvcbjmX/4O1GY
n27seNoYiqCntkyKjUaaqDjLsJWx7Rj3/7pawYaJsRuGmyiLqodFcNwa/yS8tyiRsKZ/3GqdTSqr
P4dLxbluxwzcFybMB7AzAjNg2BGlTYUpV7ivmWJxG0R8vV7k1m6ARxqu6y0o7pOct8j55uytcD8y
xtgwYW49p+Xmiv96OyQCG7J1s5b7dPQCycfQP3ZFelbHL+ncNTyrnhdmYK/604CB1asuZiMrxHjQ
xMGXfeuZuj0/Fs0Fc/DcJoqW4fDx7ZJElgcMELCtR3RBxSrO5+FH+eZq48AjQ0ZvhBSN1AGwyVyK
4H5l/GFc3i8ONprSvV/S5+AcpNjiIZeMIP7X3RCbX5Kz9uQVxvyrRK1JYXBUZuCn/NmuvQ1ATZDb
WmOH1XQGOFZoKP1hC/oDesOSbMESBvLIYQplNat4LwZjYBq5giQi+JQ2JtJRY15t/FJgHKOdCHZ1
GTi4h7oilpOdIQ3uqDJUk0cuqJQ4Znyq9AlYwTUbTNzYnfqofYUAbmaTZuHbMxh2xzINAe8+Pec7
po4K1xVW1/9QifTV8AIQddd1vlfuZVUXjYVLIOfF50ap0dLJSbq7oq2eAiXahGwqjnDIqJdk+NeY
TCYSnO4AbjFqVk1gZW2K30FPdeohi05VF7AnHCBPoCpmul2pZd81S9sGEXBoIUhryV3QA0BCLzCV
j8+KeahgU+c7QjiCRekn+Pv/37LLVRroncr5fHCgc+vIWkGMwx/PKV6fo8+ZOAYCP9H9atUR3lN6
I3sXhhUXg2y2Xv+TwWU+j7wfHIRATATaEOO+xPwLz0eryJzN9/fhR8KA9c7+CbL8KVTEKVL8eiGe
/ixgrdkrufFzJaHUDeuJxOIaiX+JLk8DLQbMx8AoDHe0GP81O35udNCrs0p68v4iyN5uUhm7ISTK
Cw8/RW/46QNBzwYnlL/NKClkmR3eu4NhB2nkeSdDWYar0GyHlm4WyyHEVn6km2gJBqv8yWRQu27Q
wT7TJGEZ7cMBbbspypNiFYlaLXb187+DpzbGDRFQcyuKwTjdx0dGilxi4h5wnWv1sL0HlPnYA9dQ
cRO6HcyP6SxO8JiLQ4YebzLsMo1XqbW8lmVmMNcDO7jaPeGrei+uhlESLQVQKiO/zdPTrDybc2B9
eB5j9UoeuXVzRoeLydgsGlpfgV0CCQrF2VS15WMHms5LL+/iU9dR7DCTuT4OFs+LPobTcK4duY3o
2V8DL2XwZ909sxNy/MGl1FTp0a5zUUWbbF5ggotXt7mc+HvbW49jKfjM8bsMbrNekip1sH4hMxUc
1l36HgiKRVfNz+EDfSqSkw0RLnNvGLYqyhub4+Eiv6kVrx6xIIs9s3j/b3Jqr8VZgz5rkqEDdB+E
ipU3NpFYsv1MQj+OTv6DjAAD7A/WgazQdFTAA3pJMb0++EONr9WNOXceDP9oiBlyBQiD5tptjnCE
RbydozXsFiYukwP3DjuEbWbK8GTByAJ4pu3M+FKEqtzTguKsX6LbbjV2+wiouoDEt43fzREtOuas
bpEHBJ6LMswtDGViEInULQqftmBXAut5Xj66pDgIrZod2ALKwkLmqFnNk76kGW2FHPGCVLuSt5fQ
y66aYlUkIPCY6ZWQ78IE8LUqtkCMV7OPRx3aEGc2MQ6Bam8NeoyWmLjQw+FCcir/DpJDvRCmo9ma
LmFrjKGxqHmepMmSfG22bPvDl9uwAW83QYhUIbWewZMKpKyVBpR88suSLwCrM42TMiF0m4Ty6unS
EBGLNlXyM5j78I9OlFA4orqq31PMoAsSDJ6ExiNaV8RmxiGtb9pyKMUKuxb8PBuwEkH8FLBkLQMC
pwm5m0fZ0czj42HNA1XaBwvv/zudH1lCNs6oMuvrke1YAv58AEbqolrhFf1fnITpturoxyC7RFyN
0SK4a+TSwH8cQtkPkzCpPJBTzvv+qL4ukUjVk+QEOZhHHhndY81NQkxptWN+w9n2KU4bq8AOk7fy
o0rttjSv5hXQFGqMu2JdZHWNVP9q6AHqyF9dq05Wcz1+CjkT0VpnLHd5dVJWNCZGWjtatNgsuss5
nou+uBhbKrAr7Jk8vmH578JMRUf/miJ9PQLvtBI0a/20GoJTBe+s7HCqDP5idzrlfnMi0AZ8Up6R
SC1laqqfcFAHmNYpza8AKDXuQc90GqAQZdBgNsFRbipXLgxmLTf+fkXp9FuLPpc2zpmSXPGfwDm8
TKIEGq6THl9ELtKXvnESKf2zZot2meNM6tiNEF5mqJnpsIx6+7Tk6KVwbLwsSI6qca8uWcFDm9qo
IoPd99BIyHsZolGeAYCW0DlLwGjhhNM6IQwZUdgW9He11kliS7cjwhSBYL92RDSklY3SnlssMJr4
seii9yiBZOD3LvajSwCLJjHIaBkM0wfi9Z2LSC3JSjSdDXEvQl9mthiVkYHcrS3NyICJ3SgBRXQc
fUKfOKPJKsuO5S5uQoC4sjZZTPjkk3Gjk8L9v2O84X4SE7CME3VtAQYH+fT8rx63cVVT3F71JWUL
YseKwiNjE80tlAOT6Bns4ABUYmPBfcJ/DRtW1wG4leNx57f9p27Wiy7JFEROwO3t297dmbCzmdP3
wZ0y+bmvzGpSqmGSDGKHWnfha/jaxM94D5Jrwbh/HoyJaBVhkStwOcbL7uJssQeVkSRTUlWbAcXn
0kPUPM7fE9QOK/8ugx9ZypKO4MOAvqD2uj3yvrjjxc8nzQuNKO5Bnlc5Yh/aUBUMa1Ng6zDf+RC5
+Vc21LmQrn5WqBYmkVFlaKIP8oPMavnqnflMtAP8N2soV7QRqllg88hXQM/x3gydt6Z4LQXa8wq1
JyDTUxXbtV/99H+Xp3EZDdyE4BUvjZlr0leQUeQuDFIkm52MROuW6nuw118VFmXmeOnLzJ9dmVbO
c0khPPGs/PW5tjB0joSVg8/1qYmRpzNkJ8WNod68GEHJJwpvtXf0i3oT5C1RpgNAC3TD0XdJQ/rS
aVxMS23nQ6y+IYcE4eBrPgHV6AS2r1HvkbksYcLKSUkD6QaEUtnd4hje7LQSzAcu+hIuLxbf3/Uc
nLKXvpGZNxr8cpFFU4hycw53+pPSKLT7VwIeaXtinThmx0HkhUk4RLfvWHirhM70evk0uGazrh7B
LeUGngbt3NaIny5Po6WPHpnp4TVojgg6HvFeICjGwDeyuStBd7VnCVU/VgJ4llqgyT1OBpRRnCVE
YK3Fn4vVgdO4rQ1I5gpoN46Xe2OpZThByWwq6NjYK0xAnM/bj23YazL/AGlAVctVnEEwmnO9/dh8
y5aQOLw0K1H4zl0Hb+H+gjAaMwuPqu07IB8UJLoqa3Cu+YXWPbYjTNHLJHwtCynWnq0eu1BNZA+3
2cpZPkC197lmtBSBbQDU6wgUQuQqp/lFRHjVbqjYDHBMY68GErplqYf5/gsBhBXgQTKCu4XeNSiS
z5b+PwbecsBkHJrAGgVF/zuFlv38pmlMma2Nqn2iHc0KB17JtT7iod6Oax11ILFZac5PV2VcRBT2
vmsYQxSolFHeLwisKid0lQpYIou/PhOMvARgQD5cDBtUL8LPSasMcs/QA9NL1A+z7DEsZ8hlzvA5
K6oKh7gJH1Zjz2xi21Qt8ruWQMXs2/REPfvUfHHEQVT2rr2n1lrGJmA6vxGvZvbpRf5Kx3RiSOKm
o4xevvYVY29Kil+N0CnfCIg4I2g2uo/rHJm9YJj0D9t230XetyqzAzITc9hJa8oGDnbQvrDuiVJg
kh1XRyzGbiQxPse03P1SWTEfk32i9PVHKliz780CBzgZ+urRnonMO0ujjY8Ttj4DgCrU1WXhj/Gh
7S/ZGTmiTKapUl0OlLhyc4DiAi0VikU5o+rTTJx+XyySsrLAVs7sg8A1Cjoxf35WsHv/9waCPF8C
z/wHOv6J6Njl138mvhKelHLkcPZsURCIIc0273syVoc+84+/J/QqFEBnzCBizEaY4OIyoNNTZblJ
Vqi6EXXCfWSChv87NdWkl1E8sQ3vzi3gg02HcTAsXv2fqjFfC6f5HxVTrF0JOvenwSTf2zHZqh/G
vDEQwHmYFb3m5B2j34K5mYevKjzbML5uMqYTWqht3HLAT2wdvWj1cye/TIwy5LODsdNuejo5r6L/
XpeppxbymeHlyfc/BCu/Rsrt3pDWLMS0t/YUddGVdRynfnS7xoEd3iCE0eki/t3E1QrZhQEfINPa
i57RIvYeiqWo/xZpsr4FHthY2oqoBIau21gykUdeibnNKMC8nSLSKOX8mXSgjqeMIrcrbRozgBbC
xDiRsV55Dcb6ktkB12JPzAKZFVWaMvnZFPUZqaqG63zwmKp4BzQPiMRLHgT5gMGk9ldEHZ1h5CYO
ZQ+fe8pdskoVL45DNLaZhzB6ps5WMz6R7VHN1SnATDHSXnW2b0WUQmPaROyNA+mb+2mEAYue2pD3
Yn9XJIeiylRlf204dH4JT3p6765cuLLrzAAWINk2z/pvbWvemPm/JOSdiddW3F6ZuCSaweF8G7Yu
jvPIpfnZHp3w2cWyygT7jYYsO16FBKKquC5CfcILaIjldf0hgAkcY+ufL50DThLeOpqL1nFWCI98
ExHi+f+bN0B6fa3o3/Jd6kGTD9HY/ykkKp64MN/6Z1Lb1oNx1dxvLbvZ1AlcYGxSjuq7R0ZnHv8u
l18JLTszu5XvHSZIYi42I1XqAQ8XUlswBXPjQj8NUnT3lQJoUsQ8i7O0GYXUdjgCzFijDRwdfCev
lMULQDUs73fw+zSyZy+XJUitpH6/30MQ+Q2F//pOLTr+UF3B63FVNzZRs2CSKOPUjjDkxIhW+4GI
pqwodHvHg97YosXydddqeHxNqSJ5FE6ls1VE0/0FjhvHmgP4k11/ulH5qETqPuzoB5jkBDmy01CG
l5+FASPzU6nlZcxwHbNuArmNKRZN0sq3UQ0KRTjW5Qv/ZMojj7HWEJyw2k0oRkYN8EtW03w9oiMJ
dMm3QaD2YBkWuCkUWxX9A43H5bw0BwwmnFCXfeboLwGW9BgSwJeE84kZSM/l9ujoOutRoWxxXJLm
4vFmRyLB+J41eT4wp4krcQgxQdlUNI/lOjP+fdhnOvAJs+knBcrN0iP+qzWJ6hagI46hh84dRRaE
EN/LQnLBRDAR3Nabk7XwBe1i7N0FTVAMwJ84m9RttWenYk/KfMXtZ4c7554dhj6YtZR3WlCSIfNJ
VojSuArn9HCTVN3rjC/wrzweyV+vw6DHMsGq0h5YIQWh0ypKsSiiMpLzuE8j2dTqDga2J/K1fe3I
FHBjVdPQCQlBYMSy+H4Tz3qHwEaZ5jU/GbMfQrlXryXhK2u3f3duoajXlq1WNOoI2Mav7f6aUYYx
Lb/bhlmvsK3vxsd5OqHNnGsGEtqedJ2VSHtGUdRfDJAyRXAYmP9Y2PW/ABiXO3gK/vlB+3hOIO+8
ffqWRceEp7EVJdoqIqhF5MVoDic7udsxBqVqMuVPHd/WAi/ekGpXX4/VC5t0l0+A33oHJ+0riwX/
9ZJjo9q/4x0E4j+ycR2aATSTZ9+CUHVXMstmdD11Dh62wu9DGwsx1Xq3qsbNHeX8wRoW7o9WaU0H
jOa+WHx6o3+ARTjc0YjYvNtSAg3JVC1tLPlfn1O9v9E4kP0aXzCJUe5VyDAN6G175W1g731jGxMU
wHIXPuETnTz7D47UGK29/FRucykjr69k2chtzhZFLNM52lJIJ5pmQQOq48HkwSzdgs5y9we5ldiP
kxjQGrJTHNuZpy7YC7GDqYdZnda7nPL+ZqcxBJBzLc651QVU4bJjPub+qcTLt0t2u/m2Y3h6WqcN
YAIuL0eS/c40qM1YyzOuUc9lzsIMLoX8g5XnlrPadz04KWrd+fU67YLcvDEla5vcUf0FSgbaqKDZ
hmBgKnfhQ+Gem6cShfaqD++5mRWeohz3dbBb7izPtb1MwgfsGf8/PfHhWBbIDWok1lBzltQAfK8c
vFG1BtUn4EdPJaaPqwKQZk89QZ6xPfFYmlw8dRqve8PAghC3WHQPnJzO2TwpZvgDXPqONt6y6TTQ
y+iPdmCGKQvHo83sfrJkMPlPAX07BORmaahZqHv6egVzXpqcSl/f4pg15LfmdOGbVTQ+/OJldKim
ls0NNfeaRdGa5cO+PV5diwGgozr6LkBwM7VdGpIae//fjYUzh+hhNzvWJJukLpowb+nzOWk58cZN
mZk12X8tax+BnoRu/VaN57eN8UklIEjROI0QOfgxIaE3tGAbb0PLYU/Ki8BJhG1qVBlijUg45NL0
NapkJICpYKXPzPhpvVWsK1OonjHwYm7tr3uaNr5L7eSjaiGpSUDVZxqmBKPW8wDUz/ZXmU8tdZGT
KcWKQq/JQGUFQvv9WlmBtXbSyaeW5a7YPLWDSKPaVmhiSAzkUk+TZAt4TEFsggGs3HhdUE9KbviK
7iXkaKR/msB2bmlWPNFaBbcimpOgOKW0QoCqws+GWg9qj0FymeARbdZgPBlza5AX7YPo1zAWy0Pr
bh7ZLu1SQxiF1JS69ZS9FsWSWWz72EePsz2G5JRI+Vvw/oKARpuBT2rTaFbK8KU2caYIjAZj2b0G
YssOKE5/Kn5VgMCjVETEp315oh6gHkfK5AzcIAACyaHrp/G14Ybu8yIzrvpXA1MuIUDneUNbsSWC
XnXgfYpuBJhqzObkBjRIhHVJLRuE6f+Sc+4ylqMz9STCSWfxs+tLzmT43HIbNW9X9kOWs4rFk3qS
AtSCPU8gIVeRPJzeklzH6sC5z4o/m0BOVwaBE2b4zdlK+WjwH184vgf6r/lkxf/q98BKXBWbzxWy
WHC0h5YuQFvtM3A1XSS/lGwLdJFN8JnZNT/VfmOxN9Bh/YibxoPoY/clbdm7s9ftZiqTmrGQfNgT
AbdghkAadxPPLltIyEOPnJTQOXQqnPVGo9rJAA6uLE2DlAgH254rqcm+zeGlF2oCWIitWMlqhGlR
SaaR1G9gwT/Jnq9ykxJI3PXrBy3mtgU3S18sYbbPKQsxN/fqt+FXrS4fT6jgaSjfBqYRkoh95hIQ
QKelGDQ15fOGxEspLoKeXCvV5YEaRdY/+sVZPZpCylU1zoU9Jaoj3Rhb/7MjrtgO5SOl49gSzNl0
LxhKCmG370amcfQ3vabk/Fr1qIOcVV6/uDxgyJ0J5irHrYWGo1yXfrKX/coCFbk/zvs5hity7Hp/
lkvwNa2Qwp5X6Xcu7eHSyx7OZOQ8ulif48Kzs2+fpqFLFZFirUsMTPhcV0qMe2tfp98TGQKEI0yY
53+fItGfKL1Gb1onz3vjlGDq9u63/zTY8keXjKp/L8q4yOOaaMznopbPugJKu4lORj76nsbbJPcS
e76OhDHLKXoFGRZ9tzYsbwdpRwvsmHsPR35SmDISa51FDEW8jCySlESRg3I5EF9lHFgb+kqBv/+n
5HwqWphTsaprnKaks4wsj46332YO5RLkhlE6ZB/n9IuNTn6YtqIqBMtNjM4NTKAv8+6RRNrozPcB
eRwAlO9usl6q7iOdEZwa7R8Em5HCbX4aYO30j63bojhwk0J0QwN4zRWzub90UzzKE+QmOLlVpoIm
spGaqMFugXJckn2bIlbayJu8yE9/yZ38P4VSDjmOFMc2d3dtb7KI9V+WGNY9gAb56mrizRlTg89e
8PlmV9e0Y7nuChXZbMU9D5m0PDKNFuDleQAOkjIob5Y1AR0XiRt1OoKTMqF/WdY5qzAgb3BVGeI6
6b7QW+reVB6sqcPWvM6EguhSb48C7eAJjodNk4B3Oqx8ibj01B1Pkf6HYHOdUmw8Wx87PwbOIGip
XrGMRPSjcICnx/NGz04GtwkJY1Yg1yC75OSPgLRx/JdcsCLm52/uxgUlG/yLiRnk2WpAfFGgbcGV
ui1RHYyncPU85xO3cc2iQ8LdVFiw1GdhdQ4opPEjLBGyWox8/G1SIMbPySmrKOKaXcCK32DPDdbB
1nOW0ZjjBL723napicvn/KPk4vJwoGDSZHrQ7yEYhYIaWUyMHiOzSoXspS57SH8KE0xv8ra1+xnY
Sm128wb4D8pRLnE/eozsNZgfAZ94H4FX5eIqpD+g2kG3QATt6vsz8tcmJ7C3ruEhX7db71Esx6/E
hZ6UniZ4IYoL0RIGJqbeY36DzPhh22cJBVgue+psUZYVQ96TCO8+bxREDEIHZ7ryLMiHsGQow0DO
9jSCsGCe7yEzXbb5eg2ABg+pjiCNrH68zzWlt7/7RgwdQDbKCs7yDviBNFlNDNsTsdk6ikLFwrAf
odsCiYEIzOaEV4/q3q6fAMbAn/uwQmAxt96kywfj36uIEFX6mZEk/7W8u3oQG9aKLCdOsP0V1Qjp
arJAXEHA9BaRvFOHrquRoL4KAQ1P0VxqVMA9F2H0Lr8sIQ0rP3jtUlbapqXUnVzx9olaJgfBS90v
2s1Oy0CUMdSqAq3SBQHKW4d40in9y9UCaFmPFbP3aIMTha7ryOGjNX+5I3TP22bjKpC8RKNh9FhW
8CZCSCiOUl/HBOOrW+vORE41aVjx1CZ7Ei+Z7vKRPfagiKaawJ/wvBWFt0hSOSL/vlYd7nj6aJhO
cemVOIraj6WKTiJCuMMtYFMnwwXv1K8imAXTXQRWBAT+9rN2JQFG0Q9//CmRrIn/6LjhRGuq8Hxy
em8/A1shztEkUeIQ0pBHKtHJEheELy7sb23xDZXdal4SsjQG24ZcOfBK7UcVkjynkvgvL7Xil3UR
0a3hnC6HTI6DDNg8v2nykGqKGR9TnbUUMGoQXHc3/AdIkKbGhubP9CsD6lPIGHqvm0qnPFQH4GWh
Fj0LbFsYA+J+0Be01pHVzEOi4mfkTHcW1dipWDKV4xjdeRmicxP3Qjoq0+TEN/Don8qaJBisJ7mY
mWQJriodmKDxVh2cccFyPyl4eGLtXwuWuKY1zwSObrn+5pla1qPftYETooZu2bLZTBRVT4jijfP0
UCer3LZzx1XTuoZaUQXdMydSVlvJIjNbcSljlh4be2uqpVFLmCYgk7irDMMD9/IecbmVYYOkVd1/
r/RXGWkTa+gA9DcAd/YhUaoPKRfollrNmV32FROGfpffMAkLGFsub59pEShzIbe/vGQ0D+I2ewRs
t7+c/hXDpckMtbxLDeGs5lHICudpPUN7Wu7NO2sFA2EJHFrqtoQmvCZAGA4qqzUU0xLwtKINga+J
q/cPFtisnENxwCcyNeh864ZxNhm3Gljpr8mdWk3u6PYfZoJ2yIJk1EOVrEQLyEhEqRwU03cqRTUc
9ZytMs0kPnmK00e1R+yYjppptmtxPjkrb+tAgUCn//TQatOG+HVDKPXc3VIAw04x2+Kdonz+7+mt
uUkr2FuuED4jeANv7Z336tSJr3ys3nGYZOJdBnlZIZps3w4rnbNI1n7dedT63qYN4qeSCXyYXUCo
CFUetn6AGY26uopBLljwsivAIjmmfYNNxmq/ySffIPzE6+yLgq6kNorvYi7uzzFwio6aoeAc3abF
g72NliqesFQ9+k/LtWEXClDZ1tzaX2CakbmqnSHupEFiVI1Y72MKecfyQlDkXb7sLwJIZbbEc6Xx
0i4LeBDc5bmXqDNRWqrUGFjHIkgjwVbuvo2kudWrxKB+yn9lHlVUYPmK09zEibiAmCXPMsQ4WlOk
h/4kj86q6eHpjtqBGAGDmzafbj976GMazkfGV5tSSYfhemB6EUB1vep2OYZPjSKTKGS642xXYaHc
IWXyaK3SlKY2xtguvPWZpNl9eequNn+VcqcQq/f4iEKwq5YjbSgBvgBq/T9F0AqkHSrgknhfjCYg
OnjLL8vUlFxg7U1QvkpIvgsFceGD4+A4aXpw+HXYxvIgFr9f7vUZjpvQhvvaP2Zj3giL9/t0bI66
CNVg5ZyxM/mmXK4xSalDmXhiw8bccfuim732HH7WNH0rMA7U5tYxaYGQj8wJxwFTk9Xjpm2mko27
rXV5F6zxljKCUsNhxIEwV0hVrC9bcsOpF5M57EsW6OJGzd+kq/bzdC240Gqf3aJh2AHb+rW03ukQ
ORrx+SMbb2QLd6q1YSFkIGj3qP8JRYpb97tC1B5w6M7ED+L/ubgkBPVqQDrNlP5HB1IQb4Ash7F4
w2TtVE5x7wRLM9IyRrJiZ9avSMCwwRsvm2JVAcaIMrQodEgP7+Ud0SjeVCToq34ZIFDJpIKhf0LU
3dIVGzo1hxNsqhrPYOkrKbmEWldeyhzVg+/kFrBi88a7hIXuive1EW2SwMIREz/kpFcW7YGaTGgw
RV2ejw53kLvve4QKQWhswQqQge+yPI2HyiDIXXRP94c9LV7PJXNbmgpMgZAPjj8eMjYLXRWKqgnv
cWRSd14V7SZGC4vVcDvlPnhFhhkUr4gXVjj7oqnchAWLHP6QKS4rTJMk75DGbNI4w7+ql9la1fjO
ygoU9eYB9EXM5MJ+qgJRm8uBdyNxHYyIDF0LN2Fy5KKItKRjyr9uPPhZyaglGGH9pAMzoE4cNO+4
ZmToNMrFdBHA01tLlk6mazK2aB49Vw/8magMKCXtrlNaJZ7ShBLUpcyJtXSsbn+qFJKV/LtCSPfL
BWY78fns9VVRjhx6UzhpGvn6CjvtIs9UbF2/cfjAF3W06Ish8WSiX5EkovCE/hNz3Pr5zFOOlmge
c1UnCOqigO6HmX5Dw0o3PxDhkTPFtPsubMACye3b3Sqj1yKuw1r+Ai6llZ7SYqTN+E/Ew+g3K1g5
nOZh9gX1GUlIIirTbV9D57wzlsbuJyTM8IL5hjqqvBh0BgxjBkebFw0TvL2R+nJjMSvDs2GfukeV
5lhlndB20zQZVsdef8uCA5kDpAEaDJPaeIifZVU4QrxMDj3za/cHqXRdgxH3cgpv3uXKa4Gn3Bmq
DfdQNmZFTDKT7nyiQgdysHD4JnjBmCU5umb49wX/V4EYOQq+7VpPlTjduiZHVX25xaoj+MAo681f
7DePqnw+oxPQQC34m/1CGEzz+/esfvr6lPbpiQSCjGFpJKO7Of9Jr6l3TQ6i3/8nEoTVp4ADbCYB
y3oZ9LVJTBF1S5IFxp+/f0fEqk0Vh324YLCRPMVu1u33F5I4yw6ssdgIeSp8nHyIxMYx3F5KhYYz
N0efRr1rsCIUNT8c6HYFhUj8mz43e7LJ6NOakcIoUIQ+A9LRwYGKan+K23HKwcIG3hOZdeWHhpoV
WGKdI090ZrGStobOpcInaY/IeNygIjBaD5Z2OHODFfIph/7NsbOJ2/daxhWHh5OUU68O1W/w3Dsx
ITtzcLai5tOBG3YLvAMgkZ2+iM0fIwEuV+A/k0xw70wzpruXmJVje7HAhjTphxpc/BRxTLHu/J0u
CZvcQmqPHdRJboKgOxhbog5afg2Zs8k4qAvJ30LUsQZhXT8LY5VSVJoQYk5zIS7cAF4n31svxd6O
9uNKujwa35OG+NyZhjBYSGzOtkHVrenYwzxCH+tJwBpHgdP3OffOqw+dl1P6bULNdrL0v1oYoa3G
foYEWjO3cMFYsz8qquGTLUUDkWTHXSNFdpEzTo73djDc+XvxeMrjSaqDHtSoO6eU6EyFuDVhAyvB
YnP3UVjWVuhr3dXVv/cAI0jeoF9NOqnyzeWgSAN6FdNhjgC146jksK/tHKJgc/w0U74j1Dk73HWg
KPvIIJ7hhq7YFPfTZy+wZvoLG+MPimd7ktaJAKnTl98LbzIVZKSaVnhmrGvAB3/zXWTZIPABz/mb
4s9hX2z1LVffEKsNUGyHjuNB53oSLx+yg0JKC355POtx1UgUgri9+UL/rae6227t/C/iO7gSkbO+
eaAT3+jjXYVyeiCbWOHQ8KTC4Ha/H9xYXVx1R3ndUw/l8PKkG0aPsCLX7VJq9TH3zvSRvcvAPtuy
PFIrQYFdryzEI00sYZERQDxcic0Z82ajmxXfbgshJS1U7iIwnHlqhVcmxuWTyUDb66OydbjUP2vZ
0jER9fxvoQcVVvpnYlxexS4IVV7OMZvPc9IKFi5Ij6lptLWe0tL5HMu8ZX6SEcMiSu7Hi3d3cqCU
+lcDIBJHw+mWUPWp1NPnWBAQoGIZvG8cF6NugniEqeBfSLeq93xP6RJTep278Pz3sPdaEUTTu+E/
4jPLWheok9i7FLUcnEm1/kwExhJ+zD8rdxhWUf2nuFJW5PbECYPpzePIT0Zq1pyIF3AnLh0G5vsg
fdhYwzrKMC8UQRn3Lq4xhFL/XfjAX/liTWkjQErBJAvhKVskxwne9s1f9B8cCRIdkhcBijQdkf4+
64JT5zHFY6O0fOBb4C+S62VJ//S4jteDS1hnOu5aEPo+IxvBv3AqW4lZ1XVhWuQVZ2es5YhI2s+Q
5FW7QRCmkthgCAZzt5uLqxqOPhzqmCmWslenw+n1UM//UJhF1OimTYwT62HZTSKxsck3R3Dw0LrO
yOYsALv9x9UAPCxv8bmcr9e/ZnyTZQwk6NvBC6Q1yje+kCl36nMzZ5Oeevwm+bqjzxQHrKRU25f5
IvZ5QvbEz1DFM86XUF1Nigsu4agGukk1vTvHBTPsdtImFjxNuBeOtBzx3fafF15n2s+C7D5U1Vkl
/2NVPPZzT6RCgZnQQSyr9XME9mofvY3+0WHu9FMtJ/mVGcs7t8HIxc2StBSDzuRMwDsmvZnmgphB
acCCV4+6wbZJmV+OlnMYPjOVbzTkZAQ6kUCpXWFbETXCKgV9gOCWRfJWvvBkKaQiS3rEPDDoJOO4
lRXob5dMozTIyGpXC94007nZ+TD7N6fgvk+rpjvfD77GLUFhsuFWRtCTkzMEPTkwFofk7XhTP7bH
KQFEpYGBKphLjo34m7WxvS2OW89DGkbcqWcHu+5W8CbRn0tAq7pKTQRmDLnyQB2h/iKKk8bGLLad
gOXJg3n8xETpMk0DmBRusVcOEuB2wm+L4nckViTILY5bg2gQJW5PK7joJALfS+pI6ZF8j59bAmd0
q0WzzYzUwjCzqeV4pmvfh7t3jEmnoDTEULm0wsW/NwwMApSZf18XlSFsZAUXzVVLRPFfsy+qGWaF
oHqXM0tjP5xCM9zqo6pdAzRw4/iJuBBJOj3ocZEhYKp9gjmQFrwZ5HFV833V7ku0HgBMfXOI+xgp
+rHPC/6fmdZY6NbwaZccr44aKCXwQN6kaxb0/+/eFMnTgVLXt52WlDZbo310FO0E/362b1g+uT9e
mG9pV13lKjnK9JxPpAOlxWMVcreLNDVAcT8BAXcHImQIImU50wuQOoPysETxuqoTIrsGOc2lZnYx
7WMQKED/OEpOTQg4mGyHhMsj7M8JzoVUb/O7sicRJAiFrtLguS8r8N6szmFxCiv/m/RQFxx/eJRj
Cj+stpG2DvH17WojnQW5r3a5bJ3X9dm/GTMAGC29EDxum/azi96jIjxmxSq+t24g86/HbnC4jomj
oNoZgLERilwLYjdsy06kg6ShnkA8qWVW+BnolmWcxJDEOSJPX63gnwM26BN6fK15giwy14fvNcFb
tcogfu6+C9AH24knzbGM0liF+J3APD83cozlBKsz76xWmQ+4VQGmDFLUQVAzhre5MUzTLNK9Ap4n
yuZCHiCAsByknFvsgiW7og3N7d2SmY7xDfxajYcpzuzMnaeylJcKFr0iLMfEbroIkikEiTCi4xO0
xoBpsgXVcQIh9Ftag8SyVHOn7ET5ZvOuEr9RUkIYFSRVHS0vf34UJInmeCEooLm2caTtsNbh3YNi
/iY59LmX1EG6sle7qDFt6EmevUIJ3NsLSUu1SMc2zjG3l5BUwolOqRx9dRKfs56S4cxI3fb9LrTA
gudAXoUNIaWaPf2AxYLC3J1FyIywaRc8cxa3Rd2YrfD7VOe8s0w9ZU3CP4bdAnKP4fWohfsPJEz6
Kon8eDOSqi+gx3lCIqpy/TSlaJBLI0UJvRrJ/2Lwmv/uUokdThx8/puQa6lcrpuOnAa2H/xH2j3e
CF3+bVT20GiPR7gxuukSGbcyvlZx61RNQ4u4r2hGDrCL9JyYp0fMnklA94DiNs+TObnB4EaTBA1f
HJmT6zJkAq523fEH7ZWua+7QjiD9AG8L/uLiibrjyyvaWzUxHyRBHHfAtbRDJllAXvgmVSGHVsIH
wiMarQQaI3o8cCcdr9fHC+wFJUI4aVhrcYf8EZ+401ppbAUqGimqW93qopmH0uWOqVXkQhNt3SR6
o8O+c+r0GiBpLhmoM1sMCAzMltjM/nuiczwf8KsRNiEqvCG15GxaPMKfkYTzX6t/+JX1LM9OS+52
oXs1AARdRYAEQb39yp7V8T+MOJ59nD03bc2FE2dRaCEKZIF9Un6entFlFBsqzWe6dS3SVNe0Rw8z
p7ApRQGFIJC7HO1ZaI1h8kCy3cYCfoqclUvDBbwcetYAwDhZiV/svIUjwUAjH6wjUuAwD9nl4NSZ
sTTvBpSy2vaTULwVegi8SLht014CdhthpmvpWpBAwrXXwiFdzWdAZIv8qmQSD7PsULRfq55HEYaa
0n4HVYbwGD2WtlIyHcuN+041lMV94MwsyJSOqlKvXZvEpz7aA5nIEESRtlNx+TIfhV40Q8wjYAtf
pwmy9TwSJ01GdWR4oXtBRxmG1RCkoyMiqBSlikoYBYzlaDIAtrRIlONxOoA7in6xqsu3Rd3+oG7A
asfzFGBgyvIPBCzUgMA50NYiTxqp7tBKaPulDd5IGgPSinGvOxS59s8a7R62e0MqKvefmvoNZobB
F1qHBqY5uZL5sP7G2r+BrjVygq1WuVW+FejQUr/rRxcRaqDHkfqAZJmldpFfuZ8O0cNiE4V6xhwQ
BMc0lf61oSHvgxZNXqoIIADx1mG/AZWDI8cfSPSFJORwlS5lH1ylvvYIdE05quvfY6xD6l66mpXy
gWyuFY5kCCvOSo9AHCS4XRLqOSoGwZpdFROk3HDAXSpJiLrtGypMae6FHWJiGr/6vHh0AVlWKzVI
X9S9bLdg626JrcseHGO3tx9HRyjGHxZC51NtZ7LCTDOI0VDU5M5/3zRV2/61q33XtpVL+aY87hfW
1Z4V+2pP9FpmQOy0vLJ4Tu8EJek+67yWaEAhKuk8sbr53qC3D1Tj+2G0rUAZIaOz0LkMARG8IIs/
E+EZysRxecpZn4liiTH9JGSRHAmOhnoB4Z5NhnpysIxVJBr0K/1AlItewaQoTuJa/FBn3cx9ZDfV
5oL8309f0V1jfFzN1mlzYpqKmQ9SXYj1A2la+JJIMukwIiVhB94xWUz2r+n8yQ5l6DRUUeDXo/Ew
9FLEjNFmiJsgQtViAVbqTQS9G+mHCHgyy+mdeUSl+t38mqeQCnsn+SQZh/U5/JmQMK9x64PdX7a/
HWnEc73G5hXjs9rOUxlYqYTFm5g46VRQ+CYQNXCzajG7v+5cJKrfipQs43kNZn8ytmqP5bizKzNd
KPdfEm52FBgAUbRbdErnxBMoRkwwfeGt5OwBSHOX8BoSyFgSKZM7WcoX5TxOi3/ef1gegxI8y7EH
/tI22d9nqyXbsW2laIUtwJfW4E03tggYhgBdPRrBoJMl6c1ahKmxVsYIDyXhjawwlf7Sj1Ee84b1
mos1BeedmxsraygGR7ZhnDrgxkY/I7j+smzCVtBhV0evAZNnVTuvHiGu5jc8gTXL6WdCgcuBHvb1
aQzvnHV/EzBaTIgimOcb/7N2WcUcXVT/St5O4RFcsEGkG7CWYG4D0ORfJwMYEI031XerBZ9fZXar
ZlHAifmFbIT7WBDLV6RL2gY2cyrVNnc43gua9n/wZQx55lldKYU+As/ImQfaTGBLpBH7hNxrfXWM
RNohBjt8obALSslFh8qq/t3FEQSTbH4AU/e+SywDbTgbIQLcIa+KHE70MdKet1Y1uYqJlmvLQEMs
FgOkfjorv8YOHzopyyqlzR4FEqWgLgcKYtldVdjq8bbQb9kKnOIpQAdRJH0nkPbjGShYFrInRUBM
WvP186HnKMN8SS+r41itlmb3evQZpPHNTep0uXyJ5y2n3KyBdSVNKoIpDlGDoxXz4wvgUPErVtL2
SwwweWP1e5x4AeE8M/ibIj7UYjF45mEb2ODTGUnSnKgSaq2d10LDCoTg1brppVpzYCiYHERl2PFC
qWEDC2QEuNOF7/ZOrYlp8VHs7k9ZUBF6GHbkdBStJEDFoGuTtSbG4M30Ql36TmBp1PfLq6NnWdoy
rjZdKFUDnOuKIetdlAo2ycu6w7SdxEVfwZr/My+urJxPsY6q+iaMbNSJ8MkE5+uchKXjrjPXWG7g
VSbcMOhcubg9gRK5oEAftJlUR9w5UQc9e7sXsabGaVT2qwlpqe+iA7vel649Er8m2SLiFlFbyVQI
4tCOFGgDoIUzCx68XsBZ4RlSnYhPkMcg5eilC/IqB0dfm0dSSvikswUm2W/nlmYXXXg/7VW+PyCc
hpQskSJaNRO1q+8kZ2F6oUFMFiUAnTDaUKFYWbidKo6iirqiZP1/8SNa5ITBrrIy/rBaR0e2spOH
m6WpSbvX3zsysLr2yh2MLrPVk/CSoZ+10JpWiLTwlJTlKr0jBh0YkUbDRNizd5SNVsjfJ09BuQi/
paco1zlxWCCHarBqBvmpAGOad6rJQmm1eIAeSNYlmBNYDVeYk3bRTdtvizJ9I7dydsMqZZchcICV
peXg5617ZPfaCvjdcVwM31yebLoI62LDO7HNGWX3/AU3OF/0H8w2aBkP+o8aMcQgn3wU6mGQs9FN
BjiS0mnNy+VIo4geXEb+DHuFtCUYrvwEzlBnq168nxb0gTS5BFshpeQhMCOOi3XZx/wOitHcsthQ
OjAkUg24kT1AkwPf7crJWNrwJRjmEA3Cjet+3tmtARPOj2fRZchCY9zjnwr14BkUr69l/q/A6ECp
Rqa8vJJRzpxRa35/jsit9CS6mLiIznS+T3JHM1bEUxnGrqZgoYeMzimL42f1t+pJC3KBz7Gqp/AC
3JYJCwRaQyYex2hTNXKxy49AczVPC54q+IyJVWYnsf/zeT7cPRizq/8j++jHtfVOz7EPrPgBX0n2
UGac9SvzdXil716YS+n+vINzkOJ+aVx4hxjb21+jNR6S60wwqlJomE3A0LuaHXaqeFlTLBzgMynx
Mup4OXcHBj1Tod7BZmKybycI4eHfvpWqjatMHQ4Ra3wolrSZJHzF/kT5nBK9AGOaMbS0iZo7JEkL
T2FZOe7OZTW/nwGcsGg/E0T67uzoGSrtnHF+r/E57/ZGhk4Ee1dO0vrCRcCHXQFZcOg9u7Ur14XJ
60f7CvGbcKqfgKAjC5TK0VovL1MXHOJBS4j9UT3F3WOXgaTUXx5HmS6wfl9MdkWewB03kmbdz1NC
yVa/6mv2m/t5eFWmalZsMlwtltQ9fmcGLLaDoQl6XsWpS3D4foinGqyOvAgwL3MeEsuU+5YqxdgT
YRnvJ7dgSqFqxu90n5sfHbQCJ4K+ukUhIYc39J66Jybi6t4TnMKs8Blz6XO3qksS4bAjAFZbJhO6
8YxpGlzRJQyb9aNQCA9hfK21uPG7XgKewh9OO7Z5mo5Ci9N+LimYUx7ejqmRNYG2gkqkMsP4vvaD
ZBJJy6SQkJd0FR8GFBxb/NSPu6/nst9g1xKdDk1nkXrDBsXzkCS+igRYO/ScubPJaKcczTik6cjr
ASfV94JuShf2/q1Jj4tAI2gHpxR6CkMyPgp+HOyXPG4H9oboRGGbsZjC2grF0FySskwZei5BdTfo
l5BPGNGVBJHR07AiFoHocp80Vj2HWNbEZyorIH9BKYmedJOa5h2iK0w/l6QlsSafS9pnVz59nL+l
3sQpOgTlb2grkGy4+3b/8Pu/qTfHwsZN2/uOZ6EPQxgpaRm2LA2uxVwscplCbjzkKZISLcZFc61D
AnbYBTrG6RCm1ujW/HFq2PWB+eF7h8q0tqxwcwJDy0+afVpxApR94gEuR636SR8Xe9OxSDgWrqFt
r0oixv/VGQbco/xyX1WI3t6YEZ3sYr2IJyt008GCl8SnkD6d0MMZ7Uji++3ZyZScVAAG4/Kk2lXX
gYfHGcZluAqcy8lrJwb1Ogdzp4Yxr4k8CMDfpLf8e568sX+6rWE3SqV8TECWpvp+PfQN8PxddMA4
5rW8ka+k1174w5DMQJ2JQg38iDi/pkg1Dq51UwCgIlnxtyIgSyg72o21dYr/ouCPy9lqO/Qdnbgi
shJI3Ua5Jg1wpzSA6jTlUpveWTBlmo1kHMkIjtY6W8AuK9NQICPc9NqchVnG2Eo375HiB/24xiOr
zdB63lBYuR3Q2xdizo1MLeKp/yDL21e2uCJKkYDrQ8T9/xXhgAcPiRnzrmAjEwAC1kiW2RYKfRl7
GGRUxokKoc9bwNhB85zRBT6OwkHJeaMS0CRytXSDFyj/zV/AmJYercfw4gh+9MJftx2+efVtXS2Q
tzn5aitct/vK2onshFnaopJHcthayKho8WNnP07Jh9QWZgC1kQVQZZwrq0nwxJyb/BQ+wuylgOjl
FXft6klu40sEmXTZBXR5vAvUclBgEUJ9DADl2JqasCi27xHiwKNCZEyrU4o7MrR6CLM2vlCwaw8Y
BuaE0vR/rpZb3Qs5VhEKMNt/wr+jJpJIcWNP7gIfnXilfO9Fth1Mys5TvC2gizYMLlOvwcJv9isx
vP5e0O3688HG5ABYpD/QutS2w0vDKNJNf8Oj4yaOLx+imrMEHK1A+U6M4Nz7omXA/2iLY2g9/Lnn
CVSmJqsI3D0t5ofVUV1SMJ//1WKZnfxCjX+m4XIxkyew86xycIF3F6iOFxfODA0ZPMdfRTEC9qzY
8zenrsG1tUnIyNxxQ57rMldgWh8V8lXdGmuHA87xiL4A936wssJ4XVG3kDoHht2bvNPDfYdBkRpY
ZCQUt8eXzcogrTJH9VKuYnClGHhkM4/v/mAeET3yMlcSEpLN9MmAl4mDe7ng5/qqKKAHS21OTJV8
yvijI/3UcGhK+CncZOB8J7TMq6yDmCre26C0aoMpPMV5OuM3IxTVyo9NsivIv5X0ql/MlX8VmQ+V
n4d+QMj/+zeVLg4FOC2YJnQVYF0KYKNovm30rlgvV2dJ1JOTtmhFptr2uB4YWEwPLU8N3BWUsw6R
DXxwhgR5gEQMb1jpQuwSNVDt2RVgZn1hCVKTsUamt2ncjFchb4rJku9OWE5/GVBFhsdShEO4h5YQ
Lqp283ZFtVl/EIDK8TrqDor5+XgHCl3dP2bochCX77PoHzztXgUQfYc02cRvlnWGbjsQ1J3bDqly
/MLdu+3hrh/Vv5Gc/A2w/UidER2rv84pjbSon/f2B65CGx45uLPCGDnvp6djjwX0VcUbmU+Q2U93
aCz+hqf4gx3QjuOsfsMaFB4x4i+flCUeaiGRSbaoYwHsV1agQCr8Tz4jBdNngQ2Wj6L3JUh+VKyp
Ww6Ndrz342JOOvm5GeDA6LoIcHGgsW+ygZeKFlOQ6rp0IXrLtD37anMpC1TtoJaeBK5y+DSV5wgn
eHeK7RjcXjEGII4vVqKkj0UysEdT2kNcX0caykrZbkcPanUEP8yTbA73v5ImZz2i3DzcQrr9J1On
9uga4ludu9zN6BWNTd4e/20fWNoJW5k2V6fl9Az6d15szLwPjS2YVdRciAnv4OfZ3T6Ebq3GFzN+
MqvM8T1Ki0N5zWB2JwwIcW+VL04vRM9yDj173LLnIMGd61EH7GwFL91Oe2zt6rOThSqjk8YGtMnr
hovnX0f0wMTkfFzAFf2b9PlPFFWyelIhk2NlwYWGiEZhCgQququ3SfSLmdvq+1n88EarJE+6zCP7
LmiY/wmVu0D+/zg0EQrVJRnWE3U907IYfrmWq8GTa2rCVwHAGpqnpqzYvHsNonsAuW+D6kqXDOPT
cLlDfRhYbZJ16WlCWfQI5HsEdeZbfVk0EuMN4vVlFgSP7iwhOQrIErnxpF9Sx0NckXWzTY306gsW
V9jTNfYpjSMpCJwMnFzHo1vIznFN8z4f0/vL3TnyHRuvr4VV7rfo86brUtSLQtz8hCjQcnf+ipGx
lkkyD3yOqSftv0XPLn5q4u/SBqSDPltLAmz9WA0RLrIBTEvOxT/Ch8qKia2NmpPN8maARuErMPKi
UATnah9K3O5h3Zj6URG7N67WRKfmAwBtK4p3vFD9dEfIzjmpZxvPPbMB+Hl8qxJnsAtklGSBSsO0
5Ia2wQJ8WIRvHsosSR4ZzCf2/KEvas8ImM2UU9d3Nnupv1amET5/G39+oSG48JxKWo9Wsdit9PZK
BoVtKG/mopV6KVHx4WTNCcNPid2PtMclj+i5y+g2DrP3BrxqqbcM/9e++wqHsTFFxOGRjliinjnw
TT308w/X0IIseRHGqIVWbDQPfMGQY/x3n8TomCMaoFprb7QqQvf9V3e3d4Xj9vd6/0RagfkwdInH
adCuPPGLQd42KNnHrqDqDoRG4lFpOZVk4lQq5a9ckHnbT22M76o1u6WgL2QsHg2GiFMGjz1u2AdO
NnWwGOyHgg/9lWkLfnkU05tHNeV+zprhEdcK2kLUvAuV3cyl3j7rifHqEjEtn2uAdG/kKfWQOU48
KMmuPvrwxkmVUkg1FhaAEjy3a3ykkTAL+0b6tYrSsTJQ+HnGfF/HONewj1y/N6NIC5uF+PuTcZx+
DEAgJRgbmzDuHSud1mGDFTYZXUbWrf3ry5lT3HWfrvguJwDNu/FhVF8s3dY455SaH/GVqqD9eMQh
Nrpdt8IKDAs5NLb8TPh8ifFgfpaaqmh6HkMTnrFJXQvLEhAGvkickGaxHSVBbn5EXZ8Y606WIH6P
83hE3rfc8BJqqNSOWSxrytNUOOH4banFMpeBVh309t1TLiVnSjH8xf0kzFgP0E/hdhwxajcMK3Vg
PLuK4ZF2JUwBkbZA/JfHjBwNrtVAAK8dWA69jkOPNb08t3YoQSRRa7UcczpxSsfu2hxVd8LeF0HS
++dTByqCsRpMCTiMIwbZhOn3Uc1yNwq+T+iMh2KIdL/VJNQvlBpGyk0qvDflLMmEUqPxqTrkRZCg
32QFQ/sUVu2LpYHQde6FbciROLYhiALQ15Pw4pfWHJ1qbor5phsAZbal4y/lB4bioQQZkX4LzUus
KYc1GEzed6WZliu4HbhlG7njHWstmsU5jId0VTFy8dLVZYvQl9NuFXj/UrSXEr/Drnq32OV8//kB
RScYWdgNye3nxK0jVjB97J4xcXa05VA0Prr7JdXMf0pW3r2EqtVmClNLCtJY2KWxEiJgdq4ZEzBc
hEDQN/DjAFk2KaWFixMezvMq9i7F8+RxvFWiND2kmcAlt2rOdyvY+YVxbAnM1ZXvZRCJ7h0heaR7
fPpGjJ6JAub8Ty7wImHtyT2kNsFtOdZndqBY4jvxFqtWTHFnTM5wDWMixPf5vnuFY06bD3D7qT+A
UtGlVtiMt+p6XeNxEU3+g/PeTcdyDHqVaZ6WuJg4yEGeq/UZy3JHvz1H1X8YFL2Y55osQ94oORf/
DGATZ4a9s5eSPlyIzPDxmz2A0mZjMBVVs64Mg6bnv2Gxx7ITk14j8NMJ0Aj5z6RPskQzvQRFpnly
7kCqpaIqlH0RvUtB48XlXVlLWtk0r1BH65KkHkaAqpX5jj0fFYqmEk2BRt2aZu1WHSDPkcXM5Tst
u5F7U10Ke0wa61yiA26ypO2KCop4EANq0URzZV+8Ud3f/jWoqQyKN5T/grJ7+ECe05BoVGSHNwcY
+/ndFkvdFyATU+UzS0Am21gEhviJ5Sp3QIpSs9mTsXyPq3Y4j3O4I4Le5X8Bn1dtlRncd5K91tRM
IeW7SED5g3YHlSJoekkY+YwDU4/kQ2uGGl/qUH0XD1fDtDkxc9ql6rxh2Cwb04FzXgN32jt3ULtF
hk32uPAb67jo0hFmCrHRrcysfXi7P2CIMYhyNrHUZ7obJV0C0agrDJ5354w9iIPDoYUkkUjB72ql
0M3v6XZBF98uGc26E5hxtSxp/dmzPoxfhJzPsxyv9P7TNs0+2QIy6ZJAeLskdzg0R8fTcSJLHE55
nwlr+NltEeUbJJVjqyjvusHHxeZojl8sxoZefYYcK5qejrHtQluuWwC0bv933fcs6MZ0O8JQCUMb
WbGmGwcB+EkxD3z6BxvAnM9IqS5Hfc++tXHZiFBd4YIVyfh4Ltd9Ven4qATmxYCN+/kVt/UMcG+i
Rb5HdkozvykIDKIby97XG4DcZoXSAMdRKY9EqmRTL8ArImj5L3olaI57OLSLp6tN2yD2qO0ck8HX
P4qZaoARN1DW+CvNCoaz38pR7iPLv5cynZvfwvYvcw/YBbQpMP4b9qAPd2T7gS+5ogwrGVH9wTIa
J3+hUI28GYRc2V41cn2TEZUjVlY31AGxPuYTR1+ogo7+/G4MLN1xNfWDE5qg2AIwLZLqNuHdmZy2
xR0RMzOpIR5pccE2FHe6tItD2uwDcDR/zeVRj4S2RwpinUyB0TS1Ve4MVWnKCQYBr6E4qnDrZa07
zjKBGwWVidkii6dHgOMrhB0oyL1ZtUzFYhrTeRqPGCLkrygbsOkxhIAFtyEA0l8yyWXw5oB7Y1gV
zFu62zIcgS2mwo9esjMf1B0B0DFCKMBqAjDZWfgBFlVmsiTDkcqFQJj8T4Oz4dukPXRAvG/Uj6rB
XqLGo1DKO+l2t0ifEr5v3pDo/hXX6WfeHRnmQNt/aHBZJ38cZgU6OcDZToApvcwf2e+9gD5Zx/IJ
lBNNzQIIJahAp8itSiWZTrkzlU/fKI23kVHhndkVFsY008nxvBu/JYtjVFHh922/MtQ6Qb7Z2dlz
LVbGlqlLMZA5raI1uMmFX2dP3Y8UxFDRBgJ4mIvxom8TGQfJKWJJNOvWPmIuM8ShC34c/jlUIbCy
EQkKyISFFxJn0slHengPmFbwMhxjx4RLh9yVmwCShI9rE5k+RTa5bpiOowFF7npkYA8rUtlwmddy
iycfVjZHJX0IvvTpzD59DS4JYzh4g5wvPPRzSRZZtx2uRl/lFZQOYGfA9A+x8JrKZIwoY6bkk0DL
sseP+GnTinY1aIuaJj/krbxdkQTrze+4P1O+052gp9/Ty3X+fa66Kdv5Z2Q8B3d8AiwJjnS9MSq5
ipBWzYFKPpOb4rszSyODMysdEbCenXc2Lelu5jUGv9nHcRnC2v+p+fsmd+82QPydMgMnk7UBb9TG
Q1/lRAdiP+MQ8O+nVaQmcd651xZmBTbRbQm+L+JfSUuXIR+fGBiux9HcuzBuPdG7AW8gT9tzcqvA
G8UhOTDgefVR0D1Qm+3+pilzhaPQA1Hx3yw2fd/pSYP1I9mGvKI28V7Hkeu7aCWBkTGaFIX+4HvA
n0ljd1S+TmwvqnsfbGBhnWYkV8n4x6x58lANHWhcdwT5NohJF6YLYMtnVAaQrNU9A0GY+7r6S1gE
YFGRSexw+RBLbttXTLEe6MFYu/zHzsS+0P2Cr/VrxBzBz4qw3vBJzSMLVvR4oq4l9eLT/xz9CyAL
Q4HZXRsZq19Mf1lwEbDVmpcbb5ANLqiCe/AX8vLVshRAiK77hasAIfyLqkpcLaPv8ohUNQtfqqqu
dUHr0gpUmagDBnTf5HTHRUQtMz2ep+FV8GiQWz4sX9qw1plOMpWRSe1kKM+1WAkoF9GqTbZach11
qfxRN6vHGaTHXuwrDBNFmcjdjvxHu6AgAIznO4/orn8+2RbWG5gAFLqobT/Lo4c17KqKuVmggMAV
xZWucWAvgDuQwLRWQpGbHWdTEHbzINW6ISWncPjScho6qQ1YgyWIN5MisCDlYn0Ka0QyW8K65Y8u
Xn8Vkwj8u8+4yyRupZJWdQ04+qYhbMbCKZ20K9wlEZn/We4PXX2DoS7j3i6vk/7DDR8o4Wbo3AbL
yMrXJpWfXefpMFgb7ienmbellR2VfakMOVC/Iv+fJ8i80Mg7kTd3uVHN0ZddKStQ4TL0U0hS4yiO
oYHll8eccjQWFNoyHMVtilR2NP55rtClFA0C/ELcdNFOR/zJOwxjSq4Par9bpKPYLITr2bixZvw5
ef/dBFIo2E/UOe0spc2KlbuixFyhRJe0Tw6ChAltQ5ZKLGaq+JALr8in/q4xFUh0hAaceDzWTEiC
Z9vv2rCYhAMg0JABFsr8tMOa8OidyX3vqRHTQaezFGDIjdLt9dItAkbK7pRXsPbSULvhRttAuxCi
VlVNbFbKyef8LSfrwSPVfekd/i0XCP3+whPCZvbO/VaslMrJYqP0mVWTHxTOWt4wvv9FU8G6LXHy
xTEU7HFW+LhpJ2JIJ9AgAF8RojKAWjbGvCqF648q2+4U+HjMC4MHpkVqXJkpo2U6Kt1iScbiQpIC
WOVWpYLqm7eAcEzWPEiKk5YeBQ/Avuyb9o/9KlWI9Ex790YB/HFwaUNQLqIq5QNyU1+P2ThgfXvC
3EgsMbFhmSblw20BariF3LzwWh8N7kR0g2gw9V8YmggDjtvB6GM8Nwe/M1SuN58Y/h7uoLIbJ2LJ
5U/nOwCdwEF/aDFWCYvn/jI4p+BCCDQwp7Xzix17w6yDxDzxWWX2NjGlLM2S6dyqPWMkD1l01/MF
UuKcmByynW3V3JJY7k41Cx5gPGo9Xc2pCLAnrD+0A8kwR2CVPM6UpSmSz8t0gPJobhGvnW7aQ2I/
EFbI9Ht2TIMQb9C4QDtWo9lZHENW4NLUSKwVHFUVJtm67Z/AcuCphUhFHbPYkKO0tgOP36amqkKd
zqoOthz/0LTRnKCtGOn3j/G2OP1mMhRjED6/CBf9mEyNIpzCnQfjnQextWftGitASldNtJCReCj/
Pp7E3/um3egkIACaMOgEgh8AVzwWkSpxeEsGbfbc3Q4GDbX7MnN723aqXYJmiaV/6sy4la4m37Eh
QYmx+s8UGARbgjnUKKcV86nl+4lhhcLytqPG9NlkmL6280fufqulYrd9AQVe5/oOufNe1DutnJFS
mhT14YsFmgCJDuDbEX0SgotTHAaUMGVoqd+HMRBYIFVfwpghcBTBoHr+uIHTjiasF0B5WS821YZ3
oY69l6GE8H1rqzAThPgrP7zQ0yDxMAIAOvX3aBpxWX42HLLuQGhVJ5yOa1b/QNhzeaFwVMRFu/vZ
a75JTqfD3WJVukqupflAhaF4uGq7n1RzQe+7/zNr2Y934zD8tpz+sOALKQR5tZcR8z/Nu/7UZ4ng
xBTMU8DiQ+oSgUXKxUpkbp4oKOzCaCWRlSbaSyE6hoUJ8Gnh9ziqsUNrjZd5CIXUTdeccugNbA0Y
STYo0exTO/bDHEeFiiXwv59CgKYBo1EsBRkTZ17Bu5OHrvFGQ3uk2Y/94XqHX9Gv33Oc6F4h7qvU
sRD4fSc4uLWk/VylGtd00fcfY7ewqNqYx8cEUWkmE2fOHXLGrlPa5plv1dKacNJXwrP/4k1074Ju
KQts6HCCIQYm+rf757iZ94tZseLTtgI9e69hX1spi+csbGwwo7yqAQAsg3Sq1e+1iPKgYZ6FFLw4
Wg9K71vJY1ltyehvu6L9qjVt2kXlDA5aarprobiOBKlapEH0mGfmgqOYFIw/oaDvE+oOUGksTUTX
xhwaSxl1Yzgup2w289IfIOxhpBrlgMNh4Af5j3ckaylpRXK3RiHh6fos6IEf9KUsHDLZGmEocLrX
J6h4+QEkc0iwwlXTNsSO9wBVfBA2YcKj6j91t0R3n8zv9LvOzOgaC3YUP1jngRgjwHiT45GXAdNx
9INJ+G+ch7SYkgRRE64jaRFh/QcNOP4sAI7m+zNkklCHuRXfE7ZkPvA1OxpTv5SBMOk0sANBZDJu
qoBKFry82jli4KV087aCf2udIzGNKtBEBpInipQhYJJECokKxy6hpf9g8CsUfxVAYg+UhiL4XRTo
9uSW22+igXG29V3g/8/XAg86b9aCPdR3bsa76Fp7vp+sfipKlfxSm9yEXl4SrOF5DurumaluwQds
Vq8pMSV4zGXHZTv3c3qMa80nmPzKjNwcGk94mbCEYmjFIRj4urPZMX71LthdgeJIL2AHwOcUUpHB
4peL8lfPTQAlt/jFlNMq9kmraqB/q0pSX+iofjPM27TlP1Vss9IWHYzIlme8bbFQ6R8SpqS/RWUX
ZxzMiEZHcuDLalQgiH8Jw7jLvyJrN6GZVs6m/GYSWhxlgqc9dNyf1JNawvtxxdoPQ3oaJLfu640R
HenaqeJ7WvNSPIKqh4/OJZP6tNECnyX1hP5Ffgjz5oMqZ6Gyyqe3c6V+PnPbNtgArwYa3/8C9te6
F4e8/ZIIM/8tM5GK8xP5jBUupQEWoQZcwize5rTza46GPYTyEl2IAj4nLAHFfjSSdrrjF1JaLq1q
ZNXp3ldLbrWF/q/D+T/AcZFzDsfi/gHTDbLwGT4f5GLqTWc8jwHo9F/LN2VbjqIlEklcsni75GEb
1WvyXfUxdJYcOtdT9EGZtjYW+MiKEEcbc/3NgEdWepkYrTgXMlS+yEUDnC2ET820SRcQKrwckZjE
HsmxqoibMqXfB6CdzfOTTl6P4/g2Lrf3CUtWZSHRvnZ67Y/wGD+yqFjAzW2UBaeguR9xrepr4njs
VyeOcldDL6/9vmG3hr/UIAnCIHl5Yi7DMXj9qbu1sKmoH6TqNLyC4qZuO0pEeci3j8C4XySjVg5w
/WrRwG6opddfGEcGWJJ6oEbk1kmwAGIsLGc+jl5GU+NOUcjERM0W/SZO66+s79+7sZ8PeC7XUlN5
sRJR8PG0HhSzbLJ2PoYi/29rtXekFtcX1xcSQIbUjMVJHkV0s22EwbibfMq0rTZDrz3JZRIw0cKY
9BajDb7oI4gOeR6ALgLQlp4Y5+dcHUIYs7wK2gZA1Q9DBoqhjmX5zHosNnvKbrIPj+mKaSL/zwD0
rbWvlnt2j9kouZfTDVfeHgaqbSQnxrwSkToZY2oFtO3RgOvHBXRfsScsik/FlW1YO04DhV31kkAK
L7EqNB6R/pr3o67PgZjPucOzcNOdynyd4QC3CV/gropGWTX3htNWCpoN72cUntfwqVJjqWx3sin9
TaG9TcZCruCJrzk3qcbVGrn212QiO+urIVVTOGvyrTOB8XSq1dvkzGuX9zzLVL9j7+F01ThfH94p
DnYjr51prEXBUCO2b2ZfpQHFHiO9ZNYq8vc8rEQvQGG/9JKWEWCc1NESJMrvpfN0hLTt62lvhSlN
/bmVRkO/thkv77zxQZC1WYZ3LvWa/3Fn07DbhwZhvezx0REbDAcuuwi6b2bhlFZWFtTx5nIm4Xcm
vOx4Ah+d1qPq9iloMW2ktmQ6JukxMTQq8pLsVl97z0r3YEieqCsOwqutjul+rgYcBj5xUSA205w7
Uxu/mLUGdghhdErjB08IZPIMVsBaJM0u6GBS4NJTx9iejrnLlITk5J6GIerppXqzhuQLXhMvr2CT
DCitiCd3TzK8k3zGzEr1JYf+nfHTZDzglDDRMHA414DxSNvj67EJwGhSE7REDYK7y8ANk9veLTGn
QY4rz1RbzgEl7lRhdAcUEiByZLDUBAltUmoNNLuB71n3qmi0q6pg9bcnBkXIs6DNLKNHofyBkRc3
3bCSAkfCLy++N2yQI8PxJHjIkvC5J8Inx6daQ0JxpUfDc87eNYpLeCh+3wpGgKnQhYxv0AvVPlWn
XDA8eQKNcieOuksTxZfuXjQkqUS4khu4m0xxpgZ2XPvCbakYEnE7L+VeVQcjgnpuITa2BZ1bLvj/
bXF7C8rF2xyU7HLvvhmC5pABhQ9qzdomcwe36erpipjLIPcLeTNZgGrzahZN8+AyrAAqisB9S248
zY/sZ5UkDDS4PjZBN5FKn7OzE0/yTTC1s5k4QvDaVM6j7c3hy3VqTxTrI7JCPl6cdedko7Ha4P5E
Clob7n6H7vVb7Y/UzFN+5tyefy5O8sWwzDblGkHCL6O0BesDoslRYlWohaNjM9b4IPwKWNrXfDj2
0dlY81nITwz+r+GzaozlJ8VC/oewHm3a/5xVip78qAUTqiEGUIv5iKa3VT73oy1t4DrYBjKQ2igP
36ZqaDRILAmtdf5GtmYwCZcJ+7MhcrRwII87r+ONDg42uhhC/B0+cheQl4iGIH5sfD9n/kHTCOGu
JpwIaKEnqltfKkfijcBd8UfNKLabQcEjaoB7ueGnoDXHUW63JvwZ1UPw8PyffGoPmuYdCrG1wwsj
EGmrCOzYiC/N6hkN7HaRxIft7Hy2KPwZzRO0qQWc1spMkbcMJF7jHvH+0qIVlmG+7h3WwqOf9NlO
fY5TwDgQq5a01xUrd3f2rp2CUzBqz+IGUqvr+kBB/scjRRslb7X2ozJ/FvRoZ9EP5eiO6joUg3yq
lfLK2ybibhv1F1aFOTIrnuDw9cJP/hwXOesIUkD+zuBqOcTjZ7jU6obZvIWmJHgGxoA6pJrm/5ZK
gWWaSTXb/Zk6lH4ZGGFAc22oICqQKok404p2ZXUGlBIT7eOLdldfa434IK7WPixB1s9tk9BFiFNU
5AR9hYMG/UlqplGq7ull6rw+HebqaM8QVFou31wrwGj4ri4xam+nBgi2gAXyNhcIkl93HTKUiTMv
DsBf1CjbY0KIcsagmRlOCN+blt1NWLKQzmGZp/bRmrsyLrqP2w5dMF6CEYEE9VC3qP8g8I+KBMlI
886SLm7GjPHRKqMRn0KA29kVMepLQ8fFT+vKz5FOS2/DuTHWy6X85zAKspTx/DkApxpb+PftU8hR
X0ojXozD0jCwbVWTYsk65Uda0ioXf/kxEuhfp8zxzhQEQ+gK+QTnDkp3Jh04cFGWbDVpkrCxnYow
siDpeAEHA8lWrNfI6jQ2pjgIGPoA8tYW4mbRXIXFtQiXPWrN2x3Q+sm1G6Kb5WmbZ3ehin+EuKlE
EXEBxVHNCUgWQQ239gu7Yo56bkuDxJ/iZb6rJoahTilpCOkBV8fSb/mDLN5hRlvaaqGRkYQOZMMP
qFmsoq1C27vN2nSIDT65TxGhSKdWYjnKoz31FjRGkXhlkZQ/qSy+cjOxbFbeCf6PDFmM+iccCOGZ
n7aB2izDLjrl/g0idogHJxggdbnMkRKEHKRDwNiq6JTnqLQvBbIV95/1irLawEJ2KkEMvHfzXulm
2HR3mEgWuH9R51tdCnsLoX+bUr3d1LeFbXsLmDU/vYqL0LEgbFV91+GThtJbFogzn9tiohvTW43K
4bi7Ez+bou81DQnDp0ayLePkDMOR51aaIJbiT03sBUsIM0WNIIgSUCMmCNvoX3tmNtTCEcGIcdAz
NdrlGggVhrjZwp9zsZ+SQHelDtEh5k2lwguzbR2s3Y0QznhUN0g0VBtVJCBmzyhf2g9GKV20DdOJ
hyV+F0kzgprF8v1wcBkPhpIrnce7yo0RqzGDZMmu3s/DFHnTsdiXFJh31+CZfN0RCu3ccwnqTpSS
LMGj7ztybpb9r23+U7Ew+9n2MKNPx/f+mb3p0OK/axfwmmcUQDeJLgL83L1+NDCf98ON1PuX43Fo
Wg5ol2ZT13rAcKjHGBrdrRhMXI/sBY5OnYNevPjfBk/O+MsSiFvUXh75Zp9K77NGcVCQnYgwGgOp
gzfI/ih6w7g3lDPJDInftya00a44UjkFh36Y93klFX9/cFPXUJ1kO4brqzy1/PThXXCBZmX5S5p0
WRrtUXdVwLuRkJs+DK/XWvdPBvj3cGcfl9pukJXF0BAXB5/1zbMLNripIJ+XSAsP7WwkCSGqPns9
SnsOTMTDsc/M3J6JfmIex+rwRYmu3ne7NuFypr0mz2j7bg3CJCgug4rnHE+842H+P9f0u8OcyDCu
DE9aMH8hCJsYf/8J+Pbg8uLeKIfjrvbBORsulXk2cn1r5Gck/7OwYG6diGrWxGXvDyQcluW9lKgr
rNLKu9ulaB2bBSl0exDYAvyCjawKU1OG5GHpk3cz0pOfRB4k9aEwD/2J8X+Q5OULU/JVRqZ5Um62
SBnwM2hfqkyRxwqjYi74F9To+r1PR3ErQyX/Rtdql1+cDhx/TrFxmKvr2nwRH8/gYFHPLy54o08C
ACVoehup8ySI7VJCWLKQjG/eVNqEiaJYsxxpwbdz90s0JSJfLtm9QMlQcQcYc9cbTaeb6iUfjIps
/Hq/KLvTOwPFWsKiXDouckl1ON3s/d9oYWa7W9gVyPZ7Mmsy2055VP/jODUngOH1XnCL0ORUquHk
HTTe7TM0ukFuES+nrl/epk+1BVBAGqldJ1Na/JOhBy/EKWOA7dSHQhSXepJGRPqGvx316PDdFM3z
9usjIVnUErPFAc2kO0WXCayxZfbQAIrDKXnyh/j9IxNXH/Hgx+OFgxdtw84lz9yCvTpxM9HB60Lg
hwMraJnz9WdJiIuxepV6oP5cFVEoSjNdyUr3XZzLYnR5V4PjkgGp23naHc/JofZCH5qvIK3tnItL
YogUEiJzggQfoQgJ+t3EYdpNTT6YIDvPQeIeyKHaYesJby0j3myZlSQmNdfXzEN+TL6yyLngSmh2
iBkmx84rAP44oiXjB24iS1gIcMb90qzoGdudtSMloSjuWMUgVsL5PbaLUSC8GqInRSqq3zCNdLh9
hdPhGT5qs/Yu/7IJJf/HK6U2DNSqmMn44Thx+YY0XkBUJpiP87IsjoNebna/dYRyh5LrpVfwEViM
MZt83f6rSMv0nnYnDGE3z3HJiIInsol8TrfGc3Lgg0CWOjsTHTG1WVmYiUuZLFQyYbAKs9qdzUR8
UvoO1gAAp8GI3Vt1NO2dbtlZbiTqQo08qlImq6Kw+oYRqWWGaPHvtpcCCR7UUvgouxj+JK41i98h
SXXRw7C62OPGwfP/eGVo06asx8BG0q6wWCJJYgRJc46Djw7LwWrX8LoG5WEkGxpv34wd23qr4iPY
ckxpbUYl2RnMx/J4Eeu7NkYkx/LRvjY609yIc+k0pJeUJQE0DICLttOzaI5Lxf5xOL7M1vyUGxCq
dV6VbBKn/ABBeoBCfFcy8Dyq0YYaHLZSMsu1GdTbBcpKPP/4ypSDVCvO2CN4D5CZLxZj27YIX933
zogiwd4lyoKi/DONlIKdokB9nawilHa9bbf+buYhRWidCL27zMe5W9AEJY6DoK5LvTs1MhxZ8ETx
RsQH7QoTpshKH73fVc2vA4Xr7Z96cUHXDimj5ovtvWY3NyHm0Va8v41Lp1sqolUP32IK1VBfb9ig
uzH8FXsEYRbP1AhWN795ECi1aQiC7cwgmx8H5Sox71jkgadP+wUxZztRbeTRQXcB9JIR8qFBKNjm
HsScANZxwUK5iTisKX1UQ3+fBrqRuGEtxWcg9BYO3Bido7o0PD8l/xbUnA4ht0Qfvn36qBVTtJiF
VJ8o15M39A30Gt17fug88OKXqgiNYGFG7qnoSygTb4uIZLuX+Inp+uoCJWn1St/C2isBlyjN/e8T
5dz2c2SOYAz/jR7q81Mooe+LVL6aO7ajJ0UcEz5N5lOhdVmHB1aV3tIevDlvKyq8pSTzutG8dak1
f4HRxcSOWyNynHfKM36TTsC5ijG5Fwq06NGWTHYbiqnqiMfTvVwzynZwINqQY3xsZHE46ww0Psh/
P7hbjEYIIT4cYZEIw45A73Et0Tu0eBKaCvjHBOaKV7V5wFB1be8/vSrlMvfX2wVHEHao3+65Rj+n
BzWCy5AVVK/VHoKfn2Uew0JqAb+qe34ByEJHBhBJniNN9Z0cI7JY1BUNtrrzkigszAbZTVId011l
kFnvsn8M0nz+3sTpOn7D8UColwdhPgW7tpqNdLEoddIKZmirQ7cVRkjPi7NLknvJm4vQURLFnGQt
8XQ8mprDCkRhGeMEF8Nk4nrBP2FlVFhGiOGk9Zvt8iZ5pOxaoiPlQ1D6UJTrQ6XU1tUxj5Uy5G2n
kfJBLM5BMHapLBHs9genUJdckF0AvD6mMTCV2X+4rk2K+WSNmjkTjvExqjyGZTVYB6A3a4oAkwaW
XZMrZG7e9MsCVnjTZU0qXyMNT3NTOu9FBuvb8xRd/asIa0IEREfRJCoVU78DpsFJpaWzLBSUzmSv
JXAVm+YRyb6rwDG13C9KKRac/s1DipAihXdrCcTh3176utf2xScIlLNz6W0aQehp7wImev5o81PF
i4lEa1RBY6HsghOTd7YfTPGEFHFmA5BqwYRqVgZGzL2jbvcm9DcItDsa0dCh7toyHrFGVMTRLmJi
qjgr543m0u0MUfzpPublaMgGAhJVvnjUdDYp+dTLHFlVop2PBHzY1c2E2QGuxGQ6jrhtXxYiyoxE
5dSB/OxVP++yZNlRxbwT4kpf/gw4u+8YqWcvkk+7Lo5buU8+mRNphPeK4vRtjA/nZeenlBBJoyCs
h3nxZ8x9AFyMsulI2SbKzpXn1ctDiVbO96qxakObYTssX8gAYl+viAbzF1Z5Y8Ut/ekVWOeBxHJk
1wYC1hKq9DE5PgGnyDJpXqUgrYtPUaS6CT21nrJDj4RGY95fT4P1popyYhuF+v327ddr4maRvAQj
FDR5dR543Q46ioikTBjx8Nt2oFp92mj9+RzZ+HrzqozEq+lgqHKxGpLNZF1SzjLhb/6ncxo+lHAk
pCTI7Kn9sDJauxsCQDnPJoyTT8X1XPF5sh1ABBk1hMmyZibMFV0KzXfEeez1JllN94KZUv17VaNr
BHlWB8czHXt/FvPQbnh/jshpeRhrIF1LZIkhfyA8ICXe9nvV3dd4FkUZAljO0Up2ygMI0xC8pSMb
SbVNlnWx+xExgwCowgrJ3A70nJ0fM4Wwerk+0e+YgMxo+8k5BgRwYoYsUcvJAclufBQhxKrgGWB3
gsAD7kPGNxs5mWL6xA0mGmbiDSTXjKxdawXzFoCXgFFtgC8zFz7HP5jnFLMQlCCQwC0nJBkT6ihN
XOGe+rAGwz2Yijp+KIHfHYGQ2nirEPRzsVBHUDwJ8x/gieqnex6JNk6Q2V+ZenmFzdfVF5r2QtBy
ABlpnelKvcdc/2UmF6UMdmL62B5vikH33ggQveG/cLfdudh8nsCBtwIvcgoLIkz5AHOX1mqTMs1B
ar+u4bfLEJ+1XOh92GIuffQD6i9i+b7o24P9ETpuzZttIAPAdgJZNcyMQMdYdeXXxGbZfXSLm5u0
SiP7HMCZGB76/DJM6u1uaAR6pa2LzXBcMdpWJZkf4zgSgz/GU7rfJexBCJPetyTgccO7jkl9Hscr
t3JG2OFWmM1/CGwGeQhlQHzBg5WHf1eCAi/iKaJe05qIA9fg2CRVU1h3xhXmYQPEJDlS2CIBb39i
UpXcdBPJqRsvwi1o7lntxHu0d/a7jNPkNHbbtXIjybuC+iE+75Z1XWTEdaobKYZQGeDiV/eJBIf4
IO1uNIM3DtqyvRaSDYo4nbQbOKJ/E+5oc/rFaMXG1JNpkvK+tAbDwVs1ZZrwg7+K79i5skGk/Xce
W9iZwXGl7xf72AIISLyLuAnhfyT0sdGNBQjQUxXCJykoL5XlCNE85nOYvUJqVjfX51C+VQs1iTlp
h1YBw5b07ZBZqv83ybnA06hEpLCB2E7D+z2EQL4W6ZZrPZ8tZ98fQSMDX0akPHWpyc5+HJIBJUht
m2HRygecIltJKtwLP6jrwrpCpQRskAxuC+YYFPJIZu3jkK6CvT3rPPUTdOSmU1a553/9g43NG+Sw
3amQjnBqSYWG18OvfOKsx1GYQQ5h6SlddeGPC9ybrAgC+WO0ayH0VyZELWKOwfZCnZ8wVVay/aJr
iiRTOQe6/huNPu1l0yTTOuIwn0L3QQdL/SPxVYQTxqOkVNdBuEDDE7qWK+vw97aJkYEb8N/aIfpm
pfMld9uGnxswHrSJBCZi/guafgzYhW2nRg7dUj0kOVduOTeVIzt6tdVnLqF15prIk+1uJKSuQ+ZQ
pDAilFZyA/8pfsEU9X2q/T3ldbR8SKDEnXVIi8RHo1CWL8U4y6uRiZViauMDD3im5uauJQbozseA
EciuyOyIppcbCe8hlD/KgP3aqWs3j/e3aVsrx6sjSde7NGI+/cGCVPzzzhqA1I5eQgZHYnXGwsRt
y4VS0CqWCkEsIs9C/c/rTnDcXDEFmEtAyv5ndpUglRZnwSYwBzF0NAjw+2UsV/2OnttsJ5gBu7Ye
JSYyy7N2urAgIfNncWo4z4obKRjaAwEG18+kxIZNEax5ZwoEG5W3tuWNfubORkgvmMBW4yscoZj7
tXIca2q66QJvRJDxNp2yvO9RsbOwzg8USRb0TyG3c9R+tHqNl6UUmQV76p82rCRSxmjhIDPqbKsp
M/CjgadrXPNp3E7PEIPsxi+WCS/LMqZrgF3Gure4M9TFW1i3mhs1GJ9wb7yUPrbxjrWI1O+d6r6e
JQmLQxkvfK+G14bhH3UOQdOAcFKlOByIQnIhgfJnRsevipovNQxMcUBsm08uvq3tKTtipSzmqPEc
zTk1QXtFKeIkUsZaHcTtKGZswmJY9mIdp8j3L+D8DTIz8mrMGWoZpKCwJaS1KiMf1DMnV8Nnwf8N
LpiTfdczSP+QuHT3cZ/5IRG1VB+Y/ZKBWbOfBIGjCGSR04U/79Fpe/5t4fVev8kmniJMcnBzVcRd
282ym8jrO++OPulAC0pNkql/XQN42rxKKcC5zQGcxY3ChClwcMTo9d04ldEbh5W57QdhRflQCXlk
xEv04NJziGoJb6yQZwG3aSRDCRy5BDngwDYqhIAH76qE9QTh08wBKmyDM0OZE0CDdlW9njS28t2D
wqlKkH1jZIdmM1OYePIShNdoBfkSIA0PswlaKpXo7mChy6sO2Fpd/FAG2z31+0rCMbaEuq1v2Ylw
f+mwaWibMKff1vT/KCPLtoVseEaFlEbbTSKnXj1RLj2ey9nYEBWdOeDlrPcRPj3OcWSWEA1LvDVd
DfJmPzo4pt9wAHek8Zcx2i50BQ59WCKYXCyuO/oTTytg8X35AwNACnLUvEdJe5ibeN1Nw3YN9Vss
F9IOYTkR+zeax3CPmw2NrihKjUlmhfn5M9EbfnJO5PS7gQS1s7gElQNT4VxM+AfTZA9DBGE0oATl
O6FNJQ96IFylUHT+qT9ibM5sp5agLew0BLXTfp8TLHw72cmxI5KLBFsBkD/NPAi0u/ff0VXUxPBH
I/0nirfFLkDOWkRXuJs1bPbcYKRpsHJxDEW7SDKC5MbUCmfd89vk1o6+0xVq74o0d6bAuR58PhAz
yuBhmr81hnHZpM8uSQzKJjL7+kCdFIYTfAM67nA8NHqxX6PbzqxLCUd1h7OV38nADztDdYJAwNHs
kIsDRt+NkBYjE7QY2i7w7E6miAO6LkqNpHrKLJpeMFpqZczUsazW0ZSWs1czeL/lyLatmnaPDBes
ehqCUbpiPiHQg+bTrDGWaYQs7+X45KXbyx810ot8COnXpRG8B83X6qmcKXG5EHx0K/7b5ncpmja0
FcACrut12N1AZP/9SqjNZ6pfkvxEiUx9DO24AszV6Mb4wD7rrAOmc0kttM1f0tqb9crKPct/ELxp
sb6A8Gvykkv/TUk9oJHYb7bO85vDz4Q06NxDSoDGPnmezTz0N0tpLhikAQh0zUt8x7jCXtqBnddI
EykNR/tLKjlE0jziEaSUsr73pCHtExaq5aHzNcXbxcK7UZUJ0U5lvBUzGh1WucgKKREobHUT3eia
GfbmEXdTSC4vGXjy6yWez+xZOAAj5wo+Y+YAqTnbzN07asQW5axHvOZGFu9xvBPXoS/OR1nIWLas
KVTeL0DfzvjQ6JvM/3a5heWUK31wy52+qCWI/sEaAKipHMHS+g338OT1R0tSH8++daCfsQ8WhiNb
6p3ka+MTAZfrg3uJxdjY2Orm2S/tfKT48ynWmaarJ2iBMlVST+iuIjasC2dGMbKpnQyCqF3ci/FB
bkza9vYhKU+Iy/aijMaSx/AOPDbdVY+C7ciBt56vP3Usp1loTR25yLDYGEwRjho9SyrUvhFgDQEd
MOFsFvdNB9yHRVpaYnurd/rGzGXC9/3g6eS3xn3APK18/t4peQBMphV3yA0TLTDcBtYTJcOVLAGj
YkSru33bmUkc/HctDOav+y2XIOGSvg+2f6uwuhwSnFUeiLQ0ruyQS11dJvoO+2auIuI+fhkihOZO
gP0yQG1FI66VPNLM0L/ijGppKIDFLN/Y6gmn0ZHzGajlQuWY+NeknPRwMBvUdp1oEDDYWbaWdNBP
SX+B0TJR4QjvG4ZMgznL6Sj1aZd0Z6kBXU4lHalx5cUjILX6fdHmpZQtGc3atpHlZiQpagAazdiD
gYK7Hpor/Bf2UZaucj11zlemPmuiPPDWSgcZNuimRZKYbnf6SuLW248qHMnNZY3KnZt23u6eQetR
5LkYaazpRRsG657Z4fU839Q9ZRFndR7hoQGYYnJNrUzzHyLxMXZfN2vo9ou+22WAj/JL/Oe+4VFi
YrOtOBdwPoBvQzRdpFns2LkPPrQgCnTsLzd4SS7ldNRUBeIGmc74vXvwhuuIxO+7dqP1A9nd3ZwV
KJGK9vlZZzcRSLWXtWabTP5290mn0ELzDWOzwrbpY8UH10glaATzYMm3ucq85plF8WiqF5XNul1H
bwFE4Iw8gyN/isb2jGBnMfcZUwBQmbfsOTyphWkUWfGaqn6sccz6ebMQN7RiookILprkrQrK72eo
J39IvQ0xj825dB0G37rpAHHHc8/D5QcTY5hloyEIhzK6ljhFUavf9RaZOZ3XeouFphweSu8MNNqr
wrNtaSJPYu/j6yqfpMHL4NbiKARFjbOFU7Tp9PqgBA3G1JnhWzb8tOoe3hLPLgep6cvDUcqimYVU
mAz0tcZ29sB+9h5tiRUP69Jb8ifpkdii8xwA0EqXiwLBAUBov1oUx6getpAzUyc8gYnJdYPsKyTE
OjZErYOvFbFDYTS2MKekSN619frRe375ir8fbM9QupPc1yHscgQl9zGh0wr9DQk7bEGrWL/pz2w5
vKaJRIYIMZhKcjygza2TUj9oe2Vma1wNGTfCGgSdOYxZEfWgEn/B9bezUONtDbCaPMhObNZ/cwy8
5EF4iAMFGbWbDe7cme4Yxys9i/heYMBaOMiV4ka8KCe4p1nKBmcqrkoeOJH4FmJeP1sRH0YpDDXG
R7VORVDCYkklwnSbPoKhhlv4y4nqcsRFKKAgcFa12mJ9Wthfz4HQyXrG5bM8GwpVUg08BdGOP1ui
vNRqBMP2VPK9H7dmWBFM+R+d1kY/A4epOz0V+6C473avJeAnAjn+kGXJZmI24o0eQ4833LfvxU+W
7mn/P5xwhO2tRTRu0hVNIarYKlqVGdCztiQ1ZmmVLxHtojgGI0UL5SOhlayabpYWbedcLjobe+wq
2NRPwbeumvzUey8g7xlEAyo53Nixo0u6dSQBwWnUoilaay/irWsO6TZ/raXylW6XGVX41N2HVE0L
y6GiUqw7YQyRlp3xxUQY6Vnr7LGOYQgcOqiTDfeAr36hbefg0ctmg1GFfRiE5BRSq/d9VpAhVGBx
+FvQPMyOoXIyh4luVXr3wVAmEPQGApg+igfmJeW0bjUEZgSxUa41Wti8MkqoKmhVQkZOLbkYCVYI
FFyEsHBdl9A1h/xFewNkS4cdRP2v4GPGig65uc8MHasCToYNf2sER+ptqqDQNcQwwQjH++of5o5w
xgAgVGc3bRNByAj0RalYyxVFteNgL0XK63oM8RdYfUBig97Q2niOf1jU0VLO3x/TGqEhrbjVwzfT
H4DkRJMkFKGlg6ZmyRdnJ4Pk56cv3gGxFlJCxHTMH5YnXK8ra/8MBxP4UYVvDcyVBD/uv8mGt08J
IsrTxQRp2B6nGbK/r+elUQ0l7ibM5BgujtV+fekX/IgiNXsnX0lsVOfMqUDlkTbHxIEfV1vxKquq
i17JWP031fHfY/os/rKnXeZH3XDjk+Oos2o+caay0bLmLJXW2xTmm86Fh+SN5V1zz0hyB61Wsei8
Nj4JENo1o7tFbJT8OtOJIqT+rgj0xkte4xiCTEZaRPHAQOwXcjPuA74XsMBs7ABxmAJE99+lb+La
XR2nWhT6BDHJZwWsJYLCQ5y8nPsuLyYwkhYmGZuDb7nhkDfj9hjfLCtQSvshQwMDsZVdKHpQCFXz
4fppLH6quyxwypzG754g4zGzmEA+rXv+NPfs3WbOfZW+yWK8S5272DPAbUdDYpze8DhrNyMcTA3I
nxwc+1i8cbFNWqLafdL+K+OBOzhKr2r55zQJB97FclxrTmFAyWGruLSEg+1SBzFFJheFIouHYmeJ
PPSaflqPNsZVW2QpoxbdiOP+S4tV+LFi4ryoyHWa03NmzQbpmPsHcZeI8XV6ftq+WMuepXoT+6mM
kowbpNfjpfn+v8OATAvBCD8AsdpGEFVvyJ4J1LPaN9oH6LKxUfUoZXW6zOGOL5TfnZum0uk/GVjm
SnAAg93fZMkpwSDXqx7vbMeYRpyp6Z8VkOm/4vooDtV/ouv4Dyx6v5Cld5Tz9qtHXeHyD4NJbXnb
axpoArjE3fQoj1okJTsMgB9i3zDhCfbV75s6irWXAAqMfkAaaB9mykFGrHJr0fsDrPA72heva/x7
0P3qeiWmHV2AuTI8JXYonXoflIFot86cZy9LtXefuRPyhjkNWOK5qUDO4Vh0HNcQaBh9kms+k1U2
y7d5R8bXzia11K0MloTXisUvq1EStJ6XX5lRI4bs5FQh0dblibGFAXsnRysiNTy5iq9QapzJPURV
4wTxmXlO7SdOp63TBNwEjanji3VLMFu3t8n3QxR6sqOXsI7oNqFW1HLBYvaqWVo+jYUzdKBxs99Z
ooc/XOhEf1pSqLxNIdKL+LDtYWRJLelsErg+P87KnzEASf1cYopOJSMRXhdKx4VbwMEnZK8ZncQe
TiOrz9b8QDKA8GqOtw/Qw0uq0sKX55d4p2Ce+Y8t52Vf952lzbOPe97FptEWlOss7Q09xI55+xRg
F0Eua1YIpLpGZTFyaryK8rp5tJihBlUcZggnnxxlR37coezs2bpY+AqFWioxsdbCj/jXc68SscZq
XFETTKrspBvyOT+ZrRjv/Xo0GesvCX6e9oL9Ze6r0P/oJEHabpifGI4DTl2C4hFBEYi8WymMGw4O
otKrXpMTJhP/G1LpU6gwGTMwoIUIKyOG6J2+AmzwTxhEeZ7oFjGWU+GfjI7nR0mB4lGirhdXEXxB
WOyij7fg3DMF44IXvbdJMwEZ4R5Rpb9yQV0Zr2Z/FaYAQ0eUlBJBNFZvbqROcnJBgrSwPqWFr9fH
iw5J3Gn7eHgON7rOZ7jXnGApF1ozHD+cNQN2tgycatZB6ubrOdDtGWr3+QwGfxFxJ0YyWeNpd4ad
77gjnRergNyPdoRwD8MewiWn1XkJaeBXEKBK6gZUrE703Mt9NtbJsl/ChjfSlKKnV9AbS0EhiyVy
nOQSgJyneBvxyPUj2wpD5y/8CMm/xd6vxsOlEJnfwv4S1/0bP7FgnJbmDVAvKMuWOjgyqgz9ftyy
eDQqWUb+qkwtZYg81tW3x5eKCJGUsW5jqakGkpXhDOIi+EZjClNoZMq9Je1pXibcXmqgzvR1X6n4
keTv3JEBGJXRZuIloVszXRx1OEox8OJ+oIfVka+EWQq1RD+f3s29dm4ieQpmUtQ5wZfqYKYt0W2l
Uo/vYcPujY1lB2IXQcKPjpq0rxpzx8q1qGz4yZVRa0ZjIeIKmNllb+PJfrshyuMY7Ahy4toFCxsp
dWIGTQjSkNDTYPx3qjO/LZ80NMiEB90VnYGhrNVpy1DjxnWL/qg6hZw5zuPb7MLybAIuoivUhLT9
vsoADXRaACwXHRaDYOLVw8qhwhNmo7QCJMovmfIO7b44Dv044TBwKiaaq1yZsom+tU4b5rSXYXTW
AFEZouQsYbzJQpbCp43kpkWKUCJKujQbVRVRHFHDoAOOWj13fOGePrKesEMk/CNX+dTy7cyIKAKA
ODuXNWicqv7IOaqvzQa0fy3GabrrRL9k+S1U5EDmy/GGAykCSt7h4rq9Ii/TI/J/MVjIOpwl93Id
ezxA21kBCZOc90zwYw8k+v2hm7nUmIddC/0n750Zp8CHa12kWNn/Le/oKai8jvfcfkARmceUZTkk
89v5QhM6l+n9vlqiRGS8IUW9hb4bmMKpeOP8bUb4/+bCM63HtvDcfPz+hMffUIj/OqGtfVZ1Ndaq
APG8kFzbAWWi4AMrlLVVrewpWIe+X9+uNGJ8/96EYvVSiaqKD86ktym/aMuwoeLw/M8Hk+71ecVJ
NF4sWFrFzKPIYtbSwOdoCrn+1q3Bi6PUeNWldwAAdA1QE9X5jqRn+ulPiMV6G4HwAh+KNp8xOvsB
hUX/CatI/YJFkgD+uUZvw0OpCjx52w8j4tYvAiyTmBLljQchRsgXfIQTwVUD7XaHcX1+qZMLLeiJ
keQFgt3+nhi6zJq7D52tSpkR52J7aDNNw8pzVu95TQrJ6UeAOWUGh2quA0nqEGDJdjMwzcf/I02V
fJA568GDgZ3cUaQo4vFKQofPz93i+xWu7EPUBbAUmFHR7/Dxj1cYlKkJscXeq3xiT2wS9wzCDLYH
OFpjRJum+tEDCfgOOIz3XWq31svM1k88CD8hlOypx7nkeI+CK7dNDiCZEmSqp1FW2nezDCuG0Mc/
HuYHE4e6D5a7vxZoX0CAdsjyjijLVsn7R5Isg6VXTyq3ESWzSq0S35MKSAvs68Qbb5j7xAUm5tUg
zf3DZglCv11yRQYeAYMK5ddPkn6zNHfwKm+d4g55StHwzbP6oUakXp5UpSKqkO/dgeCi10py6le+
sVBFe2ujrGUEmpR54FwwB0IWQeYhUgirf7NBbdkkPEZFT7WIYWrZokY97n1Qx+kY6OU6PYD+wNFU
l7EdYbTVwDnRQTbl+v22lMV/0XuwkDzAwJJFgRCXz3WCBKWtA3Kg5l3ENLHYUGb00yuBS5+QDEER
0gR4E6QpiVZ+xpto65nkXEvA8O9ecINBgkENFjv5P7xyxD81BdDWFUbZFUfwqKRqNm9FQkYxTApR
uEdXIoe0AM6mDuUMgY4Yr50lHhGp3fF5rTqzTfk2gHg+S9NAYH7w9KBpQmUr3jC8TogY6gxnCfO0
Ykd7UHbgAvf4l9LXXy3An63XsGujrQRypV3vmhYJgOc8d5z5ol0cWOi6fhJjgak7bNjY3S4c9zyB
D++A8dPty8KpH7UhEXx6xBu1LursxqfY5rm6TeBTDA4uxixKrPHl67uD2HoKJz2sFQFX0KJROxi+
s0gC1QhnSGIEWBRa0Y2oqZLJFhI7ErWZ0JT0YKMw4Ik5P1yW7XL2jllPRWhoioqfLnsdph6fZlJl
B6g7BRfOMlXLIfgLuI+3CTlAYvpfDWwChHdwlHzjmG8UObz2Nwx+5/82vRrHFy6z4pcNDdp6YxlR
yizysjwYvMQr+llyKvgp0yRRydXJ0KeNFO5ADjGevHMLSfIfjbYwj70wdWGASH7F2irhdM5DbEAf
x3HEUIzSEj/JDfFGpR/1r08JxoOwgeXIHIPM3zLD+B3Bly4CLGXnnOFz1OfwGUUjFIrbNcBTu2jX
uMcADPgcaZ06XaOSq9VgXj2m/6//60/w+bey+gHfTnSQinzGQ5adrrkRYwnhYlfZai/s3hvxEqHS
XVp72QJUKAZRgvem6WKhqy41vhULIv9KPAzhMNuXYjwyIUwDqw7bNbCQYvBMvC7FJUsphuN+gsmx
dcw+tuvZ7Zi8lpEJy1G2OyhSd5eBckjox8e+LDvDxT3hYJHHWP1LwBdyldlNhRepIeeAyoq+DCpH
szzB6px44493/sTz9xh25xfu8Re/9hxYPApJMknEtAyG6ogF8ZS+Iwo0B94r9Wss26+xlY7Ylejo
Jaj8BGqXWm/8mKuKw6yghCHyjBz8tCnpSfMivBcTIBTxHbgLg0030nT7bup8yRh6UxRpnUTi/g7Q
lAy6OOBgZpckwRAm1aL4CP5xr8+1jccV/NbgK5BLlzOTf3r/8AioZpNmrRWM7Z9zy58/2nAccDgG
7U8jlSpLFj4wFDtU5MpfHmLpiE/9MOU8pRPP5rpxt0gJA1W9EMM/XWVWxsGBPXbxSHG/sARWxygb
M16eDIy6kfXjrzcCEKrNno7R85Q7D+Um6nCK1JmfAtwSM5z8H92QLk/y/PeNhwSMJ9DOZUHAzdXd
cYTg8EIk9ONdTmG7hc0LMXCEWW53t13tv/eBKAGTrTCHGtR9qO+Dw78c8COUsHphwehcMSdemlnN
neatp9lMq8tSiH64SHYAYBew3hAaaIrxAJ1MVzv5YhU9iGBDbZSILZF5+Digmg5rOhx8+DlYUFra
w8DRzz2JzmAokCAm4jdSJkwbfHwC+NSyXviD8T7qPS/YejUIZS4i8luzUFcO/aWxLngLob854ORr
R4ZvN60q7rB8L853h0CPc3R3adUn+KvuiYyQNuk8xKCbqs6H91+aGgaqjDDUlbLvA2BKr1dG/VZ7
3dNoDuIqGj5U4kfkto4QWYfhXiLDOSYdNzdSx2tKNqpyvF1yVvUGFf74YA9KZ3vXGh0+15AU1jTr
vExxfgZ2rr4K/qpZm/J+6rXbcIuuRUUPyC3NWblEl+nVTDchdSvoKRfl+mn+N/fBRyAa62YAv4ki
d4jh0GNfZFNC0po1NYQzWJWD68NRN2H+zOo3VVn1Vldx6JzRyqOUjP6zFtSVtR7g2NPjvM50nj4j
4W5xkB3jY7JdfXC7NFINpQQl6e3Za2rbQNQ79GXerfjOWACKmu9mdoKJ9LTj+4hKSjLqojA4YH1Z
XwDTD5Y3ekFN+I5cxk/U7RdGwin3T6Y3sJ/ZCAhFy+yb+Bv/HresnsJ7KIOMl5zjYcjpD1G9HmES
q5dF/Gsz2P9a9jegkZtpsJLHHccTLB9xgxkUW+x08Nu7tY0lTKQ4BhGFC6hWNL1OlFBI70gGjDs/
9rm4wqavL9jQPyo4OgZsQeKd+pwSTBUYZMe19/XIORhHRyErXIEzVaBSccXcsSEu/+DAG2Ny3XB1
c5n6eqXlfbUohy0jCBlNoVKEL3DuKNH+i7eWse/NqIYlndJB5vrQsck3B6xf+Ng5Z6RD2NupbHRt
Eu0DFCgXiEiOYBxu/KJLixb5qqcK76QI/Ma2Js2U6phvHtYlm5Htvpl02D05+vF3wClt0if/0FNF
6cq1wGBWmDCi/MbkiolvMVdEhifLWkybUYPR2eR6jU7MJ+FKeEzJiiIiVkYPd9MqPfehbG35owlE
r0Lj8CknEccrXky2Ny8e3etKVioHH+LP++6NMr7NjPlzvLxxzdH9cZKQ5nDq7yDfC7LenPHOpOH4
a+hR7z12LnplLGPNxUAk9YwKcmEEPsPJMmYXS/76ZZSVxS8gvd7isDhY0k5QQjLK+bQNxCvYzwWD
1y6mRHUN5+m5h14ji87PqKfvOt6A+eU6KlttaKeAXOgaHegmhbCX+R0HDMOTMwXl3NQMz3AK4bAk
B40SEHPN9el7GZcYOxCGcHwnbKhqDIEdR1wIokTbS5QHBv2IMLg0dJnjbAvzSB7MQ+REzc6lzH4b
V1n+W5SbmJWJ0GNHswFZMI2l9naf5IYqEcu/0z1SaCyptnaMZ8UebPJA/qOOmgJ7VC+QDrWRhdGD
pB7bFcYKkCgIr73RoSIBpxtFQqWgq0W8JSBM1OxxGdO9xYJlUj9IZurKwp4txSXSTwVhQWcok8wS
q7S5rilAJ5TCg6IQs4F4DYsPIlmQbWqocTh2R0A0w0jkHm+LD7VYpFPp3+5G0PKC5D9DIvxoFkAx
vIeZdpatq97QsjnN5x+Kv4EWqc93RvLkQ4CTX8KSbxopw3pAYyvA3mBhdULf5tKckY+TOwpVxxGa
3hHaQG/HCK1ZJXaOfI3wpHUbVkfMAr/lZQW1HPMWvP/KO9Lvpr8xQsIWP6PHMqXtjRr6sgZNLgxJ
qCOJD69TFFv7p0nFVxyQS9L8cTtNBEC1AZf9GpliRpawBNO6Uvud2AM6ygqk+80qA1t/Q129bECL
0HZ8g0NLZa0jf1c8geyyLPfR0xE+MTb6yCwbqIWS2/i0R+WBcSO7hZ1JAaQej3ZnY/eq4mmChqkB
RnRHA/uL1U0a7gRybj9fs0iHzDIPIZTOrVc9Q0sYbGvTnNY3dKmbkkvW+R/SoPgabZ1BCuBthijg
duPy8BgHpbyz4jbxL42UJ3h/tOzrNsVh6AUXLX3UybL5Aai39LGz+3kzsTqIWnlaG4fFK4cUSoKV
gjFlzcD82i/WtyPVE+njcyYqgmVmwte5P+PETKDegruPQ+GEegE4Qf7hmCizRRSlR9oXG7il3rZc
PEuf9zxq0vxtYMXVaZ1sD5ZqedViGLgrvuZTD3nXN2jxZnhEyk5/5bY7YVHv5Wtz6YuRsAnQWw5J
Ghbgv2Qzt1CKxGXl+IzJSWn4hsBgJtRzmcKP+x+wdWXq6d/NCy3opubgpuTco/O+zqujpWR6yUVC
bd1uttiag9kZWzSS6ZUJC2WrO0acsFbxG367kA1vbF6HRqvvgPmdc5SSx2LjPPYO7f3sGpimwoLp
4pDIV1AvpdPlY3qyP/F9JHnE88haHwTK5A8/xl3JwApCiKppPRwk3YTFBrqlMALLfdt/BeuSeB7Y
kDboMhulkS68lzLjlK6ScWNWulw+NpXx4JCa2iTH2bp9oK1fXgbDq1TNtJedZVpcCtvWkHOr1CpY
4AfgXzZs20GT+D94pRhFP9nVPXjikNGuavAE6JOrizaUpYMY30yG+VSbPLH+5YaaDt2CIaRIqqLK
fU6ReoiW5teDYkGj8Tc3wQcA5rXmB/jbb2tHkYLiIRPbBHWhMaNBrt/22SqeKMFRvhdT9Lxz1g9L
uW/CQCkCh0KrhMGUyDNTjkpLNJuvP3eQ8QkXAr6XdXeQDbXsCLXFajq6qwG6rGAJVEfJsX7lpLfC
N3QN47SAJ1uRyt/WjxVWEJsWvDi3uEJm1p8mQHehjXs03MktRtvRLhYEQKo8We9t+c9NuNLx4YTj
UH9TgiUqtWO0UFDL0hakX2WCbk8IYKk2CqJbapbRPNJjqRiog6oySgd9NjofxAyfq+/HkgEF4lMx
y1jKqFue34PJKHuIarjkNO9Ik1MZBUDxpxKHgRzdq1hGuryAnQwkFynOzwoRTRuFxCce9qVycUQy
KOswvvGHKUHlQwLkdy9qRvcOg2BN7ccqD+nxVu87MDWYMn6cGZgr8oWzyJZDm0pzGrlSVq88toiK
7PdMLOn+r3Gbqcb9yVhSThvMrCjIP30km+BRmIQb0tu2rsoC6MN2UyOangAYU7yDkPoL/uzsofwV
z6KDguZJoI7zK1My4fc/YfWymw5OXL6zDrsLNcTIxKzxK4iy4loCI3TKrooq/E14D9QMn/09objZ
AokplzvHnNUhisrd330XgIgecNX0gO+L/NT57lNELRhPoA5sM11qCuH9Y+n1qaCzO/qIIVeGB6NB
nOCH69/929VS4I3nVDsJg3bIM4OxfFDl19UtlwyXOmLZghGd06H6uD/47NFPPIQbCk4SvgW49k0e
awb+HZtE/Ekk0WujZbzL1yculZ2A4rvZbeGZhqFO6ajvrBJMN6HELBeSkVyQiYzJ0Cvel8JH1ax/
CglLwObIVQEyYT08fh7tW0R52mReyWYIy5qeYEcEzNk6KssqeE/6PdU8bzck3Jt/8wnKSN/jNvJS
10OdfubwKGz2IRSuaCSm6IQ5yH3e42f2OXzFZxZTyVlcmctJkX6D/igwTQlshQJsr18eyUzx2k7J
i2bqkbSkCLSKlF/U2ZmmVuuyvpy7Z670rArQs5LKT4bPu8Nq34oS+AVdlahMEdtzj6a4lmG+5Z+u
S+zskXGOA4Kpq6dtdEyO5fSkvoKsCCBLabw3Np4WSCnmxcFX54dEgRbgrgIkQnIez3tl/enTj1bw
3pgO22xuP9bAEnwJ5x7N9ue8pf4DcDSufXxJ67TczJfblPvslYWmUr0+i1mIC8U0CPAgFX2YvRrm
pMtboSwStFYJ6j1xDlRs8c6M2xYp8M4MOHNguwaEnLfR6Inp0rQrFhCB4Xw3W9rwVfcXIzZLFb+1
C4YB3Rf+HUC2DUlBLGISYlU+kOQmNkVVMHXGxe6YZ312K3WAd9um6ll9EWQAr5i476sqYm8vdG8O
SKrlt+HNw18dYXAd1xjC8uVLby0xEyLPzt2QtIpXLlK4GsHYEW905AqWalCUuSjGz8Q+lx8/nU+n
/AwfWFdYmr6T2rNNXiVFT2h6AYEH5O5a1936QQi12NI/o+tKd46OQMk0ywmP9oHPxqEdCfybrkIY
C0LXQ7Ce+GG3EdhcsnlB7bHQWWC7qMtsk5X+OMg3ZBa4WJ1pHJR/XPCltoJ58YzZp213p2SyqCgv
2+6O07epo5apQh3PzlEPsbFtpHBIcquCYQM3dQHMcW1y8Y8kI6MXgnM1zLaGmSXat40gUOAmuOuD
uhueierp6tJl21EFLjHUcayxr7C8rtQvV6oXsK8/fuLHw+zGUf5rITuhv+eglSD9bq5XTVM3/rA3
lsjfCYfwWcQTQH5fyWj5vi1YlOIfnZ6uYBYTbIVYSNES5PANBUeOFqxB7vMyIoOC8MGop3lQrSa7
GlhsDkT/r9TUl7FzTdZfR2VcXtJxj1Y4DzMWcwS8fOLY4YP4Y2A912o3jbL6jvodP27isjy7MG9Y
ukHjibsb99CDzcp35XSy6epkoO+H1YOU3tVfQ2aPgryOZWVFcaoe3ybRNvttrTJqVdpx6aWAbKPq
6zOKjnvzhEidTWV5KTvnr/+0cLHOE1u0zuRMrUDZ73akiQyO2CfLHSreMNe0tNpXetAO9Kd8ni3I
v8/W5llrLq3yznGibltLrkiE0uNNEcqve+j3rN1MkUXmVLzHzsDEhns0+JmBd/7fvqeB9vUdI0Nc
vJILcH3T2ZuyJRhm/ZO+FYQqDc7MQWFuB+HGFERAk3wlYwHuBbpAJpN0caIc/zFTPeYF3mjANzY3
xt+vPCfNhtrjtt6BN23wlmPsUMb+Gp7SaRP379lP3Gt6HQuj2NF2FXnDwap6RTVJDKWrGqd6pTxK
k0o4CVmYymt72tSVxzsYYsJ1D+MBOwoBy7X0F/0t7b7vuewRpwUpUCSoXpEUKxfjRAmbtIID6Nqy
M5CItSbpKx6yeQM6Qznq8D7Nw1bVueuQ8gRNrZZzV+raZXrdj8VnhtycjSyFeVwpBe0Kasg28wOb
EDG+7aenjThB3hsfubfaHuQmusPT1mG1GG07BA4zoRPKWalL4BTvLK7BlpkqeH0QSoAaxVQKdaNJ
Bw3WyXD27GoSwrbuT6qpODwZkLCYmdiXGyYehvxxCeOhqRtYxEnrx8HFKMeof3cbBrIeGjpVV0OC
4IlIzCmw1xZchJHxSVWOO0TpQgkhaiJpQZCaJXNaCsk5SYNf79t29UarEpJge/6jB/gYVkp5shHY
YLdLnWWjVTJpqUnJWlB6SrIMv+KiS/XfjzSaRkAXJlOoPMFXGK/r3rkkAs30PJj+iyDgPLsCsgEw
JcZutfePU4Y+39pMT4xNZqccqcxb1TKWbi3s+OZYqiUV9oKUAFPXWuvWREYWWsLpJ0q/t425r/na
5mM81fJG5SKOVAaDpWuoVLR3L9C9+jtzUVQ7k3H2vHwZ6axeHusmuF0F8IKx+mHViGM0rfACugQi
fOpg9jNUx+2QE4K4q6AT1ySJFN1pjyLt1K66dcdAS9wKuDASvegL2Mby7xD5yDt522Ez+yMJ268O
cVW/RrNXjcJknLXZ6OLP5148W3Cx7651uJfiAwup3h4wDTlUoKddBucx60/2WFJiIo74YiE6IPXa
LnS8ipEVv02PU1Ol/dns6XwKau2p7vqr0LE55vi8k7pGlffyIashVFc3ooQTOil1dawBY3Qm5Nnk
oG6JHNzSTbe/sdeQKjE+1adFhMa69k5LD/AkC7UBllAsmdCvVvZF6QL0INxjhf7fjpG3Un+1gqgv
awcWA9IswfTSb+pJxqCrsaLHqjfiYwD6fnI9aXBW/T+0s0Jh1qNyyFTNT4Gu9wiJ6d+OMbo3y1kU
lLiniazfCfNHPAwrvxz9ASgR+i/pU/MoUQj7kjAA7zOiwE9/O5gIsOeTmgwr8T1z67hvuRNC91Yo
qTbJ5fz//h83StrwQHDoVTx/9mCCfEmCAMMwjLwYgc3vc9Mx/I5xYt0raPnjVCiPCOaD3qgVekip
poyTOh5mM1cpwiV7bJc+WEU7XWl/2U6OsF3dhq5JazwcCjQt0OwHHoUy041aYmRPgRqapC24pUnw
F7N32rReCguCvv6+Dg2H292dyXYMOdP0ZtJxzxG5sx6By4N/EnfrVL3KcE9UeofXhEApI0nPWDLv
ZyT5hS4+BNVnUgo1qG0EvlTk896cSZarltG1WXDWA1RzxOyqJp0kcjH1az0leeu7Y5+EwXK3m9/p
XkhtVE66N56KyYcN4ivb8618VTOYkSVTv39Wff8DiKUO+TA32aXXYXuq7mmWFkTFHosOkzoGoczp
VJZ1+5M4yUla9BSuKKWswGgoFWt18jX5MbiHej8jNvmkRJtatF2eH01ypnCpb/5cj1F02it+kSe2
iZwJTmZHGXeG6+YM17PRFW536KCl38JovsHArBE3E2Llw2gKXAKMUnHLyJOtd+lCsl5TjviCJDYK
eUvtFx3scvOui0oTOQPA4RBmPU9OtnS9ZYJ0542XhDHk+lrlVq8ywvzlI1inFz4V8AlN3UEzWT+1
iQBvDssRBelCdh2YhsxYlKgwiB3SPwz29vCNSrjb2dx9Nb+VvSuJ9Ylghdybouys+5Ir97zEtK/O
TfZnvAjrSNW2oSXUvb01jfN0hP/SmWK68mwe+OR19O41F4YOIEm+TZImFu7OPer5PT3zKyBYMLu7
eva+72wqeSVI4GUGXRzkyLUz0et/Y+wLUwjEEdehoTd+G4FoTqpJkUiIR12WW6dfwpcBJso5zRmB
IIENm534Hh43rpOY1LQfN/YuUl4GWRRAPP9Jxwr8kSXxNsK5gkqsioBWQt1GI3gJG0gPYLkEObLZ
7fp5rKfXJNW1VJz77UTOyuIGQXE67vd2U0OiOdyGHdFTqsIe8xvi7aQcOX0BE8sh4LXTq+gvGA9i
HA2ws7Nkdj7sUEVct3B1qq1sfDtLorf6WP6OhSbMpVP6OdkGAr2ppLz1rnjsnaedfdTWEM00PDhb
WqE7+2urptNI9i1K3SKrRIWNC67bErtgFIdCm1y4C8nEPP5sT8azirhzmlyLrfPKlNz+6y8nQydv
dXAhWkFS1CQ8tSRxK0rdEqs0LCgR0bMcg5M07V3sjjTOAXNimvU1WTTLoPdieygVVYcOGozePwiT
v5gZlqzsFS4sDVs7oOmQ0QEYOnNPef/RNTmVukvbYAFhLUszh55HzY7OIgda75M0I9ECsmY/6e+N
VDAg/0uU9zGwBfHdzZOkJAwbdPl2xDSehl89B8Pl+vj/XDO38rGsSzwCN3DPv7eAHpPiQwfyNeQq
ECcskvHpvVfju3BAa0DSNXdTttuUaUIyh/i7aBRKZhz4y47JllNrb03iow+O4pkkcrIo7wxeyh3P
4bW2NpkTBpQdlWzpNTtf1SmKDbNNPW2vKJeZKy/qfkZdJULIsGoQxSIeiZeT4rNp0IjCeGWTFszL
1CvuP5QYGmuvE9nPBYTXCWvjkt0mX2Axlf38AZhwdUW1GJaCtf8vzxKnKiW/wNqiHv7M1Gw7a7fM
OrV4t0eigKzwO9vcz/yFg2DbE8Yzd/gHhtfTMf4NGMfoXyGHJEcwQYQzos/Jx8rzo3OxZgQesOkU
uyNjj4KHJ2805liq1iSl3tjoC/9IrjErHOrC5pDUvIQfHtBnrA2vP+2p0fzAfs5KrKx5SwzB/wl1
gbMTYpntYqzhHWOZlyFDh3mhq3wO+taThFnIdPEO+idCP6/V5g8092GzlcRhdF1Z5KBJLrfuGqLA
InD+woYQODFG9XBx4NQz5SOZJN0NmOjqPEMgLjOmn5M+xcC4uFPBKwDWKxbO9r68FB6x7+ndLbhE
cb7SumT7KYiqnX4RaD2QLreJZEo7hRV0rHjI38hU/06YR1gd2QTwyk1V2WlQweHZaBpBRfSgn/c9
5syMOS/DiQrDOF3XD1N7Dq2Qfn2m5uPd038N2JSqfjaC1s0MiQn82LEDgV/Ziu8kZMakGL9ih1Jj
3h49D55xTFUgbGLhIaFe79E7X7ZqmGKf4G3rE++c/T0o6fenBqa/34IA0J0aM1fyOX9bBUCjtRdF
O9y2d1fFjJ6FoUWkc1J9I0rEBBRhwoNrEbqRxr3LC1JpjFEoWl9tj/gE+myCVIPmJ9DxMTx2yGl5
n9CqwNMZvSuIcK+YrvpTfbKR7jMvmqV+WjGyFZ8231MEADc44HSpp1aENjENyy4FiYJ/8FRiuBjd
5zN9CCO3QkAfk5D0z6c//Iqx5ZQAUqgw7PjEQFDKkpfcmDW3nkZPJ04PUGyqbEGms2CE4qoHIayi
CCoEMtqOx0j9ydj0ksJ4l33IwG0PkizBD+O2fwdPr3TW6Oks8K0clN+OktqzSb5BZuFNXmaZSzws
/reCFpXjjJc56XpYnV0PXrjAAVc6Keu7omhT8EMJG+WATSLS3n+KTwMA1w+MlM0FqEEgVSq6Hv05
Qyt+R5ML5Mi9kvdRmUVJe3YqTRe2QEf+ey8hYcHaAYJaGiRGqMBx5m9fPqpxzxKR54mEXDFbyruK
jf5tnuvRrmRJBLvFibQUF4mLjrkEPwb2UA0h2vYYb3/0nMVB1QWw2nK5NIpdhOsofUrUgmOakz+T
61KCAReuoQ8itS6VNcF46o4VfsT5ZHHMNXw+dyPQTCBVx/v7tDD6MybjHe6eyPpFEill5NIstCLu
X5uPgAf4tVM2Yve9RN98mSVOlSiszlByPPt7EH7xRt3SbYYfoyXicrBGkEkXZHdVtT8BuGVbudPL
AEih1jecNu5zH9cflFID2d6EKbt57M2UCPE/k5/WyiVkacPPPiBkbkbCPaRIo4LFkZMfH4Eu0z1D
rz6JGwRDisnDZMBVmk2CKSrYiIDZjXHmfEEv7/mhT7GLs5uuUwifEDLhNLMJHboM/5g2vZdjSb+K
7dW6VgMzc5wzH7hAnC2rmC+VtfsTI19IdGNsXa1b2atMCBxsz74FtatBvFYnoUQLCQQWJnc5xKTZ
ms+Kde66G5si1fwVSQabcmIXAaTqHDPfOSjWztCCl/jc3cuJlIdLmSVdt0gpDc1KC1td6i7g6y/t
w+7xk+m7Wz3bTpV/wjUJl8NtO1we/7upGWzFnjHuXMI+WWBJFWxLOMfY4RDGmTu/UVPA7OKRifOX
PwerRiTdcumJyRIxA3ygqxRIlbCJh/aSEdUA1m24r1MkAkp9IW9xFjJjtd1CW6MM7/hzZIXOWJ9w
Tx2gvFJ/ftMz7KtN5ErdmGdRuI9mrVQm9enNpL0ztyDSxEvYgmMeM2uYuAxrf93A19feIfjAGWFz
hVkORWtkprk/mJC/e8H2WhdOK5P53lY6pruEqAP6tiawIXEfiuOaU81QP+E6mOlNK9f4PAh1QwUq
HROmwKzfLCMptTehzocM6AaN5Bd0tIx8xthH/qQVL6bYfWeEY6W+NRnF1qW/uw7pv1M2NDDxex5i
ccEOKsHC1TEGW2WqV4C97ZYKbQAFRRE1xnP6XYE0ttNacC48W7aeuua13kelvAvxEAJXvlUt96Ib
3DgRSs8F+3Rz5BIF2va+SGqSFXPiceirN3shqmJa5eT0emNkbuuY5ky0zwMgiS5fTuPwTkvMOVfs
iGiTHI5Dd8KUIPgQDPdetRfhxxKwD+MfvUgIfs4kSNipbnEHvIUaTFWfP07okpdvo8uoJIUs6Dpz
VY8bBLXZSeIfufCJo6BjFCzS4MxEYpd6cHKiymJfv8A/fsBi0qMEDXWquLvA/4iSXummlRMXapPq
OcY6ZZ9TFPjJEuFICE+j1tRnHnFQCnh/hjwYFCndof3yap4t7/4fRStM5Iym060ZMDsEgsgvGpVd
xb9uYk6qt25hl19b37Q6OSCteYoNOK7QAXiX7w2YEEpqsGatSIdqgiiXsi8NTWdBnP1fBd1tpdQo
D45fPLc5zy4XHBu3GxVGM36jqjSv/3XQYwWvX5AtI3aFE7Cc8qVzKNPtphjdwKlWjBnoDJ//3y8F
2S1Y2nQqsbfz34dfv3eHEQAwaCJpCpHnVV4SRnSpxtGzqucnYdAt1cszdeT/kQXtVDmeRRCQ/Pt7
lLVSWg/xRmCgTstMA2HAWRuJrB/5l7k8n/05xSn5pRQnj/VGmFuJ5KFjoQyLplC8zvKvPj37gnlo
Z+SwJIRiXWQRtxq3flbWQ4Gs//NcMWIN+sd/1sHXoLla4vEIReEj3oiy3qQkFQbhDKDJsZ6xQk4a
DSaP1Qov07wQfozj+xZIlZ8NlB8swxVlHDMjic+pXFhBH+0idtIxYFsWK9gEnRFnUvp6Espbt6AG
esHqvvb+NR4Kd2Xm/yM8S3l7DHLAdrVJYARqufQGjsD4GxJtLNlRrLoxbQUVDuQGXVE8IDW7k8Pr
xyqT45r6s4mg89N80VcwO9Y+/nd4XavtAbDZpG98dHg159PurGZtB5mzLUKdopzjgJkEDzZlHJEm
bmrAhJJUD2DagbOeBOOmHobZ8Q8aslSSw27JJoj7SaYSZfQAEAbGJr15pM5g4gZsqVyHKuOqVOQJ
3PeQ2h10+9nMkxZ3A2ysczzCz8Nqo6thtDp2c4Z1EKPAjpwRcvftsGI3F86g/V9nDfn0kn5P+nor
t1ZydBWTq+XtV9g2tx8bTYLypOMUHpZradG0rQ1/7yY5vtManKFA4bWYHPTwgLsO6+9g0MVt71eT
29EFwrBm+UIwNw/ypaP2nN+7Skj9e9GpexPMI1719lorX+GuVSOW5XUdNeflno4FaKPWLMxXGSuw
UTWWtylbDCykSGRsEuv9kxV261bdqrW9T9cShP2ruA9bx4WOOSxHTPEJuxD19PXagBk5Ax8BJSzh
9eewUtiltHG17/yfr8/Sr9rUxho2M35u/O4EaNORF7PD6WLsXIBFKzLZQnpfgVNW8iZItBhKHxo5
LtMAnqAvgqbta02rBWQ0P8AQmml6p6UpA7pr5WMNPwlcgOlQioXZtv9U11KcMh1Kw9n/wRE0urAN
Z++Je6vmHuRj9vH/1wZe4Gh9O52Xzs+zdqBlspnb0Z9+pMHXwUtZAGlLPStfxINM36g3agCLo7Rq
ND7ZWFfMQnGlMY74iymEkvFICVO8sIhLljESzT4iL3NiLg2qAzvz0O6FbGt64v7edpXdUpaYrgWf
xh0HTTzwCWdwthMkSvivOdIGhhz+MmHMyMAOaB7lDy7NYoN9UdITvok66E8HuNhhnbJrOpCHV84+
o57TnGyFPIdEZh4VUBgYniQRY32EHgTOZi2SsAunbFjIDHtXGOEEhWs2HqCGz7XbCq1ot3lPRgoo
p2jAF44l234twpglrYZssYOkOulKSXnBVblta2nvXWd5OP4BuEZ9NV4p9oL1wTOdsgc1lli/jQH3
/SQn+Wuue/3brZA5sQBQtdnYm2vd2S25yvRriYDU4sPJFbLyu9PLlALdbuYrm8yX6xtlmR0Dvmzu
yzv/KD9QvX9sqlqC3aiA1ARSYCn/fwoAPaTXhot0XdQLrN9TkuVeLIb8Rpbm/PeVWF6ryJoPlQSS
WCU3IikXYBhfajpgcuXYAnZw1OonjYiobMbkbJGKPxDj8yaHRc6iMjwRAyJIhZ+jwJT1GGD8sN1a
uAp8cQkuJOAcgrDWm6Svy2ehnkd8PMfNSYmYrPUnTonUNGLGF/GWRuRhyLyPisRlzbqk/lBSzBnV
5Z+ekKrHTLOs6bqV+6yw5LnnTEPmfuGVGzRnyPoXTTIgHaH3HvQuZiZCntMyDLhREAXSiZderHc8
tbDLuueLpuHlDb+e1Nlb5ar4HuhxMAt9VGIHEL6mhufud9NuiPuqJuZNv4tYX66NjYEHKlYcbBUl
lc/TwR0nKKW19N41G7QjPOoYaIM4OssNzVo9rXRNNd0cYFatU86nqVwssx5gTFGnO0X3aOlv63Hf
uBI3RmIewcagssGTYLdVosB4F7rUQGqIkai5Zmb43w6qow+F4eWWnHkw5y2ufM9pr5EdqirQnqsl
XRUMJDirqECx+hEtoYIpMupNMNIrkGJgnraTG70BGCAwg8Cb7ccAPmA4NfX9A341eScFofcg2YQH
TtjJym/e0S5Rvv2vfBlLpER8eI1zrLmtuuo4F0mdEk9uFcezZRtuySeOGAJlq9er4gH7qjuF8Ghc
PcbDZkorHAkzVMd2MTeuH9/rZfFzsdwUlL703Z6F2Jvkhkf6wME6vo0lMLxR+5z6f3Yj+UguE+uL
H31zWJ/ctpX/YEIhjwzsFhb6Hn2ByOe4gwbwKgnkiMIFq+tfkZ54ZGY3wGV/g9MeC7VAGCRq5jf3
DkmPo/HXaUNmHXJ9X0mRiEhMwExhxQFH2FXSF76wJ/a3EVNwobrmR69aYrbvidRxdf5z92dLlKzU
8TQ8D6iHHbX1/MdczZiYgZtviDUxZ5tFg0qbf9Tvz4DIJ4PodzSSFG9RmzXNqtekwG3MiJEesfYg
vsroGVOP3I/AEDMZJ0kKa7LEvQ6A/LI9xXGqbhwUG/umbH1xmnrn4bN46ilXDUSWwLXrwutRVeaI
YkZ5EOt4CKU7T05l6GvSW00K32M9ZBmOJVSxe+kwQXfR8i1W/5YHJaKwGof6gIYkEWACkwMqBF5b
0TtsyRWK5Qq6RcJZoo+4hozs71sK8Vespp2BZrMahqJDkLbYg8Yz+c5v7o/8cg4z8rnOrw85BKxa
2hhaFmox6b+Qbemyx0mgLOcUMRZyBHeU7v2RckOOMI3RxEOu7LIve1srmggjEOG+fzf5YQgVSpPw
yT6DSP25svwbyYGFoBwb18hchhuJyhHctlufxvc2UsWj447PhGerKZv6a1WSlT/fnOUJlBXAFqbG
ZZGd4S1usV/QNzTrGXDNpS9VyYaAN87pPM2vfnpb3/mCu3WMOeDgecGBTL+ROvNQd/TQjNlMOP13
qcxLSqtyvTs+yaDc07rlpAYGOmfu+q844Mqdt6qoULDfV9dQPDbop3vqcoM+DSL+lvLKKHFKfzs6
W57xuOk/eUBtRMT27HCUSU/1qFUD4L5lKDd8Xqd1ivc5kIQl8j93POLhfDcTq8tH3S081rkkRKF1
H/JN9RMgsICRJvw9r6CuCZOC9mFhwR0ZqqYSQpCKVC+7MjD1fsIFpqIoLP/56FTRxVCAYMXrKYm5
XLviUp2e5Y1ihQbP6XUXOKCzGFIsuqarK19HsUSM1RkUsUKss0VCWSYG+qXJZWtTkD+xqBHB416c
lHeOjVEYt2a5iyCiwRryE5e4Tidrz3JpRWRRiW5AnoG+DUc4iWPBulX7+dyWW/Fujx4dr+76gwka
113zMMFrP1Z+SHvDg1yvqBR2De/6w0RGNJHRcM1R1f8rt64OwHlBQWzemRTfeZkusrnf4gnwodeM
VCEcxwUMd+3I2Iow+K/g5LbNS9PJqowVV8pJ0W+vGbJ5qLuh7uXwDxBEalEImyzXbXJkKOu6vjl1
GMHi7PfcN8doJk5t16k2yBlbwz6ImfXLdr1XlNqY9hJZLY+iMt377rG7DYa+7hhf2qZZW8hX+l0L
ipSfRp5cCCk9fiiZ0klrTEKiok1zRF5FhsbE2NYuvMG9N0/PHZMb8WCLtYkSq7enVaNsAPTqFTwJ
3vaUfy0VXc4wejpu0gZA0WdLM5/eHkj9jn4O2OjVqDo85hyKC/xgDCi1DuQucAGRiDRP+GfFQbNw
AKJFv/xnkS5OR6xZjRvTmtb0uFC4UqMYTWrg/btzfiSEiPzqgBEA9wCx3k9DZGv4tafKh/NujOxC
tKXbfvPzSBtVuViFyEAK0617/HzWnTMtMQS5RdgBH36YFOflrypPdbLqHu9joHg4WUYCWamLefKz
5kolx200WkXrXlAg33SgX6YE+cvVcwNksoCDc7gpgsiwb3bSEJDYYaLuV4KrF/wD+9AjriVE+q8v
X+3pJI7+FBjq+26rkiHRbHbgvIRZILgm5UEAs6ZEr6pagC+bRBN6AsJ0RHr/cI+zNLiejkLqHeuf
akqB9GcZDtv4ZqE5HTMgHAgxkIafKMwEwGzw1XnWBwbtcov3Dtt/Cr24CiZaxtdS4Xu6w1uC7C9V
c9Ft0HU1G9iklW3UGbr7eVJ5w0WacJjNd+lPZj8j5IfKRXUS7AQffuKDvpHV8PiKMIUJ4KL0UHuq
TRBeloSKT3ebXff75kSag0KoqwNJcNXQYckyfKPRXfOWE0JfU6vbYd8jY4yky6RsAYw9hB/78+RV
x2h2EVdsVvXGMCyX0tD6csks9vsJQ3X0Tat3s3MIFXhIQdqLzW6FKWgy5m/opstXY58qIqNORGL5
Tmu0CqAT/AE6pTsYqfj6o9vkpfrBl9meIb5pdBkEj9zvN49HJZMs5XdpCuNpYowh9kJjXTCDzK25
ZmkhN6c1m3gBSOkmlpz5a7+mMggTmWFxVoipO/bSVaotJ/xKEBR8XrT2ny/6uFZhT+98rfLPC6yb
btXDK9qqgspf2/2Avtofw6ivN8KePeAiO5Ko0aTheQ31neStR5KgUIGodkikyYycAEs6HQY107TJ
Nqv11aTTRIe8rZZqRC0CB0DkcYK7ptphgLAElNRxQfdyAQUmGoSbECPX5lIWBKbJzW0/uqmJUn72
GMGfuF2bDk/uTa+qNioTSe3sKKCg5oWO+uuq5CrwLCb17Zz0OFU5yn+qnQdxDfrAY47wXvZrKBkN
+1s7g/OdSSloWFfc3b/edL1/KwB7wlg95q8gTlZ2k1OUXLsJRDpkaTFMac65SC4D5gxclr8tKhrb
KRKstzTxTUni6UtvkkNv5I0lbtLEJhEj0BjfbAw2cb6w/TBFLdhr8pNGJaxYrpairAqwQG2h6Ne3
7QHzLEhWXBjTV503BWUcdh0G6iNC5VIm0YMNvlJOL8fJlAklyyN/kIlAGyV48QWZwPxuU+5XVwNT
8kxFXPfI0bX7iy9+AuosbupHEfcLLyH+c/ksjKrADHxGz+OFeYPikwTiuj89iSAxdR2Z16iHiKIY
8PSph7UbWGtG8eMWky7XdBI5v+n+PQhktcWxRwwEXMRcjlEmrOQiuQknVNdWphkjh8lp3FR1PhND
ivCp2hQO0glmus/wDCTiuveOV9eoq6IAEp/matqNEiq8CJ0keH03wD2wQCN17neyULW8eTbvfnPM
aRIob4q50+3D6RwF98fj9AzQ0Zdy8FqyIoXqASOlmKdyB2yDRw7ZYWmH9ziWN0jULZ5Th0p5FUrK
jPrzLYC3w55t1QoZuE40tt7dj46DQExzESmfnI+xIxWuJ1eSWRohBf2rS4swpWTjuJPQxa9kajSL
rqIBo4mPLvrIJ0uumxQRKx9yosS3WbimDTxZwzEEFZawSkazv/GTa2IDE2DbtmS71ubSLhp+vMNM
oUoYoODKygdMYggsYbfEgzhPP04kLv8d9babiMfLcvOcZUbQx6ZaihQqdjyUFEEZoHx2kGTHfJ+b
XLygqbOugp3mhXwMmgx88YbktAgtWl1fL77DaUj8WE1NJC6BO0I7PyCEIYQn9gObX9uZCMlARt6/
QhYUW6hjloSMg5pEitb8iUwTxHk8X16xz4ui3kUrTS4DEjcemRQzuwLfvhWSdJbI3y5btcwjfBk+
XS7AzR9iGdFcO6h5TFyX0Ge5xBPVSiA+blE3V1YdbHuk89h2nPaCKd764Aj8c8jqh2vyyZzDwIao
MAbXDauq0vLkTC3fjjA1WMcXOc19zn+8ARIrLn2unsLPzmKRZL6G3x0LhDqKlc7GTBVoPzneefPH
ZT8B8WPBbKlxks60YRFCUg3N4S1yp3SZWLwgcE1kv3JPYYj9OjhDXDxk6xQmQuOPSgkwGFY0drKR
ziD8eFy91wBChcQfqOPqfqMJJaXvC255uvRX4WaGeRcBCDzBMgE5WiduTsK4L8a1wShyuKdFR/TT
klwX6DQi4Aj0eWoOpS0SObbiLxD7RByqS+RfxWj/ngyvZaqrymxyCKNaDU8BCx2WvEtBtx5apopr
lH+ihQ86gxQdL9KfbQ3kZoFEzwp30Pb5KXUziFMxWQXqeb5kKf4By4vdba18civSt0c1scgqVwVy
N/9JQceZJeX88xpbzMoJ2nFTg9VFx7P+M622gWWTIeBCDhklbupxBMrX5iArTI4dj4lGdWoh4m4k
fu+jwUt1bsQguoWKW6aynAzDOyZWKR21pLDYSEQZa4ZcQIL2aBoT+2JJ5jjzkmONzSkKl1an2dqM
B7hvWkMUH5ikXkyyvX0fQPTuDdKjfdXSGQdwOa+CByI9ObEVWSusMDvg/rI/3CdUegdsSJdYt1F8
9b7qXTMNK/jz2uVB2i8P2ORrS+7GFjxYS2h0jRJ+Ca/zXuRWka4lt5osuJrBAKaBdesJC5ZMl55M
fuUwoqziGkyc5x52eV5FD6t21qjoSBLEk9oc4eIxUhGOAL9dtTYnFnZirKrkl15JaeM0PgT1Z9Bu
NfJ5Ju582NqrFYzFtwinb4rFOTdGYT1dQylJ+P5DlsQUnNba4TcpOgXJKZ/QWwnoJtToJZIvRgDl
BuUt1gRUeh68vJvmg2V3O5jhKMOmYG7WrCz7ytOo2p/O0ydiiMjCTEpRV/LlNNzUYS4vxnd/pY5N
6h5xgLcedMUC/JROwxxIAFdJiJPA6HyGGKBJzoE/Q2dpr5Ppt2pZZAxMURNzDxtTnFqa893yOJyQ
lTG9dsuvGm+qyPvwJtfJXZa1K2z1N8lFqiudUx7vo6Bo2WECWdBjxhH9sq+JHxH08KokuPPD8WpK
T555hYQvfNvM1vmJhXe8RooYXx8gIAetN+VlIXYR0jR+/WzdHRPME+9UMhu5B0HCQSiOtT2od5pR
6jwlTzx5ItjJ/WDcqiI0mN6X74/RjhmHUqxwN29a2aavdpexerZdvOcJaK4di02uB1PdUdmN4Paj
KHK5tkc8ttWlpQPKOkAL43x7cde9DjpYsTgsq07P51iBW+egrcS9zAL0XWOMAy9F9TPTTtIQV1YE
W1sEgbJCtkRg1SHnFw7dJvCA8m0UFi6hn8CZ2G5NS1XZGZZ1jtCkbSV2/81MC8/+FnOCRtID0pFk
iHq7YJ7rcCjVCtZ7xjWq/bkECPKVxdyGfDvdSuAIshdu51DzM+sBVOWKiZIEE/iWMGCcV6NtXDID
AZRSOjjR2Uw/dL4HCTkBKqb+xw/rhN/HFiuuWZ1AauQjhvla93szIn/hX9fZEChS2uHmiSP4nrDK
pRPryPJ83xDkBF40wYWirlTDgChK99z0a0zW9wlL9svAgGPnbbREus9tbdhTNVyL64F66eyIkNeY
NbUuxxtOmVFQckd0PzPds152nrIi0CJ90AMozHCJouO2lry7JxXO0uBie3Ok4EgPGkd/+oG4QwXY
pRjCkfJR257FgfmZg34FpEQOLNfMhFd//jzr4UhpOoRP8AHRP/OGkuDFY6JQBmAB5oaeCgVeCax9
VZYH1vz7JY5LSNLh/+356yTkmIhPifXEfNRLD+eNu30G3TYQIF4JMctezBK8ePIMiP7qGx2DALw6
7lNAJte/7SIjn6yZ1Hqmdv1TZZnoW/kph1ppUPcDsu+YZyxtKgMb+eZlSOMjF5+/C3O616iZ3h7I
dAmb+jJBUiE/tQJpEcjsWvr7FGJpzi+RNuKsjnuwwYlNmzvPXHnv4BMGksVjFCUKPmpa8T84gugO
weZdIHFD47dDnEjBISj8CzqrWXEBrbv7sIZnWMpvmPhgA4FocKbU+gAuoJmv2SOFFJ2Xia0Pn9lb
O88/Nw6XnyacSViEXKW0Ry/vclcJH7+95oy/fax6iinYMyqawwHHxAZFQJkx7OV+NEzBdL96myX3
Weds4B4j5G6rRRkVFYW9B/ZPfRvhgef39Xw15LuwqTDxzFS0WqTm4VxT67QxEQLpEDH3SLyocRn7
kNJAQzeUa0pLYm7xWiI+C6bWpS+2U1jFDfBOmI/X5TQPOkc20IaTIr1ZaXxFq+yx5QGnapyDUM3e
kK3phC6FyNDSQiRulWEAc1LfDsq9y6lzU/EQtuvm66T//CeS/wELOof31DJNf+V3Etq3qjbQjR5n
aVuz3li98hH0ccnHSQHQqxnBbb61CXcFUcHQx76Nu0MLlEYxaOrYKLq7kxI6IOzt2fA/vsvfWlBj
bUwyR7zD0APKblO90Fhlx3071DQA9Ky/sxB9ZkTT4jAEG4d4NGO4oBvxZqan3AbIVT86rc5VEk9a
bKviOukShm+K37ndmosTLUXqNWnknTS0h5EF4c1KmWnFtvScg7tXTGu9WXctZedeRaumfkYkHs67
+FqPsY1XWbpwna432PJ9U83kJsMU0V1GgEYnkY6f4KdBX/+y6HQYf4EImYjNHp74Ag5xWI2CwN8K
Ff7YG4xZhWI6KenqWeHuILG37VYIgvFr+AoFrI/2TaBg0H0mTIrePjdMrhF+wbSyeoQ82EFGKs/+
krcmthxKGHNqsWSoRBq5FYiC0KbWMTKlB/8G0Y10riY4GDrffQ/paXcRWKzPglbwTlPEOuQ3uIGW
KN0RfqAHrpbylNqv7QNwxe6COsYycipFiMbRJGdbPcasWCYg0gK+slTSiJLnTJaDl/U6Ipd4tcgU
HAx3OcpJ7uhZP1AcoM+kncP1Rf5kntblgHFn6/N5pcLo1AOtsbTan2NAgVkKXRLcYI7kL/d8gZLe
/gQ/nJQ5TRmba11Y2M0QX8cdI/dLgcJz/gym61Z+44iNzxCgT7eAVhWHNuo20N6H2G5CQb6hK6a8
Rh+zSemTyCSvq3cQgjjq73SvhXwwKiUwI6t/IqOpmyqs9YUg0m6/f0Hsa5KMPZguFYKTTf0MLAWc
fpBqLdMXuUSm/OnkLcmEonimA7Ju7d3xeQLcJsqTCfMK92JGpEcCdFsmJtMMA7y6GVzSHayuL9CI
jpi6s3tB6zApfnzipqEXEmfkv6YqcO09LP58EUgDiT8LDXK8rnXl67dwqLltQNhMZ/7xaQTRyDUl
2jfMyvtw7zDVyWj0DpJPXJAo7EcQsvePycDv6BPSQ8NIlGdq80fq5U0ozvdZqo5vRJn0NCBgdXjs
6rf9Wod1uZ30BLiHTD6/PSZXuaAHZdJpfa1Ao6dnoqqHx9tkz5Gn78mk+d8BPpWb4BMRp4kmsn/M
1m9xEeYI6UOxJFG6RTpURRp8EF/4C9fniry1iE68if4h0mjWNQb0IkNEgiFb/rC0JK5nd/5vsCzD
+FNMGSKKaApvfJiVFNcTC2aktS0pC1UXx0JS+euUXCzcXDHgGF/q+3vteB/0l8KOHNuORGqwVBbS
Ac6L90WMEPORsINLsrri+g9GAYl358dgsAVzsaeN33t43gNyAfElYUjj2j+LQCgCOvpFK0mwgD2m
W4mKILQ10CKBuMP1n527agHWP0EtFA5a3pjDtXGlWzi/wEwtuqr+a7aMA7cNebSTGvFBv291P/50
7b6QgvHhELZnBO/u4WwDOcL0zIX0WYd+Fx+qkmoebgzM20f18cT09f8JEL1vK4vEbhx5v8LkY00W
sEfc/nkjG6+3T//zAUjC5neIA85Y9QTGzg+S6h9gijO/INcszfXpAFeT9KjvVkKNd96s8JVmlnGO
jOgfJh69efmwwx/v1/efQ5Y30uyr91R2/tu3c6YQNeLF29Gk1cCdKltN9x8EK1Cm2Nk9u+gByCOT
C5quZh5aPdFyc7jYZbNMAmkU4VGDqO+yj80CMQP7pxi6vL+uQEZTvDA1kVT9ZdF7nkxOgT3T+/DA
SyCXHuGOLq0Id56tLK6JK/0LSmM2OHHUCDmslkMi1YkgNwPf8YL9alXuuMh+FlzaxEe/UHos4waJ
UnXzMnTW7/s6Nn8S3WA1tUPjxLVd0cVG5QV980zunVtSbreOHg1mSlrlEZjEUv9KYARf+RVZk0sM
KVvJiydcFemaqdAiTLxRk9qBT3a6FsCKzMPDtNEUBQCpx01rLnsvrYNLZTFwbVDwgdw9pnl/s5uH
ec7u1hlLHsdEeOoM6BdPNmR6NpgFpPwGdQFC1+rzz2vSUju5qV9LMErBBrQFUKpR40cJ6WzaulOA
Tf2Ra4SCcoZ1akUU/8y0tMiBeyGJ8jvFlJU36d2Y7Ug+t8dcGm3ue83de0qW2c78t18mgl2+/JVo
9HnZYETqkL8sROy55GzOS8SX/pCrCmY7V07V5tBCIxDSiInHuXV434pLeVDQkPrQnLQDo+T9MdUD
HJu7Wgi/AKOxU9L6uV7J4eWMmBPN+LNotyZoDy5cU3uygkZveTKpKEHUeZ3/m6Sffn0Dxxagxpji
7CeGjitlzyFkP5OIQFa8P/MsRyUKBh8z0f3FEIOR+CISVxQv3G5X6rCc2wKLm+YCS5g/bMryfUZ9
piXtADBmstIWNyOkGvY8wFeGKFQyO6r29foz8AoG8fGHMcAXN4whnicyRXZG1czZyFkxS2eyZTpL
gxAXbCWvuLs7yAHd5Q53AmJVmRy2yQrdq+trLC6LT3EqzATbQwtNZCx0Nnnf910VCX3oNhV50SOQ
y0TQvwsb8G0ybgGtWgzhlrqASddlX4RzpgJCrz1mCNqHDDEPzYnCOCnD2kivc+N+3J9c4GcXoVzC
vqn+HzxEWJi2BIFnD/LcriNFw1qgPaQyTHBPvMxOligeCezsfvThoi9+fGWQQVeTzKTcUQwTIecg
c5bpeEIaPHpSKNwlcSk7F+TV3BqNXv+LPjryvg+Yy2een6J0cK/rmRUTBrKmvlGJAAogxEKVcWGF
UBRdVQHPpVdgDAGD+itXs2SEDftuOPeTtcf/uiG7719QcOi1G2DtZf/1eQdAY0hRZBu6DtUiIBeT
5QIYddaNCWCzOxSpezo4EXI3fQLWo/wccl7Wqq4lAatBmJZZBXKUE2XUGa4je/mklVlfvmxlgKPl
L2yTF630A9ktjTvXpXUHB9K+g5WoopIP90XtNCmcQa14u9IeLOJaoVmfcnd8M1rRpmyUD/NyOhBc
9qfAwbOzjbrDk7QeM94NsbLiJpV5aXZ34ffpCMXPqEl3XsoVol7oPYas+qGcq5NMieiVoCcNbaiy
bW5nSEcNBjEFeDxPJ3sz72qa+A+QSTPKt2zQM9Z5yLQ/z1q4vQF3+oBi2k4CvZd1CRJtXvG1H2mB
qrKv1eCVb9+u+o2WT89qBPeJkLejeqvIPEnqqWAB1C0QkcAxt/0Y2rZWzX8iFBy/qcjeaAFc9Kvc
dXdjDubksEn5NCsPDti9XrKjzsPJ25LldBhBsYGypbGs2ETie+Xa+RdHIeg8YxNdmfi7GixbkKQy
t6rqaLqZ3ZhQ2+/f9+r8CHPWF9Jk6i189LSzrHnFIS8VHDDRnoCJYi8ahjK51LprNtbMXhc3OyCa
gNblrotNwH+YtoN/shxNl01hZ+lnq75GB1djBzZV3em6+UcAGtxSJGx8on5sWNIQ5ElF5Mv0iRZJ
QOXmwAgiGt/wK95FZcF6w6vu391tphSO8RkEcKlyehYLK4ArY4qqSL0YKduj4GfH6OsxFb+aaVvP
yfkJJ0QNMpy+BXbj4jjNPGOYFH+WKCvL2NcTYJV09ud95KcgePAzszGL/pled7uPRYbE/zHS0PmF
+PFlAQvU1m6B9YuRPpVZJ9dlpP3B8MaTohZS87mH81EWOSvMrCb1hRbh5R23T33gbbjeOyL3r5om
v3Dz11qFsxynJGIF5XEedOe7Mx+su1FCZ37bK17lvcq5LFzKu9TLG/EQPA9jOzt446kFe4ANkRNG
Kdb2/tXqYKsifmY88QGGJg8n1B1fg9KqWJQL4GIrNmrRzUWAe1tbMMvffwGmzLqO3kq2UqQcvRDm
SXOdz6GAO6i88oGAv4gUl9WaYCYUxc2oCysUUQ/UKpFC1EWcE/U1xRaSUc3ajR2X9Vnckcom6Yh4
os1asNXAIOzHEshJIr+q8PqEAA77HhqWpRymjZ+PLzoltm6YobWUcC9nRGah4lcVcYX+kSdqIXuA
OovVoGfQj5CtYX5FM+QtxSJg7NQkL/wRO2TNU5gJy9SB1wGM3u8cyW01cpBjpap4AMCKiqj0GjEy
S9ZhnxkoByCWu7nczNDHg3RhMJTBM5By1/rUH/jqQkyfdXwHXN5ycoezeeOsoUpYl9jUu5wYvC7h
Z1NroHb85HGQCPmDfoc03I1RPUoOGh4LuJ3G0309JNtYMzuROyD/Fc+WWt09e1dHVBL8rSb1rWgY
NLny8uYARriPF36iQRZnM3DfhczqsEg7d822WJQPQKFMZKTFbuMTKfuK9YrtyFDdNde3VAoSQJrC
6hBGp917VR2/1BcCwhgNxP9yNMgP8DpmXm2qavLP4SMVRmqroqKhRU7D+gtMBNns/DNDAmA1zmuR
vC1iaQauapO4rLeFn0yCms33l5JuMJ2jwUwoD5NWpREiOWxP2e+QtXEXxzgU/UYU7XnQIn4kOS/a
Bm7h4YyRfF3vfwofsYlDBSc/Y5iMox7cpWTYox6rP/yLIu5OPK/MYT4aZipGIGv0susk60+gS6Q/
8sIDT5Lom+9PYsUdxPzKjvsC3mbrzSVku1oZwpbTIU0BMPrQwGkAbqALGJ9njzo3F+yR1hWs/E3b
IVjCyvroN+mDpomRqXiVkQZjpDeMP68qshildFCPlupcpH5hGC1jAJiA78Mt9+YS1eD6Q0JukCqH
rS3xVGzeAC6V3MigNi7CCA1Fo5Msjvn/nOWz4PNFEN85vWEjRELtxuCIcjKGhcol7ESeCf+3RSSw
XobDXmjsKstlYu2Uoz4SITiaINiyhRMjkrf5fnVHxFqF4ProGISMkw63kiOq65myKVW/Zcz2/0cd
SShlyYarqeA6KggU6uhcjnx36+i7jHkBaex+LMF4bKnAtFPYMCowEpVULi1QYL9yjsVw7GPZClCf
cH8j3hXN4uFgxFotodxcygY8wU/7ytxpA714HNLg6IgTaPNsDl7pLk2i+VeAw5l7xGYSky24dUDb
70Hed6fnf764/oVfW3WQR0FeiVYw1xn9JFlrpRc/QJq9fyWgH3H0/0c2S9j98S4qhZLozk8p1rcI
4WOWXDP1SPITg/eYPp/mE9BwypoIRM+HKazqFgd161ux2sSJR2C9HnQn0QNnxKV+7hX6mTQOlZ0M
9H4Nuo/5jS4rHQ9Yav0XqcTmcNqBSAXw0UD1GxqB4SDM5+ZR8/txUnU6jJ2XhE75vKpJ7Shd+nSi
wSPYaWWErHng9bIBDHKcP7K/mOY9ZO2teYHy60UECiT+IRxZiQHFFDZVcwSYS7ppgqe8x/t5PWW8
tZEb9vQ+aWLghOxcxv4uNursIcoyMv+nPoV6TTjihhdiGvfBVSZYglMe4gakdU6TT2MI24i2TlsA
2oj/cdktwSxEaqH9dRSbIBvbeULsQqtwBAjsFs62InmSL6MCivMSJG3Jj0CbzXIlQFnWcCoV+87c
hlTO+gYLbkO20aIuzHcq8LlU+ZqltQnEF0FhzWz5TmBV7JM8PP/YHKlLYsL0fleX8LkzXa7QWRzX
vE7v0un/FMTAFXTugmSuPP+g2mLQ9z9RaLlrLQ2K+eItDFhDK/xFHJOrD9Ue1P0AkhwUji915Rut
tHzNVta/KFUsuy+Oz9+vvEfkHXkooYmzUbdVtqkz4L2jlDtHwsXQO1iB3xDqklaElx5F0ciAjqol
r3hSx3d5KZ0qU9zYxEjy55BkNKP4f/a6TilVwRFWD0y03MWP63bE4BgUdWdWnBFqyvA1Zzdd/eY8
gr2t3FQO2gxI4ie9iYQGKR7t+7Hv6ypUUAFEfH9A/Qj3+a3b/LQz1v9wUyYEeFlmGafaq8bhv/WF
P/3nN72SGc+RkBTwrA9DDKRtLPdRvhD8db5IBpzE6PKrkrOgsV5mkfThawNr132YCIyn3E3R3yZC
wLuRT9OvVheqiTi1jg+bV6relq7rMJbIZPMmHuudwi2631JwECm9l2K+iGSUxO37cTlcWlE5hcbZ
e7xze1/uohHMfoHZ+GASvpogdaNw1756d9BWVqzHLcUcz/OKX8Td8XpE0eVQb087bsXVBRAMAVUt
je7PYKdPcLksuwg4YaXq29+Mwt5AcuDzBzFgLVNq04atLpe9IBLx968scIIRIvebzjI0W0STZfHA
PswBlczJMmCeuwbvKQRShQRoaWqvN+5cOtWXcRG0YFg2EddYGIIrjLqzAw0RUdUpSQ2V+PrO6hRQ
zh/kds+A8BZcfA5tH32qIIW0qrBaMc6MA4IocHKEF1YRyDCs0nec5YK+WwsLgn2QQQaWtbdstFiD
J2BokMi6c4vbLJF1cBJEWqfuYYXU+zHdOtDKf5adSBhdiJvz4OP0PMQYt6wfnoIoS6gudjhu6y2D
FL568LEhaL6Soy5fc6DAO0lo5Kgsj2IpgcBbXPQ4H0TGxVUyU9OHtPMojy+hQU+ej+HNTs4AMnps
3LbAzl70N5mGjAbcozG0C1RupjBUFmwvTPARq+s8ns5Va4E2pxFza7nVjTG6rueenXvkgmz9gXAN
JXXyMJDnBpz0vQvXnye70+44UZJI/XUe/lssqTjzNl/3a100fJ0yBp+6E1u2T6JCwl1dCwq5xXJZ
5smjb3FCKVSjDza0LOV0hQLz+xpTEMHeyDc6CNIXksyGmPW/T89WtXSmarU6bPQ8RJ83doQNJvaK
OZWsura5Ln6k1djtB65sxIFZ+zLGaCwfUp9eCqr/gRRIfAu88hMBzK1/rJd4x9vTD4DyXaY1uQPI
xpi1wl4s9tzjaT0lIL9IioBLcLgYWpBwdvI3ivvEVOxx86ir0snk4zdIdVxcl2s6k25rvPQS772L
t775iToiLb6atiEtSLGXD3+D9hKeGdgyA+QYtMhgDm1xD3m83SKNxnOhlpMevqysG9pvvlHNP3e1
af/kYXNGy9A756+gRJlWo2r5XOqP9ANoZyQDyQVsg6iKwGxNvTnmU8HjJ4Kt1IAX6oZmcZ1xR9c7
mckwKSEmzwmALoTgtf3rrT7c1nlhdWGlHiqUt3ULYzLnUKx2jgAkdDwxGveBlyZ07movmITKpOg3
k+DkY6ozR94W6GABOioesH5ZgA8K5s00lrvdGrPzqJLskOyxQ4CnkiIu5NglMq76C4Dubf2JdYKe
DInkPkQuJ+VOMY8/v5K8uGAdOItZr9zRoNZjfKP8tWNqG81jNADXIrv7IRSW6UUR29MWTuAWc+0d
wQf/IDsugvTpl6BlfZJoe5R1/0713T1V3kdkRd+l/TDInlve9hDJkwSlmTCstY93FdItGm9j2fwh
RrqrNZC3L/5AwwRAs1OjwP61b8NXS5f/dfnCrlC+6Ds3f03huym+eKUqJrEkHLFWqZNW21dOxFOO
9PSPzBvnOYaKUOBS5YvpnA9nB9+nsiIHAlTCSsboN30S7jlSM19Zy3AFmtsbNx8J2dGwn57ozOWk
lBZfhDpIhvMMuXUh/YRl4/TzcK3ca/oK8DJvSJlNq0jSR4HgYsrNpKGGzzvYvLh0w9n96sAlLonl
vzdISEtJ2oVokRT916nzgfg/TNVOF8jdREFgPX9OmQZu5eDES5STLAzhRzpu+IHCiJjGOo0U4yQw
6A92B7AI5fx8e3+lhTcn2AV4FN759E+1jZMm3IqfDdTaLKsvAbqKKsjgWb4dvSmRqbqCkBURppRz
B5qIBuF0eVZnVW/b8p3MV6UweCCIwoeQook/tig9DTDL7NynDMoAqSAe2CjF+vHOI5+p8reV3Di8
zFJc7SS1VsuM7wL+ZYjnIy5lWfbAsd6k87CucxtNuybS5oLLV9ZcZ4gbgC8CJLgYjDUiS4pItO+o
G8XHgRvRPkqCZwH8W4TIqs6FOeiAyYNpkMhzccDllV/NjthSs7cpuC3DhoJNRgSAn6UmQbvMSZoo
pAF2hr+BK3Ixe/QPTJrTxhJyq35WLHDWWjLRTgpb4AMe8yBXF0hDNcZWAephrywLeIhtFTSx6JZF
AOwMphxDWpwlULR32JMfeaBYUqU8I+9GW7x+RdZIzA1nbZxXN6DOOiNUQ27eDOaYfep5MVKV88UK
W41FGTxKLZNjxk2CkYBS0BuQHunX83vWC78eVpzqDAxVK7m3AXNFWfN4WBojFYOJ1i7M7S6NJk68
0A48WIJ8bv6l7A5r9XLQlTlynIrnTOxlnoJMBA11Ve49POpNluCyXC3FfFGiRwUTwpD62n7vGjEK
6YsfyG8MvJVoZ5c1JewIV+BndaONQcGYkxduNAzNpLPX97zzAZmvgC+kNVF4aOOiFECDast2rBcC
8F2jpWdRv3zQD9Luk9YQpOBFKvCtnlW6CRdWTr+Kw90rwE49I9ESNoNo/TpVwHpKfhtaNeagf/5U
/D/d2hz8XWHjFdGIgneru/Fxns2ldGx8Kx/bK3RCzuZo5/rhZq8vpe/gKeos23T4leMGMbi5D26F
qcQf+Dss3gWYUx3eQ74JGYoai9swNg78naoVrwCu0phiPD3H11S0Gt1C2HWMCxtTbKXCt7JVg9w2
4jgFhUiW+Oste8mG4tdVWZdeMWjeAaVbjoKwG7BpD8snWDkWEQLIL7sKmM1l/6HVt+kw1aIb96J2
EJxuHtMNV0IpPIv5M3Q+zfudb65ct0vq64qYkiCJIfLyKPyjIWgpqIKZg/2STANqPPi+hNZ9/hM1
HR0Iw1rnvGFlXvV65fLZLAkJVZ5Rh381WvUMQ7wJg8rTZw/fWZ1rd2BMbVoxFbuFRwXpyvc3br7t
ZjSr989jqUH67HgZDCeA9/HZrWxjdmwP3lLBv9R7NDVCOlbZ8r98/uecyWYuWg8BrzfOONFYsTlN
ynyENiPy7XLZ5n3ynWEb4NHTPag4WZ9ScoLQ8aSPswFvvB+iX6ttueiUyKseYkPVeVPke4x2j2gn
TxA4nQaY89LUcvX0SFRepYxSNR1S/0kVklTsmhpLmHDXZacw7s1SJVcY9RhDkfq109ZOTyYIUH2A
w2MGKvXKWI5S556OnvR0wJVtueEir0UEwj5Ct6sneQwltj5RSL9tGRS6qxSttxA+t1DgQUW1LR+b
H9TklMBW45uPnLevi+OevQAiLMKcewJtf+wGfjeMyF+/G8HG6VNGiZBebacvFwHcgHFrP71CRYeN
XOY5VllEuP1mYWPPwB5So3Ba3btUZ3XIC9lma8DsqorJeLG4Mx1PQp4RBfNS7HgT/333gwGZeDDr
F2BAkWxYJFZzgyMto+OHm0c7FA5Mz0wd32gv8K+2Ze3qDSFVk5zbjXu7KRQSY571xO8nQdkJrsLm
/TOWMZzmB9frzPhLsc7p91oypCL7JCLtb9XZyOAjY+V7QIkAMa3v4OwQdWnTYqFzoOfnQrC81gmB
MLbYzzNGhHDG0dbJz4vysubeXwu3apA8AUE2XbdM94pnVO/bqD28jmcZDdePS5wyd/K+3wIH6//L
zHZG/vz1vnglS0XNxcYE8HJ14yhXu60dxl5O18+kCtfpTCxvR3UDRl+d7p3ZMQE61lkqGCA1Fge+
DmCmUD+ifPD86bUZwd5gndioyVuKJn1MN8b9TSBWLnhk6+t8QiNl8uR7J+OYsJDqdLkDSoJloR2c
HZ+KXt0i5WsGsERgeG3hvWUNquaqXqDOOivZ2tfAysMdkIB+r1UH1Z/FI7YrsHN402s/H1Ftk2Jj
gFBpH8UBQUI8Pu1rKbwBiHo8s9x9UHNaK0oCahgFbHyfTZM1QR5MvL+cP20IAc/gJykaRVI9I0/e
PJn8Q8k3gRhVB0LCrXDtp0tqGe6bfHUbBrOwCBLTExXnblKFiw536jEHHdGn/l6PWOhC486iFSMT
X7Gw//ldUcu6tucaDBOhATHfoGfsY3fcgtAFbLSaqUpH8IAQuE9dg5E6WzP8pUOjbxq/45LcDnyZ
mNfBTZbZsCetoGFgLffLt52NGRSTWwp4AEr0rJl95UsC0XK4dbWBC8+/068kh48RfjKh93ujLEm8
KxCG3F5QWKaCiySjLrZwNCATHI+E+UsekQkiuNPNfAH0pJUTnmO0I78lvYY31mQPDhiuGfT23BnU
Ud2HGW4K4jbT40he/+djXJpxMe4ZrT8EU58AdQk/PWJmm2Ot6avBj32yFKsUR64w++pO0FPmp/u1
mPoZOF057sLu5NpvjGCdBFPzqsqD/jBH+3uDD9SR9c1PDZHB5wvX4PUw829+isNEFfB7pyf1i8dZ
/XCEVTX3pDy1fiUYoNiPAelBN+CsAhtq3J7cOlaojALKluEoo/beOjgHGc/MxIZ4ZdwRtnpHiLzt
yHy23r/PEqhnJvueZrzlY+mP36QKuf5nB9Vtv3K88kgkNGT89qwLQ71s8UN/PhomSvHWUWgJyg4u
7u1z/a8lsPTNGnmkkJ17m/b4HQDpXGp2o+s5NYnYNX6W3iyH+FoHSvP6XWzYkcD+dlFMRp6jXR3Q
8BSZRxLNgcxqXdt2GyB66Wad6E6pr7hdOT7pbQBezwZXmprfqPgop6jv3GhyyO1LrJ3NG4wCZ6eR
kexrDxdDblJ++oQSEu+gJHhoRC5yphZzFt628VYd4IdZqpKqRI0nse3zsn3BXp5Pl2uJbPcqlBSv
bj3afFHN6A9577W6mMo6oRvLHFrxe6Rg+w9SOh98AILi8tlc7MPB32RG3+0+Pabuw55mnucnnsdZ
f3ONouWgGqXRrcINU5Wv11iqP9N9lBnZ3X+pixMczxzW61leHEeWbCwSDwsdKNL5reIbHYN4jBZP
sUtL5TrtmZwaZo+EusiMovWFVG1gccfjTGlyvf2cTq7+mXM3aYUNZNDIaRh76NsERvmWhPqLQLvE
8xcmbkz7N7SE7xPxuqCDZH3tRD17lCw0gLFXOXUv8+rHhbxBkvbnHhm5cC2fRLh6tChMpUm5qNLf
OQfY9rcbAQllBhoR5ERodkdr9uxTpe9WCeKboVH4EAEQbHOrRSJx4g3TmZebzyZcLmsi/cRXKhgi
r/niZWpTFrrRZjgSnenYii6PEDBf9uMnwl6kraVO9FK1I8kVNOFePExhzLviaWtn9T9VShh1T1JI
G9hXkRMWMg9YCYLXZ7WiFrXA4Vxyu8ZHCLlwNnJOMPRvU0eqxktYcAnwZNUJaZ6hk05L8O9AiLi7
Mdo6MDUPTZTfTgdw1W9bogrQdeUf6bVN8vp3nfSKALXT0+u3gi28rsayYm42mUkHBvpCAi7NRXCx
LiJtQ6oRCCAIN1fSYLP17rlH7F368wLl+PpIFvtrSk5WGnmfacHIqJq1IPtg1hVWXK1NgXwAGAsF
pWRMI1iNpqkB7y9b6LIQg5umGkyk9V3uNF/HqrA/J4zQzuGxAiPosyBtqX/BKd4NkeDD54QOv1zS
gQaq+1NyvdjcOvnBwnn0LXF0XfvmVz4X0YQg999TGfIcV0KEs24/tDY6liiJwVlS3aXdD6F8sYlz
9ixgfVEL+Zb5i0Vv7gQjhW9H5ChHdJ4D4xlX+vDs6dJWmKE0ewo/cVExXlLDcw+hI5zncoEb1ojy
SZV1Ha3HtbL3fMXya1nAP9cHYpEIOcdBTJKozdVzHu0NuKovsKb+Q/XrDqSyPPa0VpO86xmwnhxj
VDWCJgMfku+cHxqx4y9Xtb9G/uxdpNu9NwcLSw1SjchDucSaEnacL9rcbd2yc8R77k3xkOQ7YIbW
FdUhLtDH9v+lc1/QuDJZYnCJhYdW1Fi1MRxWCacf7tF3vYrPgn+DMytYt2aOAviyoQ6KKVl7HA9j
nCF5/slfo098EIgy6JKvVyJTgKJSeb70feIz0IkXfB8OA65AaI8M0pIfSWqloBSfodkQbeg3C44Q
/LPPpw4Z99ECo1kHF8selmkCIO78GcXiCOlOClV1hOy3MBa5/x4nmTwXDOUCqKuRobz8N24oxQJU
yRMRAtMDkyVuZOW5B3iJQU/q2DJah4rCNJuqWX3rx9HX9bXdwItKUoRlGnJ7UBfF0w2uA7do99Ku
RfiCgzC8NX3Xt3nYCP2++fvorko+/eFs87l+k4reSmWjjl9y8W7vCH8eIzaBvCVVv0G64mPApMzT
l9I2bF8/Lejda97Ri/6gdb+NVtTMLVOQCgLjQ+xzSSArZtK/ggnsHCnkmeUKgGG7iiRwE1sQ8zx9
6hY1s4PlyIo4ORr8ktbBDUXuzBsGGAaJJyGif1w9/OjHt6MTthLHc+55gqx+oV2cicUby3Gc7Yc+
BSxHjm633kuLfs9ze83QC1bTBpbUP1pA3rG0LGT4I9Ln4/2ghcPXvBQfoAbNEnN1O+2ZKtUVLvF4
1b7HPMbYqtiKJnRwF4E13bsz7+ejeMhvHG0y/K7bkYCqmCCKIWXwqy/AENcCz+5+TTvaypRiQiAi
1uFncj3d38p4lEVixlQh9yKYR6Bka+lcI4Im4Filmq0SXjv0ieHikP19/QjiZb1NqZuf5ot7Ssyg
HPPL5604Ir4m44t4CeOCuKJHNEZqAu6jWTbo3q4jHt4UzJgUWh/3wjCJfakcBJjolh9VjfDfeJZs
B0OmxL3/J6r05YunsAG2tSCyZT/1ddDHKMOX79EKZhrdOB+zS4GU+GeVjDkek9dThf6AH9U6x8H0
BRKAGfm9ySRbIuoJTMuTvHjZgtAwnJf/WqQdO+DBDvwMYjOIAK94z9p6mp1w7on1BnV+2hITneul
/AnnRgF+JHtt4XXpullsKzTbMqe8cZtzrzTmcDbLTAXszeGC39q8o2hx9BaQkpB73waI/SgfYlAF
0374g6DPk9/Znro5RoV+Lf/BIRDQ7Q1DDWQ1qR+ymyNF7uYrcfcKIKPNHbLpF41XaXpwjEd2ZCyT
/qHiCV2tlqf5Z0CtN8msOayuaYXEGYUwuUiBHjgnyqyup1yY66dHtJYnzNVQM8P9p6vmPSzMAd6N
buaCSBPzBSaIeUC/bppNfLx+XhgN5Gg3z8yTzSPWdw62WqdeSrBbsO9Tk11g+FOnbYVeolB7sd/J
djMP1LPzd/2tVf3117qNMuzqIbvjoToR8sNbmKj/8DMSI7RNM5KO4hQLyeemS+EQMtZU8kxNTjdA
3mtc+3zP7cQ/F1KZipnJs0Fqi5SuOdy1xzy+I9j4mMI4ih0Fakd2fqG9HacOv7BzkL9iSMgVRMZ3
pNb5Xg7coeh9sS+Wvbydw2LJG9SRg8zAdsH60Q9dOI4BI6caYfrdVSb1+Ya/5Zz6ZRQ6SEiAaTpg
rusmYWM6Ic1N+Zgbl0zFJEtRJp012tdPEaW2FuixYqQqGTKJXx2UL22vI78aWyeiv4E1BxuWLNk7
qLkKkJ/amEGFB1isQk3IRkrl9V0rciGMewu2eSuUBI24y4lNzOjWJLHRVRBB1khHB8K6tG8V83hW
/jjxjUXJyXDQXJu2EDLw4SA1TuGLyWedNZYmdc+u/h3SbjyLAj9e2lr0SLMY2DsMdPlhjHUhCj47
4xCv8nE4WBH3B4SzRFiDGw7LQ8r6ugsvbDwLpxvOGOSJPlWbp972h+Y4TMl5t99gqE5Ylp9v7Swu
3cPfmzQqvzd3/USEYMJkvD0u2dtwiNrNfCepQzzZ8uv4OVapiXWu6tOCPY0/mAOia0pu0uR4QC+x
9eTCtyjshJUnEE+oHGnmVDkT9EBahlEdWGzkrillrf6XL+V5uRc2bGb0B22LjCsygFQbMNdVlw44
dmUnJxI5aKenxQmBoOafYJ2iWFyGJiCB6051m9U+p3WxPtEL0dqWtNieOa4Y0mhOI3oKYyKVhuww
AF0dchYltcAgTHJB5k+B5q7TnkZfEMGyo0d+XIZ5/efPSBjCoNGGnyF/tV2FciLYyH9pDjytpUVc
PPFrsePTdRIwVv/X0UkaL44wApFUzvJmWWortupLHS3w4QL6uhW6ciHtgrr/a5AO+Jfd6o5KKiXM
uB3c95Q2Nxxgh2t/nOfRDNx+FlCV+sWQOodpj+Kgtp1WV04aQ10JVacZmQ9kSaMpaNC82/sRojRr
gMtwR0kpqhBwI+KgrAjzcbmXSjERk/khH7Spk5RHFcH02KhrwoiOD8/DYep6b9x53afC/YjmU7ke
Hi4xNKL/ijWvy895PAyv8zd8071FUYmGZvvdxkp8jDr541KhXd5knZpm1OlB/ViDRrzG5hVKXDIL
ERWC/9sP+fUEm86kkwokdTofkbqPFh0wA1pdVP2j8OhRTVDEoqsgK65+f88s+IvreEZIeDJjAk8K
7vP3J8Xwbk0zXi40F/JEDuaIpiAajVSGl5SNNaJXTZ99HFrEx9sfksWtAP7aSdOXEABWqHsMgbNE
ZXyTD1EaxuM6vYEwNBy6+yHvD6zsdKaaJWWaax8BwMbFxmD803i9OZVkYX2rHJR1T8CRCa1cMdvn
pjOwpWK9eGwstHs0MWkwLpd0vZTe8VPvwjgHUmoAcy1gGOtXtUcXfPBTPAP4R/2RLxA/8iGja4fl
9pmgQGbXHletUZV9kMZgzgaCWUAzvPIxXs3xzml7hALQ8DjAzK/58NvkcmxnwsczpQoZ2635hAjJ
bhXQrNvcV+6FN/ICbZMklUT0bf75JOmqUUFBt7nmW3tzF6SfP8UFUnJd1LlM40pEylaPiOLlf3gV
lq6ChF2+dCf/19wvFamhnUuXpzkw1e6ZWUZ70nvChyz5xC0L7EbE+nMRsONFhsnYSlUzjSSpDIof
nPPB5+oGEbYQXg82R0zfK5m5pXV5whrELsmnkyCS6tDiRXuBSAU9aF8t0OYZp8DAbalMMllyG+J8
VuOSa8aGgqdPO9p0bwbq18WVnuXb9YF8SodQ/I6LzObGn7ewF9NW4XinHVZYKO58UCkpKCmEF5Pa
0JK2wxW5ZocDrVbT5ZxXoFRaBpPc9vokwm1FAOWWKEcU0dzUtSoFBQp8OE/WUoNPsKtTn5YsZ+3e
M7Orf7O3VkM4yy+AxEROrW1SPB1/EHr2H1mbuYwSqcxM67hdNIqmcPNzNDynqETlOLFzn2XNKXny
8fQSA/aFjZfwJ6sJz4V05Gf7qdaaqACqvFAYliC2JUAVr5LHwTqNxcVTp6THxMseD/3SgJ3F2aJN
fqdtkmyd007o+wj1NugKbdBgQe79sb0IwHWLRSPAQR561fC4GLDW6io1NpSb8JzjEITzungAIask
bvjsANCZlHVFFQv497975ppwIMxH/nmHtzyjleIsm/tSEsEcNJvvOlTgp1YoHTmJXy68Uk1SaDU/
OalCRO64n/HYivFAYNaoOCdLcsh3LOjn331B5SG0MTZ2y7aABsAy3AW5EVnT2zTnQGMGLWRF7bxU
jXSrde6N/i7FqFpn6NarXL3PpFn37Sa3sKJZk+LiA/iPfIpIy059b1MsSPppCUeSz+aixjh5Pn+v
5yZb9tIQd3+nIeqynY4ubG4Bsx9PYR4dHVuwmOEgFflIooZuH3P45dA5SAttsppGLRE2pLZ6L90K
TW9Gil1R2BLttQuAqFl+rRxmlebQvvfL2pc2lggT/y1UoGVqjrOYYbXOiIM7Klf9hWZbNDBal4zp
6rqWGz8XrllsuJx2KIHWxpII08wfeKhvqIsh91U6BDASt2BZuTZsIZbeEjL9cMSi0/9Uk3gYRzul
gVHMWOng2pzJXdECp9eE+i9SWOME4Q7BAmun2XLuZm70TiNMInKnrb9wefq8qX0YY7036+uRXb65
QZK3mXcifIKSnQTVJWCBkVWT1dLHsMwXn8CCFU7Yb8FUlXD7dkLNGTlE81cTuPNBo+CDZBSN8La4
8cbv2jOfi30MJnryuiJLT1Lf3fpL29Kps1YOhENF43IKCHhyB6YNNOzR+ImRH42G41mIcHECcOop
2MzxP+LbjWnUgOEXWALK9Brm1rsiQyqPG9dlprEEcnhLwpBDpDODVwPT1hBSSj8RDGXLq5LTybgB
8vS431pDadhiFLndo+vO2Dq2eG5eTY5eqlr+aeoUV40NB4MF8mmO1ucO6HUJe5bjwhTIVqnC8zWN
YExChseDBuf+0RufjrHaA5rxgwFoKMHLHW97aXqbpQLP20FvMmksoLQm74RbEFH23PSVLTO0FbjN
cD2PSDQNpTzJuF21iYsK7d+6/B067eakRnIh252gmbAohdk+S+fgJQm96Jgzwq4C1YlfJNMX3whT
saRsdwnraWS13ItRq7qUhFAGhuz2QOCPBpNmUtLSHlgIQvK5VudHfkDBANuYh9cNnR/E+MftekgF
4F0kwXM3mGr444IjdeBjXLutpDBdpvTze8Pqo7zd7neN9jEoWkxo5pitgG6IN60L2Dn8YolotnLq
jhhf3zzaWIZ1jcwWDVAr7wDAcoYcJ6rIpTAgMjpiheJ4a0BojP/XuKjKX6SQgHJl5jhoN+PVIbq6
0sRGg/QVp1wHN0NlPpdmNyCtbuF9XW8Le/c4gVqqZcvGJ7+rgGF0pxQbJzOH40YSRoxJbPPy9D1t
qv/13opYYiqefEUEtlvOmcvzPmjbO2unkoparAKOYa1Sqo0OYKGV8XAIdCNBF30bh01YMdeJ3VxZ
yxmtRo+N/t/YSXBunaz5+FhSgXFmlII1chDE7nECcr6l9cRJKz3Wq/wokks84UzfC82bbtjQqNHX
iLZytwUPCxatJMmZEf6cEdJW9lomQKI0k6lTWOPeG9GaR2Sta+YlwyfnbJbm5RG94jGt0yE9zR/I
VOtVE0oAR1Jmdv9AnoPHT3kAVr7HuM3oONzDEqZ7IXnsjUzifLrQau1CLyfLEc21kFq0uPEwlhBY
7pvWRa44ggWdNSqJmQxYitT3RvV220uEAtHWM2Exvd6heEO4Z+uhKGYlBtyhWVhJD/IE5Zo1luh3
5sg849WvWYt7VoVwFpK9mj4WwkcVCbRi4b35TbuyKSXTpiUrkvBSuNPTI9/o4Mkgj7EW1fs3KR/W
fCC3yr9+zIRFLNlHt6WAhnIy0xs1dBWOWX7Om2emNsoYPz+nifGDw+4N8+/93GeGHSFxw5qggejY
Af3Uu99mjDFbXOwBPnTaPLRMDNXsspu74UuUoKi2Mxi21Ov7HFJw/dg+7+rgfmw8/h1nv507/nR1
duLBJjQC9RBhlvnIXamPf1XOnco9qS0cDaPoDDRw9zIYnP8OAmv13+tbfuXlluRgX9TU6q6YaFj3
P2wqBns99qGPg49Rs0acACbSS44dcICfIJec+V9jPpaNdsdW53eX+UU8/FV65C9RDcL1mkrdh7lP
L7wfqoNIjEAT33oltVPww1UIfIJMCdsTnjSpR8ZepFGi/fVPR3/s4xLM4I/8L4fq4tTpz1vjG517
cGGYS9d3z6mywO4LbW7hf+quwzn3OS3XCh8Q2chQ54JOdfhx7bs8Cy2BU4F2N7foZaU36V3Se07A
5mhhgyL/gLzdOzoGsBAs7yFhe/+G8ykPhPEPLHZOy3Z3iubfAWfQA4OvmkHwgau/IRwE5l9r3tG4
kavX5RX0DUe21d4WuWZExcVR+BmlHzXGfIHenWta0vgXPW+sBCo5ed0l0ymuImTaxE8Mtsoq/1ec
0z/rlnRYzvd9n+vO13U5J/daQjThYo5PB1mp3m9fthDk+YGPwwBE+MIaBE8uok3LeX2f+39oIPmj
s5L2MbtlaMvidxsNec9Xc0+UyXGYUurCvHRlLF7ak6tOiRhrNv3lWoLUrdNfJFWJcTWDKC2GwHYD
VXLiFacld/XC/V12nOA1v0WtwKX/X7RkMUqXXCX1i8OXWJFtOrDNLSeiEZ3HnFnStBtJTVmzBFX1
oOec0CzoMs5ypT5HqR3rrtenQ8hnzxLlwM1vMjR8chEjil+EiAYQNOe49sbFXMnga+pPJIF61xNg
17c63jGjhpYqQu0lR9Pznio2RCnpC2ZslzZWx0vG/DCBpeQPiVhQP1LAGmxTr+22oWLs+eqXldrE
629zkL6Zn4xKsF5nwsbF1i7cd8Q3lhLZt+iGtEPGYPgq3YkK9GGKtwSUdywxGEwndu8PQwk7ZSyX
QZ4660irktRRopy79KQ5l77k/IE8wI4QBuYHGDicZhmkScd35iXZc5wwnR0UBwT6vqGcS5+tW0Mp
6WC4s8Uq94CpWV3PZ7ubwYnIW4LM/F39PBPkjgw7vWYsvGL4eM0yuXPUAZGvskeE9viIe0V6xg58
SnLIC2a/ZUsMtv8123XOMWhy9G4JV/ii76k6cCZSZImH4kc6SDH6sXn7ZprYbZ+L9nV7rMkcGJpK
S2ZmUD+OuKiA8IR7pKHHKyp1mUwX4y4GPTEfyl/u/HQySQsLUurGdqo3kxdEJn0ftXfp7wKJ/CpN
v3d2sBFwrDdjIS8aZOvwkTxUQms12yA0U24RjwOPDxNh2/320x9bPcn49pkxGvESwWhV7OvYbvuf
31wCYM8xTwlAv5Z9ViwDlmtnMOX8qp3pRBLu/4Rwfa1i/fU/+BqSOCIHqmpVb/3CoUY7KS+LSR8b
JJDpSd8KewP6nqUdDT+iMWnM1nvltDRkJ+bzr3Pu1q59KI/miuUi7zJOL7YUirby47gMpcIw7On3
zSzKZ+Gx5VjKtm20+JHFsokJP0hACt8hVKY3w2dofwC/CRd2PJ8FaRd57MQOgo+uPhBP0a6jxvwf
YauGoh1Tcn1POboyB3YYRGbWjQ32DN8F4tk8n+nNygbN6R2hzmi9rmIFuJBWeADOtOqdyPBQhx0h
533PzWtamEpI8g5GvTqsB6UVq9NExYi1nKpkMfDv0qa8wi3wXGJ1PwWaRlZHDR1Gv5zseU8frB1j
C/X724xw0yfcH6vGmv5H//UF1hk89ltcj9HMBvOeb7rAvFgkhRjSZ2c0muAs63M8MXXE2qtlF+j3
5rIUhV68DF5YdEo7YS39+ROJ0jbd+NeRy8SCFMKhttFszLqWP1ypMXegZ41G6RrQQZlNVduRWXUQ
V+ZQ5Fanp+SHhtPX/jw7eNakLZQWM5f4SuHnOcDHMs/WgowdRzfxvzix4GxrVm1s34ScNmZUNJhW
ZhG54LQKk7JDfyJcB/JVX/+KV24+50UOkI6m2b2uz4V0mtKrWgLeZ2AyRf0G6iWLP1uQcrPrBFqa
duQR88zVDtxTNuEbr+IHXZGekprGRAJDbpZyVpksid+5izAC/QQ3PZvBYjuXN2hLNkQKVkf/3esu
zARrdqyN70pkIVRoTyXsHI2ZNaVLhVLjGtPBXuRADs4pqc0x2I/hcq6rDuW6GlRtM9Cu8Balfz94
uH7V8GaJ5nNbeFUxOr16rpiB+XNlwkfhhrxqyHv6vbEmvuaRAxlmXoshgSLH3Jbkv1CLZTHAReXj
Gx/oNNoyPismPvHXAdkuakg44rJiUS5zbjIoTu3urX0oBnAW6QfgM0c5Ce9TJuUXaeFcuOxycvbE
KZMLwer+gGBw8SLo8NfL1tAbmNZU6AnA2HXzOxHlr6g1B4dBvTIGaWmWMza2pS5S2muk+d077OIX
cwfjFZgi9ikGC4rYVEF2x3h2ONw9glUOUgUakkamYDWAhagrcjSUCTowqpxVzBqKnNdXQh4xI9OZ
YKSXrLDl0zVIzaHgJDHjfbwk4jLX6MQMmENd1yVNCOnZckQ59rI9p+/4x8f9nAmu1y8WYw8lPwgb
tAg9tKOkmYrQkT/0VphxCjXgc1xPJyo6b5FCOHazuOiViqXA7/gEqt92BOSn3zCN/Lpnmo+aMGJW
T7Yu1L+eLnRD152pK3lOqoqT2EE+qDvU3KaZ7XvzSBL4132NJvzP6r8k/sudQcU3/4WBau8cw/jK
gWwHTRLqKq/u7cdOiQxWMlx+OSedm+dFSmRZwbCjWKbAON5cxD4L7WnXe7vQqJhwgU0/0Z17Oss8
iTYDg8YLQJGj0gYntTeoINHL71j1HNHwwl8B2FfoOtDCgotO907StW0qcCbLLoEg6a1Qx9jTOmUu
cgnoTAKSzQUJM3oDIOsbPV1IE3CZjLxSh26PRCxllZQf7l2FLyBcVVFhm7NvOBhpu2Jf5upejRcu
/vLdvewAiCPASbTY+lrHZDsAyz7BgafWD5pVhy7zDuxYneH9+1sKH9qcpmeLaVJ0nwxWYB/zJG+E
gwXmP3Ea6q9dihDxdq14Z0/5Est+AgmzFh6Ly+g+rtqxVDvxlzDuko4LW88RMWkjojDcogU7GIE9
zZJ3Jax+9F3RJQVU5rHbTGu2f3oI2kbsKrN7rKS55/O8gJlXcLxbiGgoHlxF30VOLquA/0+qEYFG
WmKjAGjCIEQ7BzJ/mxlOqdb6Fo8RgxjEkU/qQLfQ7bgaAe7MZ/cRk7eaG0n98ff32qbRe7S+UAvR
hIZTAV6MrMeR9kfE83+hHn5QXaO3bRfn4ZDcUDvTTXCESvISw5OuKq8UV9zoqAjUKVhuHz/ZUMgB
X5UkSHDJ8oinOcG10mGWs4KSzzkMCWl5S8oGa3xHjJv7IO0Ab8iyJLYJxqCOK/7BH/aBCk3JXd+4
uTpXDrvnkSOKE+GrXQEp0UQkjG1fhN2SJtiRwzF5PiO7BbRAafGVTQfHTAlOomTjrDuf1exOkp60
Fs3b5DCYMwU3Pzgfyc2pMpb1vPrZFtZB8kX+Lxkpd5U11Tj0LnA1o9JOcY7fyc8iwZ6QZ73+4sCL
0+XbFxA5KVjqNNKhguZVeTTX/79zcLIJbisLCVSFMyJdOVABcz7+xriVXsTsl0csIx6nVHaxDIyG
hhE38sSlNgtYLV2GX06JWum6/FFIjQNf+9XQ9Pbl/DNKVMsuP8L+sufHnXZF8UKppRmcnzZr2kET
reUdubM6Lxqq56PjNNS2pXsCBdy/AnQSdruEnlPcxQCrAhdTa/RU106AwezlUzDvTzua+cAGNb7o
ZfQNUMDH1sRfIzs9xdxyqTlH5yNLWqnXt12DlhawvBfPHFKsw/wmsRtRZPgbXISYdVWKJD/JBtko
9ZyPAbVqE6/ZRk0uL+aADsyFvhz9BMSnsLIxCPJA/+wrF5eSgT7IXzwGQV0x3XNDm2xeSB2bg5/f
imSdJWLGfnl1feMA0w2O8wGlwTE3BDntZDT3ZILO9t9e4XGqrYYzWeXOVIw9C1DkiPsr6zzoA5Iq
qSRtzlF8pD+qw92lK2uuv1FSjBfBNLGhd4iT4x/s+2TSOLwaR3d8j4/fVTYO0y/D+xcBPVblockG
KUfanvpLIMV1kb6eKAeJ9naPp/nq6gVoDRuXmFXgP3AoV6tAbj7nmUTGq3Jy2rhY2Ziq/U2bbBX0
UO6PjCGsuvczjn79xq5e+9aX7DRs7gOi443g2loFpz6s0txwDMvwQtZ6ZYbev/YWDjUng/GxIigb
E6c9FEFvrKe1O23lyKkgXSaNdXGQnp8MHVDe6Kpkbv+dMzE0pqJUNQOK6De5MMEzi9lR5Lz85NWD
Te3l+I+h5n0zk7KLqmTFRRR6KeBZrl3EBm4RO3cPKh2z0SHthdoauuvpfQf2Xj3S3cmy8HR8QKqC
2jEa2NSOy6XWNHXUKFnpgQW1NH3R/bVlZVt8sCRBGCXVJBDMLgPm4F2UrOtuWrMpWCbqJyxxbdnF
exqsJFvwuhtns1GshTGU1mTytUoJJjI4InE+RyJMrcaB3orVAQ8ModrfXvL7FoetiSUtqofbQnGA
OQQFFraJhXni+3LevmpeV6t3DdowTCtZK+zvzqvwwkXgoYR5fVW7GVYHX9n8AI5Gi2KTNn4oseaE
bx+Qu2fdrj/1pEAfP09IJXDT/ZzQvuadGCO10WCA3sE+d1Qgs/1pY8Sk/Yi63reQBS65Hde5mOK1
tAB6VQzSNvbntO2tqmpJ4/sauTl/nm//StLFtpxQZMJrdaP9WOz2BsasGJVSH2VsuEzU+KW9fNsg
PNO/1Tce+rkiWtwn/GTIVwvNM//F9nfdbhWjWVE6NrMbAYX8QMjsRlHIQYAyfAJ1HEQd1o3KXjx7
QOCjon0t3y83SHM2HBEb16Pb5zkG2DKc0fpL3XR72aQAnX8dppsk/Z7FJjVeO2Mfio0CHqc0ifkz
Kf3nKU2REUP13/L0jl/Msr5q6nJ8zuGqBDH4zOyeEzu4c/wzDR6kVQW0ssO/6NSR+AZxVv/GmeEo
wUTKaWIaXdHHDncHJ6XDj9S9G94TrnPEdJQeUKA2wIvpKLFfZ4WxnzlcGnK3860wTpshVWe/2964
4tQKfnX/xCsjClnK27F2dFibKXRWNb0JwhZwWf/5nSwzi6LOTit7I6qwBOpE6Fvx72FLGarTKI24
QDNUqSLopNJzPiPcGgb7QLoxJg+Dqp/AxICKW22xg2rWSAriNPQ4YQ6VFXng3OLMwOF6lI9YApG6
8X0TkrUvRBjhLiv1xsFthLsrDjzsViEo6icbs38LF9wlc93AeB2ys1lvpWKm07ogLWjDnOMoCX/1
uniu6O7KlfNeWdSej/gSBXx7YY12Sy0zL9viB818Wm6Fa8YRoPq4TKxxQXMx5B7+0O4jJCyXxofH
RNgjKxuXXHQFZajCt3GyxuyHmzVchwboZW3tg4ZtqC0QYv6v6WJMzjCLwmAZe8I9ZUWOdU8zhrpo
FHroQZkwABqyecMcneh4Plw0Cxu5HgQltJPEBQqUGpoCpMZSw5CVD6CSECZC3vH4V3TuFAkZRyxz
/oNlBB041bYx246zDYay913twv+MvweAsdsXr55CDU/77GLoZKZhB/w/GSPFK4Q2MxQfEOv/xJKu
ngzYr3MnifUH+Pn5eltRSHbDLhEE+ZH+PHonoCciQb+ocLe5zldDEhvZxgACcA5m/ipZk5/ufatC
RyfNOBK0cgvFppXv1hsVyfL9xvHS+f06UArBNkaQy0TKvtWVYZzaWafh5N7lgK8bhLXW360+OEDy
8AtsaKhyrO18owamZ3HorMUTrijhLuh57s9KnGhxv4CKpogYXtsxMnKtbl2tZ+vBRv0BbAGkJilx
TEpTUs7f10g6wLxT+g/jlUCgjztzWRn/oV+qH0DArW3C9o/BUjNPz88N4GvqKnnQ55e3ZbskvTwP
HT2aQotVDlejE/STtE+cLmX2vwOyO98lxjiMs9CXvPzCuFe00fmppcRwrdjqL89QupbbNIzKibu9
5l9vUzvsVeWDnnnKz9DBf8xI7k4O1ILN9dyE903lWM8PmBLij/4GE8PjD+65f7/h7lVlvpHuYYUw
t+HEhu3M7Pu5y8D+eLoj3+Uk5ytpwt+TmAeN7Mm5bXo4jdmyOSHZmW8nYCQ2VUSpfnhxOcsMjFj4
75BUqqs3C7pqWa5sStKlXurrCUI5SAtDbHXm9TjFF5WvhiDdYJyLfrQIWs5NM8IKiDYZzku8gU4x
72ZJ1gbRlr8NRjvZuNCN2MRySKat3ZZDcYkQdjVtmut9Xlqxisxi3OEVFc+ERHZ+AwbbftpUQi7S
d69xK2MIP7IvYkjlJzfKdiMiNXDPcvABnRwR6QXRDlnb4QlePfiADAVlIK7UXi8SyombHuCBrnVm
lmanAmCNEscEjp5dedK/jO1yQ4zuNfiFdJrUklNnRjDthnvu+EFxfaJtNAzabhuLWwxEwpx5QnQW
taCXRdRBrQIpFKICH0pR/lkqynCDf10MAeQ1o3DmXiEbpYPGkgWEMrJhfi1fhNggozWawuWohDF5
LMxnjG/U894tgtI8BiIQtn2A97FR7hE+osxchPvzlrNkJbq9wbNeegM8Pbzb8+cB0/vsddp5im+C
AXJpNmKUelKcHKYp6SGzJ1lciq8UMullJiyr9E8DKVS2nIjegqC5i5HiBoq4n73gjwApAUg3MmuO
DwHc3oOP1t9lYh/3uFQOB2NwSm1UR7aAjOMQ7ZV1ym36tFCWft/UGfOnrZUxDdS0aURoxmzG2K61
DSyMI7I9X0IAEsV2M2dXfVuT6YJ9Go7q1+OwLqqtNVxOu33vqJU4/9FkVprUa2c62DA/OdzCIC0H
L0xCgMKfonc5bp/e607RG9sDuVyPyrC6ZMfq2xuoG6p0lDc3mx4c5tIkRBBIFHZYpXA1U58QdIZG
U9bTxyhqjvsg3tJ1VJsa3dS4UteBedqjFxAXw6ChrbxJCV4T1D4uPzz9iRyPR3lb9fME/WNBvz6s
Ev1fzpi+01sqGIOc5MZ/7yJamZ/jL13YCZews9fWUoJElCJbRjYrz+akiJyji8OSY9cY5xbBRYFZ
F9VcPxCzzBlUEWyGfnHEnEgjz1r2oF4+2ZGpiqolGH0U50di5IwH18RFNnoxN/i/2FpFRJmdzvSh
+PWUTes+D68r3xQYGzcSLGaMMnlVMwTIHovgzCbwiXPtJBy5agoLJHXrQ2uipWCLpPAl2kEXyMRH
MHfuOXMHe9q16fANXvsIJXMhz6vJT9jmtUwk0+b/43p8nBUFhME831BoE2GGM6KCkzWZsX4atNOT
D7GNUVLxKxcUJoQl/fDiIV0/pXfNjNt6dAJdwHOAV4x+zrhb6T67hZymn0jXt50aiXjEqlS++kaM
fzTt24AgJtze8eeLj5R93wNbmIjPqG6kn3BAtWrTOfbr16KRh4aUwI3QE3aQV3lSQslm0euOlJk5
Z6+iSXSaJGTESEbh9HTlyxK/djr03CoYB/IN70LS105pG8GWNP2scJ+ERh0BbxPzkR7ohrjkorUS
w5rCuMrCpriWSnxsiGLZI4R5Lo8U9RqU6w0QR0/Mdx0IXiESbexSjDV8MfglLMPT3ZEJ5wlRn8+f
MbLJeP7d4dPVQZ48hQhN5wkh0yRggF16324v1bqCpwgslz5REHRCOGxzOivzEM/wSsVo0OoMz2Pp
1pHNp6PfzaRJA/4vZAoCkXThA3bE61yhfMZuT3Nme9+CabQ4wQMJmSSohO6eiOoe1PxakMRBPQnz
IFKHnJ7zs7eBqHxCVmWtamtYxOkD+laIz0VaZmT3IW1uc1kqA7oVGt6C5FTSCDVQl0y+jyeX/KIC
n7PTM0sC//FkkVTlB0PVB+6JN5GHSa1KVqi/Y5dNkuJBELdfKasIfpEiRKJ5yAK3UahPYXoBQzv8
1gR+ukGDjr0QudeMV7gJxO1ZW8OwWPYPH+yhgbw2p8Bk/g7BfYrejL+4Dn2kqXRjDLew7hBkPUKN
EKnr1sbZoQXjRGOp8dhCDNaFSwExV7oSaQyl1boA7LxoCDg8SlA/KtzDAWa1CebXwY7RvIUPgY91
tIfD5ScMboa2QLBsMRMdMUE99N1GVZ4mRa9CBtxjgDKeZFPNMKcDsG0zShDfq2Pwb2yEC7mm4z4V
cckTiH6V+pq48+utluKSzkDa9zoMc4xalsOdqxoOyJbHQgJqgY59zzKJ1grWKRRnN8fbBc/BD8P2
ZRcvOXgFWwVxmyUPfaHYyYA72NUUmMNwuUENOkvruDvs/HgKpwWAzo08VELay5eI5hSHJsoU6+qC
oAOhmiGLH2N5P8TcxEKOEplyLoSjrw/31wYJx1+QSa+we20UOk8JSXUKwNqCnk5G+n0Hbk+lhy3N
RzS45hTvNyRDpa0tud1tXTktsdxBF+8tDGs7I36IIctp7VcqV0d3sp6Tofsg5pwSw7Xj9Ahlpzwt
93SDmoiqeG6cs/AZ62NTrDPrgk8ppooJrDA366+R/7QU2/UyFs8ou2sONO8F/xwII3wdAJUmCL1q
yg6XPecMTlB5LAR8gxnNWswprM+BpyZ+HcxJ8R84o1Ymz7z5IkHQ17jBATAiGGwKQ4vieBtAPCZk
UMr03sDPOZe+M2ZepClZLjzRr0E1fVKvf7poyF1UuokYVV384zMHf+DbejJ4qoXhfI8u55w6LI37
TrhR+7EMIO6BKbRIDTsZoC8lEYhK3KPRghSNbOf5CAetvNDQIxnnfgN0Tf9zlfytOUveB9TaTPfw
+DzPbSTisCtammFS/Au45/GLZbvDxPIf/taaJtQg5PwiAVEssaHNPwCV3JnOduzzeOgAqWDYdqzy
/HIUYRlY6MP3S6SzErODq5UQqZCGHwboRG3KhFNIpqrjYWp3Ag3XirIDEK3pZZCIZ0IG+FxfrnYE
LAQK31M8+LZH+WcHw5rnem55bOL/InPThFJXcD6Ws0cnQi7a5eR+6RwslkPsu34HzdRebF/aTFWg
qOe6aKQl5dOHjZeYe6pdzYxjqiOrpF/JUnSxexibJ5LCMzSkpvNZ6pb3hfdHYDAe0wReftoevzuf
7hZ8s2nAuni+1+zA+N7FHEUEhvKV+W8uO24aLRp5/cKbAzXxUDCXHYOWbnza4zpEgmxMT0z51+Yl
k/1sDeE2NAyFOBo8ckszN/VtA2iIW4PPDQuYvl6vbyAJYw++TGnqaQTjqm8fHOh1HfO9LC0pakvp
l/jY6Nr7Knk0iIa2rY925Go86IyIFfls8pOVCyv7zvFkpLq1GzHgXGR6BbIMVPYyhySpZbGUGzAQ
ke4ikURQKJlS93QHQ8xOBtGX6hG2t0PE1XkfoM31z0387MJXeup6izFCLw8YzeddivDpxU18v+2K
/E24GlNGvhZbb8fnvzUXwYdGejOUOtvdIhkUXhDWMePbTNdSUEb3VAeKsVlV9CzJnXMgV4fd20lK
axwZphmnVD2edibrrEs8ZU0mPHqvaARoW4zF/x5irf49O20jgP1oQFGh1XyqqtpqBYOtm0LEqhm0
NFWUhHN2Jnbxx+PTcLlkrh82yRQ3YID9a9j+L0Sg+9mO9i+NlMqLRXLsVP937c+VrCwxOlhB2Uom
59pY4hKq0q0lTens9hECw3LhxZQfgFCuOviht/s/Inw+nqQmfH36Pcmj118kxoBpmpfsETM3A9CZ
4VRpnG+wA5W2oZ5WcxTXARUo1qAqD4R0gTv6ffuLNGCJTki+Yws0WBywhYyN/kHgV9HBOsKF6TFq
zGZzFV/GfE76jupOnQvuNvvWn1T2OAOCEulASvVWP6TpdlEAtCiDvqBX990/FRa9JrcVF4G8II1w
GgkfpPaU8KTrww9yHFqL72oR1DKDA6DMv4In1kxmXMj3P4zCOC1Z33LPweykiNFykJ/8bo46am/3
WVdauAzLb76/mOXKnpm5FjW2Koph3yxQ0qlIUSIqaDicjoLCJ+M6XSKb82hS45tXJ0brek7hizwk
VyFxIN0tV8hJYdGTrz4tQ5OU7aoBwuAk4x3GWGNZ4UcP5axd2VqzGHC598QStvKNAJsbhgDGFwwh
UZuw6YbeX2qVV7WyTvZfh0R5oC6oa10fQhV7spW44+KqUcn2GgwUke56jK8FOqLGC3+8HCUaN0OF
B/eoWM+LVQC6+EgqDGK2UY+Lfzuvjjk+nL3MA+CkMt0/pcUpEyiPmteIShr79bYrDe72SRoInA46
JIwVAMyjRDZneG+k/91V6CBQm/4lhC/gNZSdtBI20TkgP9z21uouwvqyVFl+aGW/oSmLajHBZSnG
C/LQn5CH+jhA4aAKrCkymoNvRVMXtetpRs4cvqJWLQTTJrdnl7O1ifyKZyZIwhcb8GJ9Dx+nazI0
Pqg5bXaoWd0QDNLuCYql/uyejPocLz/hvZlfQAynUlwREj2qMJNhP1yGRRHGnrAmYhihqOL2dSsl
lfkrBokMor2qHqDqwzaOybpm/S2acquQBDw44lbn4/aV0WUSRYaJXZy1gPHozt+9uX9ofjLiuh3L
IQymKnt+qh5uREZvfO3os8zDasfRxwqbgMzjppS9UMMw3q1uWSNltQoq+RIevOCpjjNlym950U8D
zRB+X3VCugodpgEwdubpxli9n6356t56iorSgh2uRCU5i6cl3WsAWmekgWa2eGaKpYrIZh02FzSO
mDBuFh1II1Z9WrM9puqRZ3nWPjo5S0dLMonbnl7B6CKeXZQkJc3bBsIbRoMdfxkepkWZKfV28gd+
M2zWzfaDjemS4qJ0a084+hc22T8MMuxXJKzhTY2b8/6Ruk7Yd8Of54FlDTz8SCrhRdIWDmqvJWbd
1WF6YF7A0oqASyfjGcI9nRBgex9v/t+i28937p4ixj6a8d8JYuSHcSD80Ie5pjn5QP9gVEa/j5/h
SS9e81/I5EAcPoImOo7gHLaAGe5nbQeS1aEg65mBVdw+4qk/JDXVA1ROWRRUcKqH/9850SvXeYxs
0NUhQpXrTcHsRATVJkR6b2PnMKWANaD0VVr+Nx2diCH56gX4h9o40owetwTd2uFj43JO6ECo94kw
wMovJXKwXfnqV1Pv/nIFc57z0X0Eq1NF5L3yi+wu5M3wKnAUQnIx/5Rd+UrKqWEiKfQcb6hQABfe
OntGthz+zO2ArEvg6p1WnbOBBmxxobOGSAyYPeI/cBbRQgYe1jTba+klvJuEPz64fgiOSgtI18VY
6mF0DdquTsAumTulz00ZryFAepANiOZPnGWoq66BJSGqtna3QiOftw9cGlXNEpfxvSRm+yS6TGYi
MdIWBn5E8jB2+LBMVw+vZ/d2wmMHAYs0SJ/eeToMUyvTh6qlW4cd2Pn45Nk+5luyuGJpL/cVrJUS
jQR2tkpzMvW41wenpz2Uk0TIgwjOQBqYB5TGy3SVPIdO6mgL/MmgIetMSxP0Ny0NejwGZnnJikMN
/e/pXBKfxG/BiO9U5bAHxU7DbGarqIy6UNwIrYgJXQQo9zDBIU0wkN+vE5ofpEUd6cJXcaqSHizu
L1FNv1NMsJ/OXz1lUXisVq/UvSNDy+xmkBBVKl72TUmfJIEclmJAcM4Th2nbHWDvoZbFpBUy33t/
JUCeO/kLpPDgzXYAcGxZQWNulJuKJPQt6DVXYXzWe9JNdTI9Qupr7NCe64Adq2PxOC779lQegkPq
Hb5ZsDBnyuOZS3XFL4lr/b8G7vTisfEm4h5XnZejLXbkgaptab0H2eUpT4RtABZjU0u7LThfnKSk
OA2ZBLKoFFDSIV4aYch87i/1KWrL4M8Mr97AiWcueaTRCOqLIFUZbsDnP9ULPzl37ksYQC09lQOh
7DS4jLd2zeetySp1655QOPIRm1099QufLRSgllcrZHQPuQeYGVk+FyoGoQZ4FxHr3PZ1UL8BScCF
IHLwPX3Xuuq7Ohzpmx3/hG5cyz36FgdDe3QUtLXuTfTvTii6w6s+ZgkyPAbZxZHkv3RZeVonDUDW
l/AeCOgiYVtQ3rBrq0TykllWSE16GGbdbnfpRtIl+X6Vcl/3C2mhZtCfVNN9V+rUWBsOG4LbWNxK
7AUdVtM5AewxfB1CIt7febNyPofqTi3bJxQzaWZZ+mZRHAH9KlKSDxf792J0PUdb15tcy2LJZ3rH
74aCFKBN56Ta77NwbWISprFu0YSJDrKGk+XDgBH6xVtVHRLP/HagHZcA3/2hRIw5YrjjhDX+1GkN
GvW3HhGYuro9pZM0AnvDfhAOB9OkkhGBk+oCy2OZtRRBJOFprtsso4JjCxzE4+Jafo9pjpJJNl/2
XnWd43x7sldJXA0RJvWUGY+iG1CFLGLP2UdXNhGKj4xIeQSUOmDVDRgeXCyO1q92nBIFi9DXWOf0
J5ayL1VxE99Xjl/Svl5PZGNGZ7PknM4cQWhYHkLBTMok1J6YsGtLEXTKbz/LPTy2pifeq+k49kNo
Qt3WL28JbQGcECpTyFH5IZhxWH/KaVihNru68r9rQC5DbWaR9PR9b0wxDxc8yPTZlSihTAnaG6vw
5b6l4I7N1S+9XAiwV2Xg+225GLKwGHUqVmiVbZOzEpVAgHHNQdZ3nIzjnVKjdUSpX8xIG45WyuV6
qIp2yhg59eWYWHipekymgnBuIwyKnGsMayc34dBJyx6cPzO+I/XAAgTfJVY3ejCCVQFhkQD7mTEv
vioz72+AlE3oAUZG5z5FSR3mHC5L5/18y8KhHOnAUFeRe/B6eOZtUzqVaCDPiEkS1R3gVoHSc1g0
K2M+WQVqTb6/JGc7P4Ylfaboj0F9aybe9QsAgmRoJGabUw3yeV1Yut7cwStf631w/bcmEtlaDbyO
ycB37GoRWtAPTHp+77WXnsC6cSARENgnzaxB/ml+s84xckOsvMT+fPlSvpIseEimtt2NqxxjZV7Z
6p5ObWwPZF5y7GoiKtX9O7GKHRmx62vhsHt0zG2kLn70vNK+jQUi6WMeAsSImcP8YJU/Pe5e+ZNM
gee1KZsAXY0KlGNag09YoARCawLl+q4dKMwjavN/TvmO05EETdDFaSPSk8St6QWDoqAaTMdXqJgl
M5dpMumChUF6dzZuG7a2qV2teEzoTpH8c3PrQrujkpa31Yo4CArSMyDzx6hbY0zrpsr9DTP/DIf4
cRM4YSdWQMLf9vAxgKyuovoYYEUu11Q7Lnb5wjHa3BROPihKxzcnW+8fOe1pexMEcOnyocOiDyjA
zQUVC+Yibi29Nnvy9yirHFmTctJ9ypqJkA/iARXuDrPuWHVa/A0b0X/VnTbJFFxumg4appFhF2jb
wyNNnQ3s3y0J7kD+9g8PfwX0TWYZScTlStra/8oCokOzcPympml9NHdd76e5lJmS2CTIjCizLmKd
TLkaPK8+MOsOCCK3CXie/PzYvUKJencCV154s5w8iT6sHzhji/86N0NbAviJGNENLcqilOsTh8vk
y97We8g1AxaGEiH5nyMMIYu5tUooj7fyRLjYpat8kHNrTks+HZPk0HsxsYu1N/1fFsz+PrqJEofx
izVdn5iIMNj1ciTV9W3RiOH/b6bDk7spupvFTb+RmxZPtkT7DVMwVoOAQE0P1EuJtjZzhIYjzTYF
klB3zeyX+4S9yY7MceTtr+ewhzGoV+m0zM+0eF1LQoHs5Cec0XqEb8H/SoFyEI5RXSXrlydG6L+r
FP2kLsTaGCQC7SQK47rrMHphr2MgQxay7R5gmsmpkoHEvaP+NVPG3IxqMoFpRlfqqQ3LtfJROIXy
rO7vUUAw/WbKwPVhtlN7CYvizjQ+yxMAqNSsjadXOWGzisDA37V1sVl5mZcaf5btQR44HF7Bud+w
ySxjx2xnmpoqbWfoHhMLttD5l8Ug1iu6meHjzXOhIg8VXcHXp7iKMNxTaw74ZdpTSGWM0ROVc3I2
GD0yiINoFWgCWMf8zilm3bRA/wmV8mu1ugc3EMn+wjtAg8topllvRJrvGFT2HrSQdWllD3pfd2aD
vdF9WJoaW7reM4dZ68WGiwcXNiAvFiAOSpnNYBLJxqBNVWXPrwXSWjTTyJTGSH8OlwKjTtPaXuK/
A3yxT0Z35EZhS16l8uvtINdejFfWC5PrsTeiJIP/TuiRkxqVo/YD3jgO33HnVyIqPLrGZkmTqYK3
IoK1cb4lATU5FVxMG+SMbrt6oxxwOT+zvn1Hvsw/OPYo43bii/zTjdB0qTq0uu03Ic749EJReEzQ
Fr7vq62oM2q02SQ8rnKgvdhaXMWtL20awoNTslr3+3ne3HheK18lipNnP8CLhehhOiDRXWEFN4OD
gQZCTxUMgyYLUBEOwFyqOvgTVCGi/gjyfDIhBN3KsJWMjRemC+k3GzcTbUJG/T1pc8atHxBQTfVG
ZFOwOQnZVsbDwQaEe36lR1aryPga4NElEdtr8EwOiyWGkTynGz3DYbYLmaop2jmTUQQwOvIGEJpM
jX4miUMhfxjxPCfW9YK3/4eE9X5KefEq7aVFezWBRdEbSfKDB6Z7I2GrjoZNEROCHJwXBHLYBDV4
uwZOJQKpZmmNCH2sTSdlx5smDslTxvk9/4MucKihWGmTXAMHdm4G0odEQIZdmhlLh/xv/2vaLiS5
y79i3M++2BMUUh6+kF8xnWpd6ufiDJ21GtZvPeVMM55zox0YEsWwXKtHg+tHyfj89b2RlHy14Xjg
oljQfEsjtXo7RoCGClfBHrwQPhnUcNll4Wwr3KZtdi+ETlegj68L6XwOUkkRg0Nh7TOR1kee5F++
PAoh++om92mpjRFXwpkBJA8jz4jWWAUaa/wLZf0exGXAEGx5n/teAoH67NVBQVDzGGdVHR7ZMGTW
vrTe14y6lu/p4jACdhnx/PNaB/9Vi7bP/UnI/yXfef90o5mrLrp5ZhnFGXXUI9htp7hHrYKaP7kU
mhjwYeI6DmWMtuj8N9Z6+JbbR76LGpe/igVFsiUmaNcuyifMyt5FfJnxnoeXaistjMujBBmyvOcK
7v2wPysWKLYPactHYiTBE1k72genkuA6Ney7Hk/RJQ5NN0gCNQZMRs8BfdUJhfrOpyKbbwFVSkol
iB1nPo81kpudOptEWUM1Np5RCD8Ud6yr+j8Bimk+w1ayes4cHP6bdIsLDYw+TjfzFjIUM3c/kq8X
K5nkEUFaOG/JaMAYVoMnzKHKnlKcvJg3RdnoTqbKhEYzYeeWAwxkY3c9yFg+pLB8v+ZKKZzYW3w7
qZRivwA8H5BtYscqQ0Z/Bu+QZopye0EFP256H99bRXkgfT/oOikHfDyk6SOp/IItPPvKPLf+NdmZ
5vnlgwc1/d6XsQ8s7XweAtFx1xrYKVQiZ6qfKbl64CAxjb7w3pzNQzN7Bmr+iwy22TwCuNPcBReh
gBnKvKnCc1Ad7dk1mYGzniyaa//c0tkom5o3sc+L5oNzURrdtt2y61CS9Lh5WvjD5kdGCFDgFLUn
iGDcbikDFwn+pLIIqDcYcS4k5glG7HxrbXzUYDD2prypBduLd0o0UORYgpJpRjNWCMIfNZUtpRRP
PiJNNIz2IVxNQwHnvpNDL/mtSysTk3vqfKn2UJ9M0U82uIahra/7ZNaOj40tK6t7waMZpf4b9UEZ
Jcr7S8SGyF5OKsFctpHU76kNDmrscvxBelbpl2cHBMshPobtQBDtSa+TcE5HC9NIcgAtMUd9c2UW
qX9tD9FptA+skSDiOnoHeSZGHC7tZpxFSzpVP4IXpwZFKT0xD06snnr4Xc1EWD7o8v6VThe4tfvz
dG3ZvCEXlLGZQa+2xfUzmU+y24HTutSQU79R/UaZXIJaKNNHLyFlNUukEGqVwcDIf2Ew5AoiQIrs
46QAYmUgxO4G9e043YWdED8wIYV+5foFIrM3kYuNntVYpok5pPSvuNmMNa8ko2A64hA02Bb/xk1f
6z+cqI3HWBBZBhUGcVM+ozHtT1MWdI5c8hGVYGOuggSSrHGJ12ans8Za89i858y12kiOI7RQpn8P
4o0RE+akfr4R521H/QLfgMgmfPIzMJb//1ix3WuCx7ksBxCmJb+opqIJAMs4g8rUQ7a+M7WdWSCW
xYwFZmvtnmoW7PePvNxIpQGECXWvGsaeqWohe0YvDwn9xaUNa81f1QSs9LtrpSFbZAqFDduvhDG+
btjIgOVJB1WvvVTBkt4gJxEYit0CVRzJ48QYa6vH1alfhlpdJ6GeLRhMrHLkOdwEddh9PLgbIYmo
2LTpvorXKqlFiBpvY+IKA9sF/4uZEgWjb9IGLMHMaMd+qd+qXZgjYFNmGUntTsVlwgKgR4HMVkcM
ydspyPc+4BFzNoRfHFGEFgBHGQLbjluaIiduRTjZvcU/YV8YLlM4B2NYssF/n3bkH8kqlGEhTQRV
AALmmr11hLp/+5tsbs7cW5JWXHPdURP5c0S5lAEat0ZXgHe5aY/Zzo/6BYOFZs9DgoBzlLDYR+/+
in+Cp11EqZV5ZS4qvYfzuTYZ4iF3z6loxG/ECwKRCqLP2agT7I0boHd7KvTlArdZFewhKA+Y8EfO
eIzRTtWFZeRpm0MiuiUdWhy2jttFOgmzNrA4LLMzlj9EELVHki9nh6r/rEN3lYxocM4vhNRuzRq1
fVBq1Y9gSCiVbUiP1+pR9yJUQQs2mgJHPecF++PowV0xMaoez8FP39D1f0o6Qyynx7c4h5jqUgnI
3eszsCzFGCtkeaZdGd8w/3NgR91srfXOrs6jCgnr9FybxXutW6MFnznKlBV29iQEFelvHBJjEpOU
7tBCgMaFDlxV5NKY7T0KOZ7hxOXeKH69H+5GQTEk1sxONpeANmoMosxZ0jsHQmQ1LlD4bvVVJS9j
Th66VG8w7bxfYO6qYjp1fJ00882VGSDUKjs/5UId9NmOqBjRRDIKrTOrV4Ry77T4Y4L7AGmFHy4k
dybgM17Xio5zzQxo07aWkQtu7gSDfZgID/bVjXMu4mWJTnRfVWsToDMm5AXhbb6EcDm22gCEA9YT
YcR/v+KoNOHc+6zSlmr2stLWPmnCAH9Ypljb1qKu7/gNWDvWAICwgCQ7ft+0e70H9mg6AOofxRBC
Nunc//cguCN5USOM9yipGr6DDA1ttcugp65wJt70HSyOx7KoKCR703+0z9sINPRw5oZyXOr/fTXK
7PqNydUe16KhNFDhY7uBOHqu2QfG+AzUMFYPn7Af/9r0YHx51ca2PQVVYDSkO/LDHXVhB4e63V0c
76b+6CVKz9Yq1nzUJ6RA+XnnH1qAHG+vO38bDpFG01cq89gGVRfxNd9NfNRn5ixgi2TtT6rW/tOZ
ztQNS/xJJVZe8xbUFan/kpo5HSVXk5gGLy/eU5cFJnOZZIyXt7LnLE2aze3wJYNtDmXY7FjGcE+/
E9dICleWmfI14gEwk+umlCqmozWu2J5Tn9ds3JCq8HCpmAqOeCI8l2DyuzJKU5F9ZWGHkEaYSY/r
HwgfGlP+eD6CqVNm3/6wHEO0vJXZsneZU5N2jpqxqWaIwaw+WBk50APdnoIbzH0DLaliRMvDgsJd
Z2yor/PCQR6u6YDOvvKkJvii2JbexpyrB86RyxXFg4gZbTaqhie/efpIGY0Omw4BWIaSvOvjDBZd
EQ2aTPFm+aM0blX/1l7gxxzpeIUuBulXqRWUXW5kk5dg3rxcz72Eto1EdMKBCif72rYY2yt88as9
jcxbLySqGj7wsqlG3dYkyAI6a8GaLlaKo19iSCN9Cgb1+34fX9W0pE5P/HGwoVMGaNdXNhzeG3i9
TSXrig/f+SZaDGoL29JkYhTRDbeSe6c5V8g0A/Ik8H1TsYJYlRn/jWjrWYUERqHyfgeWwSbGntZG
yXKceFH/SeHmSeoyE26c/qheNG8BdqOYxaQOMlip63UjoQg65OGYuaTPC9Znej+CKw6KTrxcCvdx
dl7xxz2RrNo3h+pstjW9WD/xMkvLsllI1dxdSF00GRtrumAR/HhmpKBSS0g/h9P2It62jJ/Pp32+
1N04+g20OM5c/YJwnFzKOhJGvmVaM/tjvAwJHTJ47H1sxFEj9jAVy7+Lle3IeUwlI3NQiR3xAA1n
yqHSzPtoCjthncc2RSUSBhRzaTbb6xzurzOgrFRrakU2SXH6IenMn75D6EQWlglSlEhbC1Zuw6f/
YwjzA8+zIksqT4VGI3b0QV/hqXRsRGyFsQtNR77z75GGpcve8rHGTwKVrFZkKme3+06YHFO4aIRL
36AjiLeyCv39mT9o/W/q8XWJYtnshWq1V84om/cLtzp+vVX4dK68/5yWxbApdhor4AT15+q7S27Q
puLfcShbRNmMKG2PgQWfAOTOO4JVqJdmAxEelEgXQAfzYs750ZycRcEa9MMa157CeYsA6Hpg8lVd
LpzBM1VDlFi+IUAwUc6R4zn709Xd3B+wgX0VCTDnHk3McH56/V9MM4ieETFBknJ/ES3Kb1zGFFNi
uMtBjjtdXOxSuL3Vb36jdX+W5kHF8mqx8PE4eu/nmoQATSdY1zDT8eG7+KO0TxQZKMgYYemVvfvv
4yEWI2rhwxJHN1+G7W9MaaAwq9hyCfjGnx0K/7x30S8M9rJifrp/L5LopNACjMZu0bOH7p7ct7B3
7pI5ivLfE/xVZ8Ihi1wlRJD5a1EM0g9JQcLxO+/nGM5K8wiVuosMV1JtgpZTLAazXSNvUkkUG4uV
3VhOzHGy8noVdJ99l/fMqFhplqLntDxuBSfQuSM6Pt7zd4VJZYI82QWPxj/hprbIETFM5PfPDmRx
JLKNunuHxQO0nK+2yzzrOqPhZOytrRlwDv0V6TyWmXOIgMDO66SsmWUBJMue1MF/aABe6BwxThuc
S64f/K97hAYJ6FOm//N3W9NGpzbcJQheA8mjp7dbjOiv8fWTVUccqagTtAqXQy31xL0U9w4RqUTx
oEnUCbDfNA0TynGAI3FA0jJ6Zb4Of5PzuNhWf41k++6B9QA8BtHqJ0x+FDs4xLTbJqq8vSNUG99T
Qk65c+EjrEv4XDz3yDPMw5DPOZGlcaGvkreuKxgJVEe/5j9MWLzUJbPsQyj3anIw4ZQQQmoOiYFU
z1pE0gp6iue17kN0SXUkGP3ZcvCLRJ2lZrG+F246ta3SD/xFctsO/jwnN9o5ykWdsKpppIi8yeI0
O0CPk8UAO2UUOi+ksDle4DuWIHHG8C1TYBB1+HZkJZYEtNyw6gaE4cxYkQFG9ftCPBl06iKNGFf5
/Ea0xVwxRzdJq5UiJ358N2VYp3m8t/QWKwGR8eXW+K2nK497QWYOhg9xv5U/mLfAGidS2VN66erB
BvSbgEftKLdL+TIye0mPP7kR0/2Aj7LBm2cMqWOS3Yz2jCR2daSYmRYEmB4jcQg3cFFvcozHZ/r/
L561ZkOjAOK11+AmpEAH7YvEfvUU9NcsLn45Lpi2CR+TWKdLsXOOU+83ZhlXVe8JUCCefpu4cLnj
RT8dC2tmd/jqfM1l06v474JZV1THrvTcZzsInGaza7kywxbV8DLOHzLjJLMZKhsDMHSob/5LgZ8r
9S22sSVk4uy1evUgyIhM4KEFPgJrfWsfMF56jyzyl0mTDCNG8Ib0UQmOT6KWPryvtqyTui3MeMLj
p/snDoLXlYV4ZC9zRPoCgH1tzo3QD8jHCZPZBDkUC8Q+cAtWCHFLmbEO9szc80yBVFAquC6U0rVr
w8RzTKiXqWFkPNqnTLjkMMR1inpLOL98dPRtvm9zQHMEZD945fjrmbnKiR070jobW3w6JyLzStLy
f2N/8nsC7d3KoC5xWtdJu44EhBeR5Z5K7dthQYdTWCHf/Ce2Cm0asMi1G4wwVtIrY7L75j7c2HxL
zs45yJyXmhbgum9rVuzlmU9WD3n3ScCH5tpHHNPq9NPHXeys2amqOpPSfFFrRmg9oHnWuitwdP0H
NbEJkzgGSc8u5QN+xsVMGZNEtVknGdbFT+8nGOvIqg5tjpUBwaGgqjUo5GfGtg+qfBQ3x9FbrFR3
dhfa39GqaKElR/wjuOT6cHFq5dSZWJyyYJ7yoU7Go9DtukIPJepXrAcxwjNiddwJ7P82iCsYITyB
Uh0D8v4K0hZzjwUPZkpuWNF2ganzNK2hwJxPYF5KlI08A/YVO0mVSvNDTHMLUpPjrVzsrMMx5v7m
KSOxndqVMxaAhEaGeXDBzEAvI80MjWXWmxipRKtaSq477CztoNziJ7VkBsoafMqDiM2Wn30ZfVf+
Cx+fOVSanMy5uwZDEMRGnUgHw1sNMCWes++E+IknfcOFzh4I4m1+i+ZUELZD3m83XY1jAUcwzvow
SuehOzH6dFhx+opU9Ph5uYWvwr5362eH8TcWW3+ovmraHcN5avN3gka3BTemFV6QQDFuLpFwPKRd
xXRbp7pXr15o6mHuTNGITOIRWtHt28n4+ihWCw8jQ6+sIgztumLtQaxsGQMw6485w9qC6Hbtifkj
KNglcOESKYPpjfFvT28+zNZn1Dmr8G3uYpyeZzpggQnPzt5o2fvYTywA2kpaqr34pdfIlQEsRRwn
avRSKJ2OkS1Xk5SmzvNiDM8m5ASLBbkz6f5O09f0uaIPSHPgS8RZRwuu6GX0nOwtKWTnNbTDHjDw
ej4O6V7uUjiLJG0On06WlVohS5+v4lhQQrcxuKTM1jyc9TKjLnrpCKq9olCA099GFLIoPLzmu5jd
K+kzq1ldBIc2IjsAP5kqJ6loFoL4e2dfubtH82Pn8U1FaYCzk7P+OspuW1uVOwvnD/ZoDiRV+gsv
tMZLwUqPNxvkEqcHtZlJoiykCK0kphFyjI3sHD7Cu3hS/mm/p8er00mrpE2eQo3hhH8FqKKKWE5D
qZYZqL+fO+DxvhxzNRTFiyiVayUWdNO3ZJP1wSanW/aj75DnMzMZNdH3BxY601LctmMHgwOAv4iA
XwBQpbLq8toKTw2xUwsOteTu85hmVVgSo6QWRvkYbrptDzmkYlE9bJpiaGYORT/4RFLZrQJ3sbBz
szOJcO0BrMfn38rjJuqDfqK/yp57bQDEdB0X+Z6e6UbW+h1Qj0fbpf2x9SerLfw3SYBfnD55W6nq
XD2yt0qbFyl6ZWe2d2/MV5ArIUuwUTGv1wVB9m0co8GHkJQRowzhb0AjoRwYUSjX4alA1TlEzaqj
4ybEvQKuMen4xWoxlIB3z1MmGYQpaVDgiw/pWjmElaEniYbNq+BUTJT0e2U40rwVkvxrPXtkqxrp
aJ2NrTj/oCW8L1oaOMhueKRR7IiClZm0dpuvhCntSNFaoZpICZo2edKvgBoZkKHYwzGwwbh0kGxH
vIcw5yIYPmkOI0GNYDDYR5p7USpTsp87vcCqfE3COsvkcnAtsVUlEB0udyP4cOt233F0MuqAR1HN
+7whohbwDzLzEwCsYZPn4ACk6zPKMKeSGHAXHcnzmO2R0zPo15uddltE8D91JIzRyCrNyvuXQ16U
7zQgc5MvLUB84ub5pVpMO3t3saIHtRaunlD8kXC6TWbgLDY+DyMP7+UDIjmsyWkpl3Q4RYCIyjRo
o0y162OjgKI41G9ZdWj4V7DmQvn+V8kD5Ej44yORqNxSRlwD756uwVPiXoSH4Ygdj2ee1bQ1Q7Sl
NiO1fbC+aCm7Q7VwvHSJ07sV+/6b6ypfemCauctxBW6HdXZxXQdZJVmd2dQEOXtYispRuJN+LigH
sz5LkD/0kPogZ+f3exnyIVR60p8QPRFYQzphc6kjfQlFFT6F1CHmSUt/qHxFffwwY5Ptxk0qGAzV
BwVlQu+1XJnjA6NItOP6kFzw3kEU2CQiws3DaRA/mKvn3iVqK/h2kWfRTT5J3F6ERk/IDv0Dtzqn
jFJEzpsSC8CoHG5gr5wR+y11816kSwNKsaEHzvNZOJOr0OeOBrtJQLkd5ELjEoZU+OMPWW5PB2Q2
r2Giiz9x2RsxQcmRIsBYxtV2eycOPo+y55Ie6YbYVQ27pubfWDGRuAlpsg6a53kSyzzXnizBmzBY
OOVw6DvgLyBXLz6EQonWeVd39EK8I3b7sGvQryy9DjD3EOBAF1cYhQA6NSZAsApIhVKV1x8DUgPr
O4XIbsaNgQV2Swc0KD+tDhU+aXAV2S8aPJGrChL7cktf0pnso2a6htHcOJdmmHCEwsNxuI3kDvrG
JibTuRV1vHuJLF8Jsp85dtZJvtb9j6ZgV9xU9WEq8bUPWHHhCO2C9Ix3vtl8jh506ak/ntiPiRlC
wFGaXyDu6bVSwXtnpZJoE7AjufmLZkG/QFaImY1bTwZRU1wDSR/AhqKCKv5KrwlYfQmCdfbYl6AE
zGj1DY2YdVAI7cjPWfd0u62VvRybvaOjLNYxfejQ9LyeUL3bHOUQSAeu0yuUJiZVwRz8Q1gHHHc4
Y09EvSZ5Po0Fw/a+BvQ2cVX24+sjLkpeal0N126vD9GS/jqaDV1DpyumzRxEaPYk2ndoRgQpDXMx
dFOt7CB9JrKYTiRcwUMJDwRQeDSF2a8odyd0N0+elBVpQcQeMLbYlED1bUX1kv7OmFapG26iIoKq
KoAduxO1chJjDr/tiZYQGLf8uyXSKgowl2t8V7aXVJQ8+X2CEwgCIhWvxmfOviH6/pel3S/gjDcK
A1bHkL76hf4Q3vSCRhtglQJsD7bOENZsPptPsfmTbQJybS4AVfPKZkAmaOJMCwfyTlptj58s1wZF
5Zm29EGHyCiOhzI+Mp5/iL4uCwyRfM6z8zsY9OZyQsi2C7q5wO2tpbvJtyl+zq9sqDr10RHfw4M4
1I7puO59IsWFMBaAAdbmS949p6kPThX9d4Gn1gTMIq2Vq6W3Jbe3icpXsXB1v70VumqCPrtSuM1L
c/BqvQurWRrTBTTQu0C4y5kX/cjEoPJovmdU2zV3Gmb4DBA3SkV+yg5Lkmxb89VE74eh3bnj+pgG
lPFFTRU8CDwMrYzGaJXwA3Ys+HxJLsuA7hLbzw/RK3/Z4SC3UbmEQW3+SN+8ZyEB4LCpPoQRl7Pn
b+waiykWwYDGzXFIqGQDp1im9CX1se0w33I+9VxF05N8azGR2xHZopZz4IsxjR+nrK5oycpiC1v4
nlYGbThmCFjRRf3lik28FBDQt6wSa/jl260d0JphySxmKXAhyl1I/Y6EV/R0wlyO5sSNBXRyB7C9
IgQ9LhhUB3Pv8zsG8y6ImXyco1RERLwAyocREWy4j7R/f1/vcXuxxJlCEB0uPzpsWrnHSJHPIH/8
bRZpu2IM5pMkJAU0HUUkhrfkUavrjhlV7B2vy+2I1XF/DNW5sg9RbRJo01lvbUMIrKEd7VGpaRND
47L5RSranYguunwjtfNc3SrHL/z+DkLHkAptkkX6YcRDKcS9Rah1L3SwXFCzdiWGirYD6DJh51Qg
334WJYHYSkjb8DUk7A5tsoa5Evbc6sDMS4dGbSKu+eRZ/mFo6LnHCMnvsgCrBh1wFnVnY6a2fpIF
eVAaHkEBg+svfxFaBfOD/MHHaI09ty9+Sy37HZwqkvG4iMGKPXTjQOyAx0hGi/1yZKL4Thlsjsyu
j8GzmUYkQMDQEX+ClMTcW0qC2+3C2JQDqOgCUaxvrrfhHVh8vouc2y9QsgtnJFXmoE0woZ7+igJE
vug4qFbwpPjST1xIjwwNonBproF5qDoupav+FxD5jNhYYQbiN4cgjFXzZCXLeOFalVY6//GoNWG+
OZJ7h+xdqwCK9s9j7Yl6mH71aFAA98idFTOOLuM/ifUObyrxsEyZfX8hd3Oh/czIo8iS8g4QQHNJ
pUEvP4ZdiD3UbNACuxdCgnA1h9zFlQv/UDH6ZN+1oTMSqpWbYXn8gJVz8I4DDaTCatho77rUKfGA
/VUEWxA+3ZXi/TmWYugNMGcHnFFAeukYqjoe+c/8Ep+dk9gePbxOYlHcPGh+VSXiKeFttNxs0LGR
Tyjna9rF0W6JUuCoG1O/S9DPOWIspEi2C9hSjTS4IijxoetRqtM0xQgBIODckRT59yXz2qWrO9qu
cVkn39Pcxcm1J9KdbRUF2yD+HOD9RTdB4CnQTjYgsW/0/Y1m559YtF5NdLoxmLF5wdIhXXY4v8Ov
jeRl5sU5cCB2nRXdaXOC2uVnv8P+Nchh4WF+OImvI3iD2BMf1RpXdSAaM4YKPkdXrBKxLozqJFsj
u7fTs0bx1GFlqpkcH01v1NSo7nahk9e12I0kGJfZVyS/10aUYUMklwLwrVe11+QwyAIHP61E//oP
zGgKmt9AHS9Uppz5McwX+5bBi2+KD9rQcuVpt19wGTwKFLb+IV1Ylm5Fmp/KtC5XjzpOJ2xsLUX4
27pWu7fjVvaFsM4K23lHdLgau2F/Z56liNNGEsioQvR7BSMQDfKI6OSRmcW35bIOEfpRdFcjG6Pu
fnZy8ofnkVH7LTu2qTTttbTFvDTNwkI+DQ0n5dNPYxx4c2A02I/9f814RnYTSyy1nEKjFDHkGmhD
tEmPz3LJ+e2vRz70jgP3oSjjvHh+9nRlGMkvgR3ayy8OL1jJVifJT5xRRRQ3cdo6gy0p4RKkqrY3
mYQ6qiu2kul3X/W9aG3eg2v3QhY7+C6Zkq+sUwe1ddExkRp6pKmciYRwzCdGlXsj87HMly5Y+6M7
a/whhl6hED5cGAO0A1NLRR3oeb4X7YPl99c4FIjXctixPUw3W6CYH7wBu/l4v2XlSULcquWkhmrU
5w+437+n8oL+cJYvKsEKb/iGX3jPmEffBE0Ca6smjneNmoDRNF3md/AoT3C16xinZodIRVFWvDd5
+iQYfRyGWj0ILgSJSh7QPpUvfJD9Gbw8ZvBLk3z9Q96dYAupNafYaj3+Fjvn/wV5hfnCgg22CCrp
+snc7bc4e7JVla5IqIvmlzdFews4BxrQu2JqKad1QZket31DDhYaLZ8uBmgJ/zq5lcFB7u3chwBx
AsxFyDd0EEUAfIo3jLekk8n+wyrqhac+VKDxL1n20QJtQcGIs+0JBd3zwtb8itoCt0wT5IZo6drP
yRILNjveGs3DijTIdAAJUiGRX2nJRzV3p1AENnb4tRxhR/0cd0IfCPMCaj24YH+Iconec9Qd9tSS
9tc8OHKZ//BsfgrIllQA5eVtcMJT8NYAbEPcz+MuF7J4GWNHGv+TJPQkp6pfO3GEdMtWmt4hMcBs
NCftnkOrXyBAC6E4BL7pCJQu4WIVkMTcEMXil/G+sEKFnUrrCgcNu1+TcO9k4h1jrqCdt/8dvLbs
993sc4jdY+8WZj1LZqFQSOu9EdhfGFXTdnvrMFwhXQ4lbO+lB5OYiTcGohkDf3E0ndm5LbpX6VfX
MzQabo2etlJKaQ0+5g3vP66aWzgFuvrwa3ICffjlo1+JumTcDdHsJA+SOaWgw3pGnbXCNbYOZnts
C45jpLK19p3EfXRMF+f+JaotvlAJo2avL7NENOoASWnb+uK9fhOe8Rv2EdEu7HZYAoreA09SItnm
yrso9W9PNKf4qDUZf72YZRsWAijT7zDQD81Ayz1kvBY0on0HXN8CwxwQg/e5AOiDphfQhQVepWeW
13CKwB+nUuZZx18pNknAIXTbngXmIwid/USOlV1ngZJALRKX8XzHLWAKKZ6MGUe+bn/4P+myyhde
CadHDQchEPUcbFldvnWcoICunMlctE2uliyKed/Hzu05p/h18ev6DGEQTT2cx1nZGF+C4p/3u1+F
fGKK1yOSVMga4F7AXV+BTsoNbtqpyWWSbp/bV42/xO9LAnWmMK+uUfQpAmAzV81eu5aVW0hkyW8j
okWz030omlbom02ZA6Ok2S5/Aj1fFw9s3Nu2YjThhafrrFMMkbpR9SUuxRRxt93z119+ecTY7XN2
JSx/htYVaIbd1ctG67NlbFahXHs8WK2qz3ZCCJWpm1uuP4eJ8+JJTM7+lfYWa4CgjE8qRM5B7Laf
LcMelB7+HgM486XZnzAqRRFaxTzuMaHDu6mPYvp45oOg/effyxRiiSTbWz6W6eRRuYMbXBfMv3Ma
VdDjnoYCAB0T0alJ2CzUPAh6Z1ZU0BV+H3DmsKTW3fM8tBDj6g1yygD76k62lvBklgT04Mf+LFGq
SWGl8RZ0M+Bz/UAFqwWUdb8kUsUiH+YA0//+CQQ2tkUyMP76N6Spct6+i9ddhFzmjqSiiihIWhaS
tqfuPS6NaQVolmlKWfeAC73PZ+sFm0jEEPuT7Mc5/PB91LD7PQmQ4EcE9CBNtwokBBk1OCPWfHs8
FdzBzce4S/UxhA2XNpJCf5ZDHCwvlmyf2ElWvUP2HPP0/rdl6qXtaNQRifqTP5inYYfOF8A/Ia1f
Gaix+snYqQz6lJYfq8o52NJQC/uGuG7hwRpgUvvRmQwn2D8Px/Xt8OHPa5jqpJPuCIV41JHKo80S
NZ3/lC+NLA1m2tfPx4G4hva7Gm9u58ePy8SZ9YpF+N9QLLU3hk/OaMp95EOob0jy5o2rOCqOXNKO
UFdv5Cj5xlZypmXhJ2s9dw48wojmcqV/xSWxs6CJXCx/jLXuSs06xlo24PE1TDoI8bnT24eTD2CO
O3651OAbgerOc1kmt6zctXxkUzi/Z0jyyAVwDR8R2GLXYWQXM/1LBFy7QKWOEQtRpHCnDiENoy8j
pARsYZa85YqhNsN+kx5bGU6anAN+7rL/qECuBwuB48Tf7tpB3adFjU9K1epjfngiPnSUZ49Mega/
JiCAjKXdcwthztWYj1Pb213L+rGRvIROUD+BDYD9rSB2ghU8fIgKhA7hH83K2X3fF4ujkEf33fVG
UUdHXUCXq97Vlg+xSjckMnhk4PAeaijyZLzffMifJNVawyzORF+d+FNpmcQnGQXTyZAksQ4nfSfR
/vMYf+U4C6+1CDFNUks+OdA8a3K9pNtyS1IYmZmASQs6QWyCLYSNF7beBgdQ9AKZwZknvtkHcCGL
OzrrbT5485djE3Yp+H7JLYnKp3Ky0h3LKs7N6V5aKqUoGjuLb1pNcluBY4+BTt2wgDNN7MNJIuKj
ahb27JcpqExZETaNR2BlDLgNKJZcpROh9oDXtD0zJE79UdLymevYaQ88GcsaqQf002ukkw4qgD59
bhUhVOqntTcHXdIPbt2eUI8rM7GtXSam3RzfvB4CXDJyXMi5sbnhrZeI6TDm0zebcHLDM40HLAR5
om/txwxgMNN60aVv2w9x/xrjHwMn7meFmIfpmgiCvBYYKMwERW2p/ZtJFX62Ri6SwhekocFvJ/LU
cYt4FSkeMZfGzY7dqn4LU2xFJbSZvIOqxhXHk9cgitDUqo5OInuiqATdKl/WwzSxqwC4AFuRiH+5
PWRVKSm5xBreo/fCVdu/Dcm7CBPib+0mBiIXD8heqqlR8dgKSZK3RsYF5ktUy938vitcSSVhRIgW
oefY4BMcJoEkgKfOCAwSF/+hy+2EkokMrnrQOruvcI/gk/xtTUeeX3Q6PxQUt78HV49CQwoIq0nA
P8W+B/QWfWWKj9oxcOjCne2A4T6yCcwJBSnUxYbPL8cih7OkFBxNN/pUysM13K029KN62hET+6sc
jYHNp3y5AaP8MJhlqom6N6j47AvEli9V2h8KFm7/qaMP2ytrbH03FPVubjUjXVNpi2FR5XufA6Pm
pRCxFZrjWMCB6M0dQn6uGor7UeTCPNSWn/fFSgJ5gRve4teyIUkiYw4B1JQCR6Y3H028jrmoS1Ev
I0xZUphcu1Nh/TGm1QbkOjPwokVLoTEzkdF6phTVTnUQ8QT1/AFYcaupN8Q0usPTGgb7TtD/97Ap
YzYF/cQGHXnf6yXgArIbH2XFC9q6GmYApfBMUy4aUNc9Zp6hwLn+HOYo7XKTRqIaC6Mv/LVE6Obi
FZdu0Zq7WOa1D0xGufDs1jwaqS/XK91J1DtZFSK8uOsUVD6gdKkVBEd3AL0pQ4LJO2a2It8TShPf
Nrt7HoWzGTtZW61QccffVOE6heGGiZnQ1aJ9bZHfHBaD7C0G+4H/BGEwxvmL8TskdnQ4WQmII3mU
6wgVZtZFNKYFlSPagvc5rpnzDOye9mnTOS9ebhdmz5FZQYcSd19Gnu73pD2qTqh/as4wIukE2bGB
YBREfrvaE8RsKhju1Lx4TGkdqFTfO4IEoxQzfvbm3iULGmbaEyzHO2ZUKfMp+Amjs7qCIiWGVues
lnx6KY4tfv9dZ8HeCSWMZ65tij44RyqoYjzROaoTG8cbqy7gR0DA1MdJF+kyjZm+Yxxs2jqxyBAx
A+E+AYypjfmd94spEoBQsLu0nUBMi9DEN17UX6nL6ybzLOkudwVBEGbEiAbmdQH5R6YyKUqKLQOW
5aYLDnSP+YGxQNHov/RMvnala0yrBYLctIpXZyCuvop3aflTlHkatSpUIXIsz8WqDvzZc/loamXt
AGZIhpzi4CK7yybXPfYZL2KNaHLfLSKbC1gJaCpcybjLatzJAbPh0F9Fvq7BRy8uuGLj0lIODkzS
ALfnFXjPeJ5aG5KdASNWZ9RqRM6BpiYzAB9gj643vvxA7eIyB5rPXbRBUg6T/tQSghcoIIxROYKA
FvLcrK9qY5wCW/pwX9w7h9sVn/q56UO2pa3dX0g1gFrZTNuTD3t1UzB5qnobYJgBvDQmgHik3mi4
ulYGSsxrUguWQRlMFhGwucxJZwVtovEf4SLeR6Tmg9T/l75Bq+75s5m9jSIDDCVh5+VAdqC3D95o
D61bDnq1lcxoW/DEhIIVYf+t0zjiMi6IEyiHhoIOu7xdn+3pDMvMP3UgwLJqAPGDrrbsNH7XMNxs
D8BsUysWzbRNAxWIjijHSsj96yxlrBg9g6vJMmRlUcmIS767/LV48LCnxzKJMEmiDHWiTRHCQ6q5
XUvLc396ygZ0TrRiNe6O1zu9ieRyo+mh471IgkNZovGZI3k9z+DVO8UJrnA8IJIob+8SfJRmMPWO
QpRbMPnva7oLpLbyh1t/Kst78H18HNSosJY37EXWRFRicEdepohyjMvsTfymy/AdA+Pxh9ucGR9P
A9NVl4zfrjY0MUeMth997kvlQP83zHJ16wM1+MY1PCg5oFjXbZUXdiOlWbmf/CHS0YRYsc4QNMjk
GLqZYKvL2J9iYVE6aA/Nxi4RxRJ944xFZrCz5II2wWjjuWdl6eAXoT8vQbL8tI4/NY6ZGn/rNCFc
DsshY3Pl6i6kmb6psSH0EfAGkjIWf5u6tsJgxAddLFtidrGUtbV2vylV/aQ+jfJJrT9XKafAEC4T
BhI+sEKTMWc8lTqIhFbUQpdzutRuVHccmTkknlwcXgOIkIR9H8HJXTYtXnfEIUWjuiCSqhKVRN64
uvfV7eY68VB9AHAvuryrb9hAQYMdKvHRZpVFstQa6OPP6LMALTXlA+MMVKqoqH2jtzCV/gv/LAGc
bscIZBiYKNF9YqFLtLMrTxP78wcAcSkGS+KexDzBvoiGao3RGMvRiBThr2A9imXRd0vOcZgGWPUN
0bOCmxg8lgYYRtLKzxNyIcBZyXzoNPajPGFNwurxlCiN4tHgDUy8EtWSSSCA0TjGKsiRZytRzkMM
+ojduc3DyfGB0I09x54tt32FBDGE6kilIKAKQQz+gu67SmyoprvUfSOoLmeIQkwNlTS+LEwFlUr9
GYz3t2LusbiXhVCfHGqVkNxRFNVcjRZNjbN7eZKxsfFZnxBnMv0Xj2fZu9CB/gmgVZhLItX/eaH3
a8KjB30HHrqVjhYJ29U+TiNH/zy70Wm+tjR0Txfhg4vnqbBI563NkVnU/0Aeb3LIGuW8l59dzWwb
T4DG4jH/9CFwla0cRjs7qeCVpGL6kuFeJR34mAf8eyXeJsUbzeaAh3Zc+knfykB2nLZjr5BTgTlb
83qPVIggnA1Zj3VkyxiWLfGJal1gi3+D3+UOuRJnE6PiS4/GbzK4bRjL8xrg1pkHnykKy1IerTXZ
XkH0vFacoVECAkkC1VM9JCUJP9L5GcMIM0MlEd7boTH/lJDZ8tqL7405qPnQdqIczsr9zL5g1sYd
zfgURSNYFET7/lzivBLK30sRN8xjYVFKSRaNXWMQiJmS4PaRvClGqHca+7k9yUcqaRH3PFh8CbxK
DzN2OME597pof2WHD603HpwFwDKRXwSLh/IpgzN/xqI3ceRsWwoRa0VEXKtT2OBjq0oSM9XnZQLm
H6zzFkroObAHeilaZmRNHhfe1DYHJwPPWXsKbdsIk5li7CZQOTZ7Pf0jWQLZ3MYWY4eX4LTOnGJL
If5KZhaiI/zpZKQOTvoFeGJpgO3eNDuI81++MUnE/C8cgdx9XiPpreVxZmw+FaJGaaUaAbSR7NNz
rHeZ2xC3Rh5jG18Wd+y0AIgTkm4tbH73jmH1NbBw0nEAhZ3obrpAWDOMjga8WDifnn7i76HrKHU6
2p3BzZ+FyhLm1Kwbgei0/urUD9mjp68MTyIl4kDoWoXGOOEJ5zrGpBXg1aAWxETS0ijmymQzfE1H
s0TheoG/ia+QYGbPDfPz4DvJjq6pGyeB0ThZBqD7yOWf8Olm6/2UB7uuENy0m/VyeZOx36u4SZor
GjJbiMJM2saT3jVcLcgjMu+ENO9NdmYDN1He/xNFLql9tqoixi8E3kOzWMQ+ee4JoV/d58ShlLGR
EwCO0flCGVN30WEgjS3zsTfD/UzzfdngTYM/gYV1Qc5wvsiKNz+Nop573vCCQB2fZGdbRVOj1saj
veW6RjdVipIMQ8ZO05V7ffqZBh8kI6YCOjOwt8X9CRxzKGgiELVFoqeU8CdKE6PcdBWGLvr0rJLJ
MGpGDptEeRZa3nw228ELTSSKxlby/r4TzA0GHyBigRarFzvs5oTnt/aDUeIgnSlWgHt+jC9f3d5I
GCcyJfFshrOVNGWDwf/DRVBdSppO/mYHNBMb3B33q5guBGm2cRiUF5grsffTyIdN/rgm6rgWM8Fq
IfzEyZGGtJA76lvjE5Lu9n/5e+t9915BT6h4ssbzLySNMbZZpxRa0mHM0yv3luOTi/Wfq6zv4fV2
C8nGx2O2OmlAh4/sEFFrfaDeTjDr95x4gFmZaomn4jJmT4mrglk7A1Rg9Gl16HsOZ4EEg2ikhAHB
XMpGFh6Gs7sax7f+GFvB4IihOe3RRv2Qq6jAlILWghFwMWqChbc5L29L87gOupij2TdFdCnjA3Rn
jyx7QO7CmdDlDnJ7O0OoFQtJZVHWFVbvgLhd9YSUUbnbUD5Gp6wsxqrHSLJrv7oSa3dT69Xj8zZY
A/Vk3Ud0vBdpy8U4i7AxKBB6/Ka5uZ89C7HH3mJGx5N4O4UfpSDcwJw+oc46gGwN4vpSqGiQphfI
n3QEHLXPQASu/6lF5pcJdpZibbwmfYNkAN+iq8fZXFtKyu5XvdfEJtz5S3uUBFbYZMs8w/TG9kve
C8RqSBRo4Dm2U3ndRWnNW7uLL1QD7fPkfiJaT5Gqa17p8TIMQVc/v9Zujjqyogup8tzTA/o4Xpci
atKd3y2Ky1QeRgS5+SqfeDVG9exZEDbeNHiI2Lk/aPX66eX2uQgkVaEYh4z+FME4QR6QrRDC+9l5
4ZL55hHUZuxEGYt0zyuB+TWsriMmzo5RkvSkCTerunqHMVB8eDHeJ1CuCiN0fG4UstCmqfJeGAw+
LKimK5cElVp/lDT/5ZdlLYGpkh7uT1PDZjKOb/vCcHLivKVS7rTzO2VwUdiQ36nkQMN7wSuoemPD
OwgM8s//4m8WYpC1RePjX3eTqwP0zEn7GGEDcfnru1IJ2JwaVD2Yrn2W8PN8xWcnUPOh+pntpfVj
qMPxtjmJLL/Ma37YLhLpNGc4zVxAfMP97LdUop5YZtEWpSdqNojsSHmg6Jhb7u5jOkJ23A+0UtCb
N5Su6p8I4lbIne8YQzztEJwvfXTbFQsTv/uUZ80XFVDjUPzqMrm/quS6cOpEFcjeh1f/V4IYgpgD
yWx58fJnDh51Ccow7HbfA4sjSykK9EOBhHbsHLqznRRo4kAfmnQKpaR1svlqNlFa7aBR3oM7/37L
RP1p3VX01xWHDDJxkaXcQwb+e5rWYGzSnffTYnfn2GQ3ErBWmf/N0u914PuSrIQ3oN2Al4cPUOg+
59tkjNeEGy949A0MzYMkgLGN4K8Me+c9VLj9Q8t3zZ66b8ZSriJ64ddsvmxBn7tElqSS1S8qSWDe
bJ0rtVh8yDSiNriDSeb5vA8oQbzcbn0jY4jJkSmxOy2Rz76qU9gafT0fvVERHtviai5SUvnh3ADe
mB4qzmTDT1BV+Lgu3/zvCcfg06uUS7mP1K7U3+QyJ61YrONzqJx6H1ClR05pv0iKMPPVSqt2z5At
V8DR6aqgypFaeEtAu5rdxNfnptM43qMFcOxcCzlkcR+SvQyFfknkuih2wQ1RVg5uGlJseGLGGSiU
38EiE51iOhlBBPtwIjQL2jPT5eysiI3qmPVbfofGE9mAR36OiQyxZaixihKdJwPVdsDvzVulERzf
BvXuZgi7i/kleYqlKYm+xFIjuyNREYOHYJMZZ/W7OS5afIn5W6MPStOXRYA0I6b22ClnvvRpY1Zs
ebFT43HoDfmvDGFZuYQrqYIXVgKvDu43Nc67IdgPxnJlJqSM0BRM3a1KuxDSB+P8wjxzEjIqNx4x
Bh7z3AXhT27rainoTtsqXmo6r/au7XuVVttFqVsospE4jWIZdky1JMzMOQ4nSzH7QDWrhhUEaK+W
elAX2wbqr2+rc3mE282NSMlMQu0xM2LZVuZ00usZUahLz+yFl3zCAml3u+BRWKLpQFjdQesnP0Rt
st63fhIdiplTWgbymrdOQi/23qvZkRomQV2+vwbRC+s0pkUWs5MDVCS8KqNCWs/u4Gly9F69hDKP
WrdS8iXcWq7urGqIadSuHmlrPHkggplndqK7DIrqzVjsMTlyUjk9e1gPDhiXMK0VgKztD1hR2Quj
M0fH8KKm+13PeVP9garM4ls6kLtxxLnhA0vK4r9YzSLuKI783GP/SnBAUVsbLW3cFLe7k5ag3QLy
+cHhEcaPzWSgvhhyY0AUW3haWB54V4yV6xRJAkSDBLEciRUBHBImfsdBNJGRq/EHNP5w7hqpBtrN
ElG770S3ox9j0gAUs2mbYE/OAYRY8gFOqO8UhDR2GGcRaVxhTKXGzVWeioptnAXEKUl8Qh2pQote
r+9SNqd7zTMQ+7JMte0u2G3Xh9L08zAZIXCCaJ0UO6UXi9cUhajFPF4tJ9a+f2tfYqqmraGz92PD
3UpCWWH6woFuDluwJi6BZBH0CSCfUPBHxIJ7ZEWx/y+AXiY0uvy9NQL4OUVY6q8wijO6kEcXTwdJ
OqhA9LAwNIclK+Ix5IRduxo4cC+I7Q3qzRGyxSeLzk94G1J1rHXtSMObZEQ6ZTnA+3/GZHvZQpkb
+xsxesigPSewr9coIZJaH8tkbl6w8AWG/lQiedJcArt6tDCm0TFl42+V32ct6NfDStee74b6PkOt
xlegf09Rb2v9E2SzgVk+9AL6biRULJ+uLVlvP9OOGnj8OEjClvbd9Jjh0Pq0KZZTO1pn9BSiJOHr
/vpcbEcYNPyIB5ZDBquTLM22Q+8M4NmX95D2iBw8XSPTENZ1QC+G65oHyliQzvWTLuYK+JGxizrR
POen6E+JWPw9il1ZFhzequBkhbRZ3HP/T7kOeC7DdHcgI0TjKoLBudDaWFLNxFxTqqxFC45ns/zd
U66UdiD9ZnfPQQOk1rx5YdFBt9iKSbPqgYV0iWbfYCz65nckqrlajdRXt6pTv7gpEmVz8uusk0Ef
PjHbRY4Dc5SzmKxx5hfL+/dXDUD/iZmjoVB4Oycm6dsc73HV7GbzknqcObRvYDBR4HlL4JXBy3K7
So/cVUDwJRXlk9T23JCxT30N2KjwT70nzdu+LDxHxXWEg/AQvOkQx/jy/B1L7K170Mij3x8YxQvm
yMIiW8THaW5YE8ZQZIBaan6xeqFwmOBpWG89AgznEtUK9OO2A7d5QVn78+swwXeyFnAp8/Bu1PuN
uFM9Q55+dmS8WMom43qRJjZRRDxMlK/Ycmevw7aVO7G1PWTke3N4+IRWcMt1GOaSSR8zIbt6I9P3
Yhk8FyjqF8ipQda6ETAPD/xjInRvyjNqbAL7P9DK8rIKarr9onIqP51DRD5M2AUIXj/CgQyEjVVD
PxogZZrVtIBNONGIXGIaplam7Oi6s3y60CfMrN0LG2t8RqWFcEsUtqYw3D7A+EDFjMww0KVLo351
VHPQPSKc6TMlcMvVOnTO/76W3RczxD4fjDB38SlzAVES8rOSNSMqe9nH3zk8bjRp/oj6jSGo9Tdg
AMqEAItyRxDqTZZTPHPKoMwYqzkrk8PTzpb3ZwjApcSmI9zr4Nd7vJsnPaXZykC5fCK+67ngYcdM
ZsgMN2NJrcO9m4VfEKFM1varl/UWLyjea/VDa9CgbbIVAXNo6FR60UIxFgZ0H64E5Qj2g5Iwtplf
JY9HNzDVlASxLCv+1Rx3L1ZudjvTJei7NMoW1ZSJc6lJ9XM3bgS2VkU+Id3Kjv1OlFim+o2j0M8e
IPGoN4O0TgT3HpjtBrnr63VfncZ6yNpZzBZ5D3OCO89+3SpXjXzj1jbxZTb6ET0HU59dxSeMMssZ
0b8Eee4vEvzGUChfH4DHsQ9xyViDPzoEEsSMhb4bVgodffr9BPDm4uC1KW2mGMsmjjoo335WZvs1
KBZmH0I74HCgbsVhA0X8cOTQfRg5S5Talbk28c6jSqc2MxV13lJNtvI4yykgQd8SzAqG5JcnqPgZ
UOhrYpfEClfn3fPJ+x+uBDcNzDIPnDdYJytOz887poiV2QxnoY88J7hdbZkw1V8kg+J0SwFeSCAn
0y2UcvMAB5V/4SeLb4CBSNHOJV8K3EcrDVg6LdyUfrCd2fJ4GoiNtj8Rkoy4Xw2QTPSgETh4UVHZ
supXVKY556qO9hEzK6J6iuhH51vnm5wSvj9+0Dz0YZ7iSCvuONGLKxPFqwnhu+UD5H0FL6/5u2sQ
4S+W34m3/v2QmlJ3+xmlZOZr3rLH2Yu96Of39kh7owtNdyTlxodXSbEG7DOZ/pjhSp/CoKBYvHMQ
Wu+C7GyLc+YSSGSsHb9D4Ci1nx9pMCdMMGJ6l7BERtoiR4G9gg/VVK7s+kyTC1+wfyxi+/dH08nK
fUIrZ2TieGYbHWlUL903mdmrxP+m2SwTyah8aFCV3vqcqoy7QELRBvDVlwEZAYiwIhv2VM1MF9cH
Nl6iGgd5SeJVgC88eN6MCz5r8o85kFrCxjevyHvt/wi+hgG9BFQw+xX5wScqWCbMos4QoiGUtAQ2
pwcSKbUxs95tiTD971R73H7oSG8zBBXJ3W4jVMSdUcG926TzSCv7oVVsVpjAdPv5oZr9r/eSNiVS
TmMqlCQZhY6F/39n2ddtp1WyiSGz3GetKNwu7FgnXsri0d7PP+8gwzIYCvnzgTz23bnJEMYhay0V
zdjp5y0i5C9FqhZZW9hX3UI7/5JMYaZq3pOFRdp5CVB1VbFhtYbLIGbTnoTvx9K+5H9Eng4vkmYl
rdRaGPV10BhkXG63lb2UQHKJeFAQFJOOYnxfwa8LUHbwS7rGECVOtCN3Sor8k6hFzafSAi4h/r7f
vzx/o54ldMIc2fRcZbT+WoMN7KnVcVsx7Jg/0We9yWy+KamJzHul4UwS5P5a7/4vOD1zU2FHXPV3
v//ks99bWcCJQTw6LOHWE4rUnCwQ72X2yw6A6N9fYgnH/02Ae2BUe7D3+6apzybfVX6n9r+NrvGa
ppKpKrJ+dd3xMyxLRuO4bXNpKyoKEm9GVLEQSZ96lZmdVqLM6Hq9SU5aTkdGYpPi7mSedBqwsDnf
sGYqHkwydsZvSVxSqymbm5O/OGi+NgtHp5mJXKGPx/ksMIPWDNhPvyjLiP6jBfoeJlNdKUkLZn4O
fqiEHjc6V62Qo0alfugj/+oSmKn3/HxlHzNOx3FNChOegdJjSxeDLlSGAn3ljyPXXH51iZgosm1i
6EF+ci+QUszuBJL47k9Dwdb6rCiKwb6iJQ4KfsENP5FQNrlKQYdA654rn7HjV2w86Wx36bbOLFRw
viYNV2IPhKLWCrMg7tzqsCVlMMXbPBBUP99meHL0IfiZbJ5N1ycorqE1W8NuXQy5zRfKS0m4cIpe
JcZrw3gZWBvVapMvxQTWPxHfMKPVqePaRrViVGEgRNLuUYL2lQB+QkBCGnQ7eDswVuTm/48TU64A
dqnZuwygVYbA5ueIELT6EEROBGmaZ27ZPGHoDz7nhyvFz4ZolQDtCSzF9T285R/NMofyMgc2h8FW
MixtuUzImJZjnHIJ4ADgRxMwQOQZ9cPIY6c0Yv9/by3hnL0wOgBGQ8OjP81q8fpL99IrNjurPPhG
MwY1tYnQ4z19FahiA8Yq5S+lxlXn02AfyMG5Zm5jEoEXtFWqbX6W6WihLQQlTbhRK+tXmEe/jxy1
uNoPxALYeABybTBoS0R0YPoSSPoXN9DMwSPNJeZClcu8uKpJWbIcBmLaLI1HJ6EUoxN631OwZPkf
F+N12rbGdTImVYfp7uSj5eANeL0HCU929n7H5+aa1wj09bPxFj8fRHVxqdIyDM0vV6WRofxiz7d5
Onfs04ocBc8HrRDsxC4Xnnou6np4kdayE135SA6xJ5rySv+/4PL41gA8TgX4mCwn8Hr1mESV9mfR
MncBJnFQ1qpcs10RVoEVXFZ0RwSy0meWHJb2gsiO0vdYuynwaxgkGYDqi5D1JVLzHkt2yiAlQ6l7
sq5HP2DzDXfh23F+xprAvFhAmRRu51lSGaoZOOjfpcsE/Vd+6rAiu5RH+uw4Nkmd0IYVDezf3n31
PJT7LTdqI6s56TzQQkCfUNzkhdN6lbmvBMJXwhbaUW5+uS20ND37EkEjcmTQl7X0AEdrSPBCQFox
rcpej+a8C4rYVHPd+YLinNIPnH8cFnxRLNvrI+eXzp8mTm3QpcWqmG3wwaAtreSn3u093wdJpkhy
YJbm3fsxIQBpDBMmlx32Ub9aWV6u6sZH7l78nUovi299w83Jr0N0BiCFfS69psMJWdAYyV6WRXsS
OMqTprUIdhO2vIUqN+4VQVP40g5xEC8HVK4RsusJ29yUUJ1/EA8SxFLsNvDtsCd9UBxtnt65b6bx
z1+eRsrawPDfENB3HE7f2TZBtXKbfAW80gyIa5G+Y3SvEH7Sp0XH+Gqocn95E+e+5eQ4hvs8I63s
z2ZauoM5updBiBrSImWXo8vXGb3z9jYTm7dezjpyUWvDgFHCZ2+9s4Hsb+qgxAXsOPZlPSlYqxxg
Gb3Mz5iMmtBgEXBJUNP7wkyVkgN1s5vhvteFs7e953HVq2WT6UQ7ILv+hBdX9yS1y36IZhfCrS8G
GP7G0+iW/+wss3eFwd+kz7of4JWpk6BLSTOO2K5MTLaeuq8XbBsEDTLqWILOAOA/RHr6X/QySa2n
ypbCk/ipmNzrOAIRvidbgA6zB36aaws1kS3otV82RYdeRzmhhOTgN6k+ZYwDYepAqUx38MoeXf3r
apwtcy9JVtwVafP/ozpmlho52HL33hs8Pmll2HaVWP/CZYpjR8snL9HkD+CPq4HlA9zUpG7cVAqQ
ItL0ik4yKJJzYag8vT7PC5huxL23c3sbScaJ2Dk4HK/CobZD7k5XnQAAo51INA+ir3qPwDkay37B
KWMcG6fhDIjLO0mrSnI1018Gp81NURLWG4jC3pg67rr7f2HDPEQxxJVSf4cw1WdtaWsn8Mu6JO85
XBc/zWBf81fx0+Qz+qv0EDZbQ26CJ/+Vc9p9X9+h+yqRpAuTGcFG4k1AkaKoq17YuethRbP5itbs
/rxjm5o6Z0SKPb7V4cGHGx5hCpyB/vyMKXiDw4+q8K2usiL2t+ZApYlHp+nlOtDlGCsUADBK2VCA
FiSWcl36RVsQN1zfDoq7545ZD0haGXZRlzraWaaRaTMuhDutraddi3T2NMQw/Hk2CJcW5LOFviqx
cvX2UM1b6pN+iMG3BiJ2ns7u6tB3C/iXXIFCYne1pD058xwomt7/pI23apARH+inzcRro55Pkl+i
jI9poFjoChGq275V/MEW2LfMebbYrGP2R1xHXIBI5W2aWRmqUMwRMaFXbwQw5YPvbKixAwhwLaEv
NvVk5fjNuOJCdBWBW/eqEzTa6g8788cSFjFGTCBkRYlpqEedM351Ix2++qLq7melXsoL08yKYD6b
9GvC9Ors2Ky77WxOTiMOiyE2m3d8jEo0b3cNIwGuLu6bK/+j2mMBXG7JGUnZl1s2A2gwuDZKgWji
XkxSZ6XgIQDNaf4UtebD7LRATKKeFtVz6oY7fw8PuKqa8OOmDMG/W/6lo+hoIlk8e7RnNBhIl5dl
XgItZyGHri4MRVy+n84SRg25uOljGDHzX02ZERGWiZogwe8LQogeX2hZHBpkxVoOIkZsJ7n9EdYO
FBr1nUMvNsKG45wQs3TFSRl4fLOeOMuFi7tkjBGd4Ap/ub0XR1T2SZe+OEqA+Jcfc0ElibqAseJp
tgNoctROaN1wHoYAWJGvrldDmfn//KTGK96dCbZYRV/g6AvxOiscAIWKJQuoKHF8Aw3qNgp0YgR9
KdnmCkwp4OACRuIAVT8fB9YHfuw3kxBL8/QZCwAwodezlWwjArfGKIehUmBxSj/eU2ZvLHinaS9t
bFd/EHYq5UYCGz0gtU1gbVaBEggil76Z+ojbk24kOqiqJxL7GJJZsGvNfNNylGqn2TozGJG5y8W/
CoXe1hlATgiKD2hE8RLv/O1AaOV/yfWvOIQQAzA1MGZy3zVLIZPy5fN/5xuTFdtV0xPu8/5yfq7A
W07IDt+T5Nd9ANW1MatJLtvEUj08PK9PfhIbD8iziqRcrrX0rkEyL0IQ7Vockfo32TCu/VJemgfw
Z6odDO9Ex+/w09HMbo1udkD7GUkzLISWfJbUSvnPV1H2afV+nDzbidn0fsgPa8kHXcuMEhoxXV+G
H6n57B4Yx6cZI/y3cPGNBKMB/NspR9ZWLSI4lxQgAdM00a5BDgSxIjL9Cl28wlyCKPiwhf8hXUqs
vd+ngAxoS0RsoC8dLwDlEZi7yVRcDw9dK1iVb1iXgnaFeYRNfe0CYM7iZ/xtANYk6OY7dL5woGbA
bD7TYfH5WwuSvQ5hVNJqQW9O8lo0m3rgJq9y7cLkhUbomZEsx03JaPxkG0+jGDQpw6KLQzAK0sqe
vYpxE4EakkMxlIHNBEKTNDCJ5hI9MsciQa2kUXoIL68U22TgP4i5BhSEYSqWOS2dAwxsUbMKEjQw
UqZD0Cn0fpTLeUfnjGFxxdeJvCD6BdJ6YZgxhDuet5NZxNl9PuClgOOdhfLsrcJrdrYW+p+ggyVG
AV27y9bwkwFduq+9bmcJ/fvRT8W3RaK1tJ9bWWDMhtO/h+UqSThg8qPvvik0ZXoNgbH6h7RSrdfi
FzQ0oAxCVf7UqNFOfKiUYEHv7lM3Dik2lSCaXroWQfCL3sqCyZvEEoLWV6+/jyJSygaN2DYiJ5Dc
Ne5bhN99DKK7pzE/s1ykDlG3Ci0AW812fvbqrkTphqbS74rUU8NOKqVDAOvowARqjpWAW4zSBN/o
Hiez/NEvzpZb9DTnqnZMdnlXwkpjrZZgL/XDL/+W6umkk7lKF7Fa21sxlUYsvm+B83Sf3TzAM2VP
54OmZFoK1KkWxC1s2vUHdWhu7sAKeC8Oo7n4x7EtLeisv7C/fOVk2vUZb438vAOEGOFkf0IytrMn
Uj4BIjBD/R6yHvP+EHzn/zcBzHYHUcHN3cwSs6Sq8IKrpX8CFHAyOgQazHLS0nJvKzoBSiwbSOZ0
gbKFq2+P6UcgWrmlJ2kOJqFdkoHjs+11Vq2TUcqKB08Bx3jL4x/O5IAdMESMwAVrlXgOcA6a+14e
yOSUAgPcvvnJE8gbF1rGk3A/UvXz9SOPH2JO4O96kJJZUt2qZ1wqDgmWhXbNqIz2yaVBnDbO0wx/
xcOkxnGdrSPXZ03cmi0pCNz8BKyVXz8KGR2xzk72+pzRA8E1Z5cxhftb132N0Nhc3w8cUYhqtOJo
PWOAaJe9SpstG3WXSxhvyv72HvO3I/UR2l1mSEYydlbHwXfeXTuV2LkNcS3Td2u2nY17O4TAgnpa
n00KH6Dq6mnnmLo8w9qNbYU6rpuC908tyClI0LD265V2B5P6OfpwiZIRYQWHKGYjKHwc8SUCqnF+
ruha5/EUUZ1HAgTrP0IUaDqmICslOaE1fO/QF0ju1RqPRMJGRoGxE83st/iVTzOfzCbP4dZ8dlLN
O9JN5UFfYo7T62CQlHf856jJyzdKlvmzgxxWlIp/kAQi5UUtI8Odo5P2pfVgis/azt/zz/MfTYMy
WoK9R2pGHjMsdqRJVUKMhB/tJ7b7rZsdzsu/bwN93qQI+8cI/xkYJzXp4PtONUt/qpCJm+hYkBVe
axXHo1DtDcGZxbu5BGbqpBYdXuA1U7Epm5VcITmUz4PwON0rd8dMv+9uDjx3xzC6cnD41quVR4Bc
h3zmx51GqfqhdpLyRhEwSTakTDQFTiiyYMShXk/IN8uLRWUrdrLoNDSeO09GYWj5bgW7NG+GIwhY
U5UTVX/IRQLCaLPJFpFQ8ZtYFHDTLSu2wlAoK9m3rAW+BBRm2/s4KNAL1XpJjqXpbBBYhkKRpbkC
ORkZAJDS2qjvE/ubl14TIYL+4JcGisxQrcVDGLeo7uKSF4sxl8/7T7GjTtK1PKr6FM3N4R+AWnFA
45Rc7gLsDT/8BWB4AXTo2yiL2q+Kh4yU4owfdOeuuXwnM5E/O2/FaiOtGhETtoPV2aROUVhKKzgT
CJvSMo+/jvSWfiZMUdtjsV5KR6MLLqUIbtdaeECwUa+DN2wppxO8oklutv0RuVsMxLt2tZa7vmWy
GdeFuTRCX4eylP+32FXcwcRcLdINULa6UEvHNxt8ZCAzf46RNVv+KCVThLgpWTkzKCo5242fZzfw
G2xTFkC3bqeUsTAQNk9C2+/SvePWB2dv6uSWgBFUNM8Ih0bbBt82j8KpirU7i8+ptphrzduYNrkQ
d4USeAzbZl8xjaCO3w5/SeeRa2v9g0HXGNOYlZgXKau+COUy93nMFu3wzr1k8c5P3WB2hlDijRLn
b16KNBZB5b62+iZg/G9usoqnghP3rwFzcpzcKoJZH3VOmWwnRnzExV7+6Sjul4s4C6pkUm0CKmGf
lalegSNOShvk7mprEi9PGFc8CFDanoReYXJMHgKpS/vExuCDPiQWNUnGYmm7KUlt6wIlWCx/pRk5
2yY1FbRPfMyIpWi0IwX3n8tBHJIHkY7zVU1UcSfIbvBYs/j0KfkaKPE6oUnPgf/Wm7ptmca600K5
qJBOFPHONoP5QT4rafvEwYbf1yKhdS5RLj2U5jA4toTL2rgdzgRIB/Ck6ZhrH6tbLH8vXiBb1jt7
hejQba4xymOUHbPvlb2I96AnJsNx/0NtStpS3apGnt2OCuYokubeW4EIEfkdIoO6c2TMWO7tcb5q
fB8pQVSnAjISh2Pf6JvSVCPitvBowNPq8UVHw+OqEoXqPf63lOrdKt2DQXJoe4a4w0DNeIgzl2E4
07L/i6DtjOpgngqwPJlb34RiY4QTjBVddallERig5TvqY3hmXHjO7aOghh7igzj2y+yIMZw6hO/s
Fb47xOtnbhp4fZ6r2r+/RvXNwZbAzq5mNZtf7zq4TU6hsfb4JWvKaD2xUcgtYSdWD5Am0eMmRYI6
g3x3mUmEIfe2P9bD5KGI6N14cNs83EzvzrJ+E+ePEjdGhy0Z8NyugkR7T2Px94BmotKgAqGKld/w
bgC06dwnwsAb53P/VI8oItUR56a+hklgcKHGNZZMUgA9V7jTJKAFRsjqwDKslr8RBb9jKle7fv31
knLYw2+Te5v5CKOVVfO0kwgSTTvXMotkzLmHSssoV4vcavgmB/P2ppLK/3xOtayrOAGmp14glrZd
fntf8m9zkP/NTwLzhAbH8bqqDBQf/nRqMZwao2v3CdVz/Agqr/zBr7ut3zadTRu7F6U9oETxsjTd
UcYcrRoyH+a9jQMQRNTE+/p63rJ+wMV048uYcrsNiAQrqFfYoAxSXRV9f0EKZkdgPm/AUTvbWZ5y
MmgXVltEQfVZNOL7cC0cd6Vi7gLVlcsJWCHaaDQrD/tiewvpYGKC5GY8VVCn5jhGC1Vp3/vVMUxw
MmXAXAqh5FTnfY/Bt7QfvYtFrZEe7IvB9WkkJxQIXphQwrQdOdWx/A8AH5cX0+7o7kjH6lOybJm6
ZCh/Errg09j2Bh4fWFCyZlxAX+p2ogtznu0lsuVnVSCgctuX7Z2A0/MLrHVbMFcUx/+Gf6r9IBGF
sNLYF+RufpNrQ2VgHZ4DioCQP3JdXjTfmiwjgY32iJGJiMOhet2djPOURexo44IqlOlPl0ERTlXD
W+U7M/t/EzQapUXq0ICDEQgLCYYuhmNLrscN/nSplCTAUXxlOuovQy4pyLEPG2yugTM41B7EKV77
zDAzS/v9mhfT0DE/SlCHVp/UwL59xmFsd/e8z+EU3iFhskHQIBHqfzdQIjQNfjpjw1IGlgQGX94Z
OY2Uvc96KFVuLPOkdmXEy2LyxtLCnTNKEjSaQOZ8DFTjoaaSTHKV+rFcT0J09QJOUCur0WyDJyQ6
IKtEOzJCpA18aiYhSBVXTHerQ7Bld5NLRIgPsvaDhMlu8fPs7Xt3OBW6UjfjMHVOiAb7Ic9WoWJT
zKkRLb4/l0uU20n3XVgysfG5t0tviYvfZY1uOWEREB9rqQ+FW4TB8y1BoAGKo180OuDwjqswQs48
wZZQ7/4Q5f13z5gZgwDO0lb9XBnbnSMnRjY2WSHW5mrbSmGyWdJhQKfmYVHJ1ckFGQviL3myhMkc
Vyo6axN5ZI6+KQWqsWF4eHSrIKx5xeq1ziDN4ZYcjjdpXbVBpxg96zyhIg6u38xAGR/54F+UZq8t
62zh0MuxWmRk+vzdy4THTAnp6stLPndejLnrsymjU7lUbRZ0ANJd03lE1Yu8LOpXKzU1/pdcDTAT
BMYBdrM9QgoiRsxtiGH+xSmMRqXhlStPbkxrOcfMYx/rzgqbHCmU+9Gc+8qRMeusrEC+mVSb1Gi7
2yH4pnLbIS79kQXT3lFW3IncYLq5+UKsr8EZ8ESpT3K6Cppho08mREfBaOl7MZ2efGjcZsLxrB3q
E3RbLfDvC+urKUihW1JgG9eL1wYW+j6CUOSDwcnz1HEceK6dxw9IbY2EbtTEr9Ot6BGNunIzeFPH
d4Mv6VF0WxjZlD6spkN4gO1o8SQrXfwxtSxJQYnohRyV67JQvS8RFWmTBT03HE/Q2+4a64UykZgC
WoQgntJ9Bc5gObuO9SMwE235ttQvxZp2qriqYsX+T3bHoeOBNlJohA6qL3j1An5NP5Y6cWXuFZj5
lcUVj7ph+fbcinVePRoV6olr7n258qE2aVNVbT9YnH20d6ERu2wYI+jJWfbtMG3nNxbjGU5iM7s/
suax7JXt01ovjeSGsAIyUeadaBHcUHLpZATzwAuNFImbfRmoYGZtcY0mtYELXkhwpNa3TmefEBZb
AsTYLZxI4UsWMhHzfCOiMe7vnPbaUWQOyUsjaAtLcasjsJ49MPCrutSD9pOSA6dX/uK7kpLp+Mck
nKqSSdlDLsmQ7bKzQ9bV3TVsPKMA+IvnBi8HJFg+tew/U8ldNxBrRt8MbEMHmOmv9lMA/ypm2dUF
rJDP0RazM6/qtsCwQ6Un4NFUR4EYANP3CcqcBGwiNPx3zdhN3UKoditjVLet7T57yxns5HwylsFE
0wHZPGjKYt0wz1EQKFdmqq0Wf98zYg+SBQ74rYqZdvMH4AEk9K+5i64Y7W5+vZmV8WBAgkn/C+ko
uQOfzS4XmzxVOPzpn3jWWgJU5sngM9U1dGrq8lX6DWd53wWR+c2HOx3GK0S6ZUCorv8ox/wBJWOZ
kEI17kKepophqbBakNKJU/yN58XIl8TGq05skp5p3TQktLrAytJQsymZxC1JLGbjdzUVy5KBEDu5
2O935RXqt572ilwW+RpWyPyfcKlxdZ0uROA0hx3LxH7fTP40aXSKGKPMoFrI2fNpGvw2ImDpu6Ti
gJW9sB/A/OLhkWNjXzxX29HkWM4kjT9fqileBRFXE9vhCnOp+2Wa8mgbF2hRVNn35eLIW7gcTiWn
9KtP83026QsdFIwYXQczA4HdV3QODBJtxrXsIfrxu42FXN6LCePUMv44A9ypSUq3WmCDyutKnDX8
wjDP1BUNEMtIoYqWLs8oycP6Le30XoscEkLFbakSDGmmlhogbFSJFrBvSgvQr1jtxZeynViUuwkq
UjEfLbS9zMA9O8ADYos75wU2eL2XpfllRiKHl3uZI7PnRWC5+vKVCYAsOe8h7VzbdeIpqFKnGZhU
BA/b2PbLx67OWly4kPaToI8CUgW8l/dcfUQiNAhVfvcddH3XmUM9jBOLD8phQtm9EIcPoyGi4PpP
V7brXLPHjj+/8NHhENbtGxu91wSrPhpaKQNViZLGUfKgCft8Mk/q0ZTIAHnRuG986tTttC9PHeJ3
rJCVW4tvEdcPAaAfO+U+qy2XCPSHyv8mxM6AN1ow+EIUCaR28hWI6MGhxdlOjlDTgDpDay71e63U
SWs6Z8eHzR6AEtvqs+7XIIs2pEu1XpR0Q3ZoLg1NFaWrgTNRr42nR3nchMM5mGqblVnTazNcXmW7
swxKX4kLkXw0jpfuVZX3TwvFQTYbvzEVACpmQUJaAKtNisNWU5m8SX2rYx28M0KfAN7SwiK5iuph
LsGJcd2fFHE3lkLZeapAtgIUDY/bs6VUigoz8G/D14vKFoUWkE/8I0wkCMthqPs5OhaQzE7gNjuN
cibRVAxdqo2p+YiKfW16HDGceLxuAhQoeLHN5LI+f+SDyQNbSbqdcoNSL0yZz2GYsX2NQHQnIiSN
ail2+8LiqVM8KA9D4iSJ6sscGdVYZ07VqzI3aT3JUKCbGy3+C1VHvAlbRSXXDaQ6ywMu00VOPnTS
HwLze35JrqM39kyI464AvIx3aYBaHaZWI7FebldVFBSWY+GSfl0Y6Jkur4rExA222y3E4XL5x1fM
8YmcXWM8Iln+kRHwhQiVI+JhoEC+B9x0F7uWwPUNDsHWOcAq4ElXpdPzCF2KDfSIOru/gKG895g8
FLYOrDRskI1De9V+VBiKZ0YX9PC7iIMDOxSu8wtRL6AFqoJMcZqRDFRzuyn9fXXplGBKE/ayqjy6
wYalwInr+PAH15lH8jKCF/dXTSu/HFXgXA3eZX8B8iUZ7CnrBusd/3OT6FEKIqC1WbxezKQN1ELO
4vNLx9j+YceHogbV/MNnBVI8vAmQSQWV4+tj+d72xv4wjYBik21XYwl1obpYdV/uJOi/WcVE9/BC
XFoYkjdoKdTs7eZRaqBeVrpDyjFZhNWX0/57Zd8zXwb13xyb/1E9Qr1y9L8d7Umjp7f7LbTDU76L
QbPU7BbSnxNh5OkJXYkbcrW5nGu0AaXGlpnNWDL0Bw6rpfQo9+OE7Lp2Ygl/cGHzmBt4KPb0Ef1x
8J2HrgPtMwYJbYYCFstIn79hJDUyrgtYsTp/xPiqOBhmDUZP+zJ9xall3rGQmBKnsvnCyle1Gitn
piaEtuIJWLaGQko3791z4eTsSJFKM8IiyWmENWdDDB7gVjiCaJnLI9c2KMclzF0IkpszyIow9F5S
cCdkzrIk0SHqmUi4atpg3zQNAEww+HdmFAYZ4EqxzxTD8lubsW3zYre3NqrtyufLoVDY0OLQe6IF
1AiLIqtqiSKB7zZCs3EDbYq95dt+Y2zkm5cPXt8W4kRcFszET5X+Oh51HtxZHo8tODH6NdkUkYyD
GJWWf4wQEqp8Gcp8281+wWP4HC7162TapdJ5J6uU66Kbpd4wFgQhX5l9dd21X2bDoyo0FKjZkKmw
9/pvH4AWQGm+1cKAosXoVsmxj6I7/i4U+SPU+ltDbVgApPOLyJnlCURJtd5eXTjuIsR11+EWdg+c
xWktma9EUIk2siD7S4srOvOgJS6mEzn9zPnaKxWo+k4m4AeHcbj8ncgKujqrEw65/a34SAJ5s+tR
ZpTYINR2e8gWvq970xwueuS0uBGJ5VM/magcO1ZXX6JwwoFRsMRrtfhkV3f1GZO4gh0nvXvRFUau
Cud3JDlO2DayIUNxSKqVaHyCRLhd8k1pykpwl6EECjLebWhKocYUVIos9+RGn8YcxgaNjma6qbVH
Bh/hvX28hINq19Qio7HdbZK/YAMPooH3+RxkebRpoxnXvtssF8aAZ0iDSsTX2tW7vAFAXpSW5POz
axfVVJVClAVUnrxRGLp50Mz0QOeWXU6x4Z5HqsuNhSjIfFytWaBKhbHTv4zzqmgJf3a21zlCeHu8
o5kC2W75v06TFcX3eRAo0mx5GCJz0meMdUBvxG3b5vG/8AlegKOGZjOzIVuKFwbfqlCFAcRugoYe
CHB+JiQn7FTx1vpC0PSO5Mu+Qk/1PbTmVeTm5xGbjTeOk/qhDlkwaYGjRncsDjuK/gmOjF7BI/CZ
QT4xhJZOPpR2k7MEh/d5fR2H8tTtadVKpngcjy57UOXhKIhewFvnlRXGjKYqqA+ZdMgvSPxoihie
NjUb8hcZ/KttErXCueKoljMJUUY6C4kq47j7MsaVctbD2VjufAcwh6rg40FqdRZMguBVTll8E+AN
q2pKpS2CMvJBZLlQaLu7HNtdeGk9SY0KXV6VG1cmUkEuCpJ95KkSbEXGU3ACVyF7REd+NYRITc1n
abQdG1GJaJXmObrF2mxfKdyf0eDiueZ78IKQq87L8eIjKy4DVBx/Wv6mEPzfNCtmtsweTfmK2xYf
GoBPfWFWkDEyt8fXPXlpXeaLdExhGpPQn6WqcMYiY7kdjTt9YOTVjqwj4uj0mIhm02hVdNOZM3tF
sMsOtw4wn3r+tUQo/+4iMs/Ufw8ReXnf6vzuz8Mle0Lyw3lMHt7qkwiXx2g/GC53c0iIaid4N5cm
nFCbPUQHa+CyBoP6a7kweLz1QO7iMCsqCMcQRLTSY7NI2bf7TWc8O+JmfC3QsVowzf/sWCr0LzrZ
c1VOCdHVtGbVQKPrRwSuXCz/GckFRzt/8gZztlA+vpHvubmu9DYwy5k39D5C2fpIwhlLBWvfRBUm
KcemDf2dUUEMGnvyCHogVvCpmKuqW+PqX7pJ59sgemP/ifoAy1YCNWrTQHn7rzLj9w4vnPMDhi+S
Iiz0kteoUJsU8YZ79HjOGdl1al1a6J5lRCdsnt1gBLDGEiUPcApGVvQzh0IqgbbmJ91XxzBROyfs
H7CO0dgvURBKizCcBr163GPs2IsVoWESRs/LQLdr0WKJNETyvhxOAsyl8tbQefyK6UGnqrdTLsmr
g0Ddh1YELtwZiFQJ4FoRDvcj+fO4ag/aLccsgDGnbtasw/IhxpYKA50ktjQQDQ7PHgiESxkDLZb6
1u83piszVhjumJ1ZdPEvUN4lS+3BhMXKK7a8B6mC9G3a7vDa4C7ssFUqbFzed0ueeksXMDgipYZY
mp2yZma3ABBabkkPYwiuFfgcwz1LEThp+bLSHwHwhYtuJlZQPwIJKAHyOnRP1X8t0yJsxzxBsBhG
kmLzxCuwRxnN9IHiFKBmLkEhxO602t+oa+s1ZxYUIDMGiPW3cAkurZlTFeDs66lzkOdUj/jcru6V
wM+iUl6LgzqaY3WLAGCFu24LHh34FDTsEr1tq5MxKSOTjkw+LQUcxSij+VNXGgGZLfpQBy5Anx3e
xPhQrgg96Iexsk64CS6eyhnRRE2W7CA8glyG2NunidcfGaDVsyYkVeYBsgKNy/dR8NCUTg6dex97
FjcF5AXXYrsrfxzfJfHXCDD8RYxWl02KU+QKjMqErB44Xeg6YSMJM4xxWKCpB9V2EzTj5olfa8JL
9LDxfJ+iwSE9VSeP+GEcgByGVqv3JhW0gBldOH08no9MMTEcaak4k7PI/nOkjkGgh0xKjyeLgQbv
vayucHokZJTX5ecCp2fbH2Id1c941V76oKtdGPGi7xihPsk8CdXyJgGS9CWITx16FQoA1La9yoiv
6/+SxyOdcjbwhFYToMtX4ymqSuMn4fn0VBZ10IUR6Stqfo9IkxOU9edRo2Wx7s76++JOiWuQn2ij
cUwbWfMB+C2UgvjXjGIlNiVR603dSfIfYb68TMePy+G1SxzjqrbKd93dHmnyq5yEsg+/yuMdbIAA
VCP1LjNF27SXT2mmG/XQYvurZdVWjwbqFkNsjimpDpwo2o0ud/V3GCzyVuv1XL8w0fLY9bLRrU6Q
yurFdZE5n29FAapzufi+EHWz3z6chtQBsrCYvc4IFMJ985gh/D82J5ruTb6cMWJIdHJ5yCXtcleW
IqGTTVlIw97BWP1iIyxEZgKBK1Iyae3wld1y1tcuLSg/aucXGrHX20z6p1d5aQdfeTj4BnH0fBac
4ujmUPHKLuGA7GVLXDAURXE+66xYUbfMOsGmHZdWEwCnZd52V9C23oN0yqHI1UQWIrZjz/dWA1LV
YswYJ4r3TJgMOx2nRN48g7C1rZ9IlLa3TkC+7zmQjRaqD90+sj0yvHCm2o3PNWKhYaxgLeXImI7b
I61/gPvHaAPRjvN4Dwg2ZQoVi2TWAp/HySHlMk87RXJDZhqVDRinwTaAaNKXqcOkPhEvtXVw3OSQ
Wx/Ex/EnnNdQsGXsKSmmhaFnNcBqVYPWaur7omGnJ+JEdE4XqZPuZ8UF5Jd/itdLNHu4E1fiJd+Z
WNAW5zzzvbgkdeY6NtP6O4ReQslQorK+NBI+RpaDvVl3rcZc/3VvlaFzv1DSGyYRKburvsrjV7St
eGVVpVy09SJZLOsNuuWBgXeHxJ9qh9JxZgRM2Hl7wVLIfqgPgf/1yPTMDUSaKjxEGCxdJFjKzc5i
tmOTsSk7/124rQ4qHnc9RsI5Z83eh2c5xldWMxaRKAqqLmNnJ9c7fCRe2ZUYPz7DoeiNTAnFfrzi
kYuNvCQzSkyzW+TZipep8fpl87ACt6ZsfniO3Dm4GjAG5m46q7ljejG5tF8v7UlmlypBFijiTnr4
sRnQg+epUPulAtd788S9S10j5CAjnEDl2upZPFeNc/eH0d/6dftZ2ob8NhG3xNpJ4OBtYQdKjlHi
oPELBaNk+doZpLWBi5DwL33A4I5vZpdz43ky9AZvMkadWls1ciZcuIFHd9T9pmXOx/RjCD7OHr7Q
nBVU83zbfrp5u64mabxzqwyeUMLL6Am/nu1Y1uIVvl+BCH56G/QOm5VHv//bFvc+GgUWh67dzK6K
zs/Hv76zdjP92g6ZLLef4EXU1UTGEbrld2A217mKjf9q7TYM7fmYtZyVqlXkddD6V7bYn/HCBC91
7FzAZ1qdpJ9DSd7gCUQ7bXVfnJaQTZ9RZXJQjPBHy6AtRsDNDBfpW1itnxmdGAF9qPAqMTFLFuv4
N7NbU+RMEhaGKLUauUUjxh+aDvL9uNdk/TAbhzT6/l2BrCDTjKm0YXPKhiqj1ZLxnhRLJyc7PTeL
zgdd4wZwAEeI2vc87jytSulAiW+/3hCESoxqLaooQv8wRRCS2N+xH8+B6WxeLzNxDriDbo/I2W0Z
Ehmz+9EbpXfx458dmVBfLDpRBW04Uc4fT1E8V1Jzw2XIFkgMCRwO8uAmkEtbPz5qPsBfhbrrJ1w8
Kg3knoW5qITrOUiUwuIsS4gY6Akp2CzXB/CcaLkNMkl9FKr++GpxqnmLQnke2KQKlejFSgtP4qQY
7e8WPV7zAaNRn27GhblxG9nBRwBgKxAuxZ54p9FRFw1RG/PXFCWWwsuNt+BeOXTSoaTcF+dmEM6x
7uRZtT9Q9IPOmQA+dXWY3sclueg5o5KpgKP6U4swMcMZX9wji2vGYl1NjpK2swTKNCiZ2HS31fRr
qXf6Pkg2Wv4s43NmwOZHyt/DlIanQi9ebtTaV2SUpG1ENRu/LdD6F34AZwm61K3QnwV/ViPN6eQH
fg4Pv3zScKedPQL18E5Akn8bh3/27zo2HtIh60f9Y14JANvsTaZvD2ghJ1AMFqrT2BmvxzrWqgej
lX7rN/cNZub8yNUWUJJJD5VlA6aHBnRdh0gBQbld0imC6azvTqWEul3sCS/B1fr+sR6Wl8F48s6y
v0iYzaNRvWw0bNwq4zumczKVIemnrOposTB9UwRjSiw++NiQAXdmDgi316jE5kQkW10qy5gIRKJH
rpBdHVrcQERGOvaCmqvd2wFPs6XZi8XFhWPYkyituF3fgxZiOsj/ycMq87fKrXkvtr9o/aHzxU9P
mZHZbmnd5fFXW/vXV9TgfDE10dkBg/hLTmIeUsxvQwDeQbtMnwIud6tZz/rC1GvnV83NGw1kxuiI
AmAIJ5P1+9ZqygP/HhuULcSJAoDWtGuXah+kg+WqXPWtrkrQuoarhrXowd211OyM2y6aFDOheCY0
mW+hYmb2iJiBFBGOZ5jLsMYWdRknxtPh/HVQ+dYjldYt5ybK6IjbZ/yyEtcbfrxayJOuKQu2eK7y
q3ePHqB478fU/NOfTwgQ9vYMNRYonskcUY7YOyOZuLmHOHPY3XqlPXyxi0qJvwE4lKAh2fx8lMPi
fNIwSJj7B/RG49JRevZlrtcktHBBeXLcBiaVzNnxGdJ76wvnB7cdMQTTqwyc45nevAespA8s2NEp
STPvEAHLKBgLpH60/0Ga+q98UUWY66rod7a9OdXuB9X5t9F1tvjwecMhXCHTtUsJefbSPlHi6Cvn
rA2qzCV4SnehauLUhK4oU+v2ZJ/YAD9qyjapQFJ1eFYqd0TYwP5ZGi5+c+vzvOtBFMJQ3+r60Mqg
0E7VeatQSBrSIq09F0aszrWUTiffJQghksgksIWVbiw4Yed707utxwM10e5YncGMTsawmOziY7cW
nMUvB0fPOAss2KEOtAbVtHRRX/XsCBEUAzm8MK94DpbheplDNZVluCduRMw9XY0S+aVU5NOL3vt7
ChvehwiaBwXeEoDKuzFaEcp0temWBMfIVLIri4yuYJ/eoD/V7KDSr6BgpU9qfUUV38d5rf6520t+
ZXDMQbAKFsgYL+zvwgqCe6z/PnW5NDQBCIzjzm82xwLo7brGaQ3q7hCHdMFhfq0La0YI3CF2tgVY
PaAofHYi/uvkvhrH/YHEzQkUUzw9EKLOoItNWeBEslSsAuKKc3Mw6gJA+0smNFSJVWqMBVyqoPS/
s4RHgH1dRQwdY63KLPsnqqzjhqaov5WoCUagJ56w20LyqmNFIYPXjwzgkkJ5qMt8cjUJPoO9EGGL
6ldia2LNWpy0zdguXdjJwLCAO/njeKbTJBzdb1DFNA/GsV40Vbo0viweJ3r1tBVJsykVHk0DBgc+
PtADSaMNmZ2VYhEeDCXGT/oFJZhZXkWawk4Z/XoMqVRoN01W6jsmWxgHea/fnkQ5a+hacGz53vfj
FpgWINeHq9jnt1099tHd2/SBeX2P0nS/Kka3k7S1sc1cmv5h9TuD7sqCEsoqOjImCdFnuAd1W39E
GEIe93ZHsx68wczl+WmLV9G0hMW7QSaJ6aZSQzewLzfBNbU9+KQQNkBIyqUR7BTLg0XkqOkY2H1o
Z5swYK1F3lkIBJ8EURNpjdzw2s2SMMKBXPWdraVIiAyDWg5eCawK7+BcIctPXMDTXih2k8paJoMn
e7Bnq7D/YDKtUOjx95MwjvfAcXzcuDHzxIdLLs/2wSVfM7PUaAbRhYC2GdXtxUgEVPVBdLUySEqq
+igJUK/Nnt/buJjPUCyuU7spnqtYuD/tjWMMCeqYzpxzS28BEbmIbouimXlpbtjnzxiaoNT1Misy
J4zCkgNXboEDAoTTb51ap++JjocvdX/R9gG5LzCMRWsiCUrdseULANtx4UTSstqKyI4T+C2ubfKc
NZyHCCm718uX1C4DXcWE/GdcMUsW/TSl7sGev5VmEdjE275uGg2NII3rjukGjLtjdjVwSJPNvJN3
gs1GKLq+5VCTjj9Uo66p1LNtzTBBByyr4awnKo8QfSF4eqs/GzXFLks8A/tqEfpsDXLynaxkdu+3
WkVXvnQvkHUXE7uxPzMW71X/tJ2+0JiJVIZ1tCxgbk/VAAwCp/791gp1VjCCATwKoT3ufKGGsoFR
5uXGfvutHeCd1LFar6QeVrI4zV1plD20Wz2rmblw9Ks+GAwiueb5zoxbTM2VJ6PehHyk79uIvj0I
RTVEJ4drmS6CvlIGWVhiWr0fzYZ5CwOX0wNeM7e83xjrfTak3q4BnFD83MYulni1hHczUgPaCPVT
MFthNhs44G9+A7HSCeDj5XF+yUH830oYdKTDps4MbcvVFo/N1kx0ysiGCEaJ66KjWysHxbcBDrn2
MiZz1tMH3ud61tKbvcuN2O4cACeo4qmadk8KEeeGNrUr4b+IkW/KDXX4MbRVfzTl1sOhHHpWSl9o
xb992Z91RvFI3GMq4CrdW6shfP8ikpmrZwMmnKRKJsSeuthRRUpR4M4JB3vj0zyHm/mtS6YIWjPU
sTdkqYqQfoQVq1yN/5d7qI+v5J9nWCS9Nbm3fqZLigfPNpnn7XrwnsVlYDKt9tNIw7W1zhZ2WXtu
Vy+WFC6ZQLlj82xZd6oi9vXHHkzF8PfhMcfbFiJFCBhf7sHtYQaCwMt/D92aMWy0xldceEylz6w+
Y6W6sUC0dVRvc//wjyEU4WmdcMbgpJkPdRc+eHdv8zuY01GqEky0tSJfsIWBr7sjMQnRSnvMAZKD
IuJ2GdqO8TOeGs3SiSJtz6YhcqePDOYHtz0kTSxAwZ4NMw3O9z2bngp/es3+XvrxYJOQFTyiMLeT
AJoz61E+09BDZHo/RrnN4lqQI5L4tPKO0yEi1GSTZFentizffH1ayLgo6bPCf8CrV0yhUR031KYJ
b54lsAYHCOsSZrOO8RZf9KKY+6z4tb4uwDS1vc8oyovKGux7lFNxOQJyal88h+znBfTDGWlA6E+y
q+bfyKcv8GzKKO/3anTNi1empcowfxbGxZjhAocEWrZ7UcnwM0maGKOOe+MHIwtXVkDD2rvwCpOl
5ExbCEfnfJcC97eM3JtA2FccH820CshyKKXkzeFMdO2FqFCyzJG0OMuk2prNoQSS5XpJzbi3ZqsA
BuCzGX5EIEpAxQVCkN27vGIW7Y5ihSJERoQI3UBg83QZXOwA+HbgNUmVd+jEitMHLy5i6WoVnpZ6
WqfaEg8FJ+z8S+y39vucf/HYL4B1Kot8MQSH1nMuKwdz+0FJ1TuZq25hFmLJGoxeXKB37mRSGzpO
cPhW8wfRcGDC+jtrrxzIOJBOD6Xr51iwB5XjGZgpp/rmYNC6cno2i7KJFvxhOWuIWYFsHYKX0kz5
cVX58Xlg/g0+Wzx3WbJozASe5GB/VUPnoLLffTB4JxZgcosZ2A48f74edUhBwcAQvD8t1WuJY9YW
qMDOtJxV3QrBPrjwvdmZdMcshA0269t0F7sMT+BoMxzvba1qPHRxCR6JTQwuG4+uaUOy1WKve5be
XoQEGJPiMIiCEJMmFMpd4YztaJVjco67oCYWVYboQ3Pz3KGEQA0u9vFeyNauZ0oKfRZqsIYxKAat
LuEdzgxcHTkGPLeETlXS3750ZWoZWtZ3E1EXVwCZolG7QuYMdKG187onLU1D3e1a/Wv33T5bYLVJ
ltyiMEwQG3LjyXmZsfOvHO0vAIixT9tqPSk4Iytwehz40Li0BXDunHdKJ4BY7n4J3DTe9Ts9W9Jy
Img1MRlQQa1foJN4mJPWJp2JsiN0JH3m5KRhF2nWBDUdGOL1iHUNbB8lx+ZhqANOUQV8CnUIzQwP
LZY9sN8TKoqquo8f4flHzCvxiP8X4R6VKqCt7Hob94+Ki0I0VnNj17ZYIvdD455lchkSInfdy3K4
oymgmUSP3qZbpsgMz1fdFB8N3mTXkALonTH6OOiEIpYt3xGAQkted9+63jU5+3KIEubz/qpnTPsS
jlocZY4rvOn0+fN9iEAdB7dvejM3e5K2/E9h4YX1FfG+Dc9JJD3ONSX6dGtWDz0AlabjH6MP7d5i
U0JhYBOs2RoNRR8Mause8XPanP8LKL6EuQyY8WkdG4VOjV3/CNWRHSvx7HPm8pr/zn3yd0qXF6Ia
Ni7HJPBKJxZHMzOjqlfrfsBUzPbybqIm+IL1pT6GffdRkHVXGNUq7x7jPd+NSiBho+Fofs4V4XKm
v5ilI0m9/qeKNtXc0k+/CeHYNF5FJoLKn1afiYfRDyf6SKkYkb5dyIhGf0QvD7mp1Un7KQTg+olL
pdmYxonkx7QwnGjQfw7ibNBsSelfbWrnlakgeSQgl/WFHjoAIwDYyD7bPnU6dXo6l3m1gb6yXPx3
LFUNgJNmfAGWYSmPl9VjcIFA29K5VcAsbIMQI1lDPOmxf9ZBjyHroy4kUhwmjT5+35nkky96dRCS
w2XC0LMsoGQromN1HvCS44Ob/Hbt45ydgnPOiWsrNd2Ktf9vcTU2IZDEl6fwC/Ovr6zPr4IJ14fd
EC+6It0TwfFv6ZV+kldsJEkUNMcO5F7jnpDdaRAHXGQXKzi1aQ8VBZYFSHqFCAHHjzHp0OIJnDZ8
fyKnnZrT4f1Lwnn+BKS+/pSGVgguPx/hiK1tEjn1GZAgqdXXVEETbybSwmiSseMzzLYyNm2RJOrK
n8FyaHDr7zL/fNvIZp8UhJl8Vtb6SMRsYyO/2izD59WVE2iVtcVwmupc2O2ootldleeva2HYPMIu
K/6JZOsRQPXez5/KQllj5HLUPKW4w3Jp+NN8bM7PoMaZOpn7S8rhbe9g2hQVSbipXN3RWljURscT
EBoQ6lX9fDpjhR2b15W8IZhiFWYa5PP7LgafzN4TWan7JPsf67CZljxbvxhg2TFaC77sEZy+cfFb
cLzmW2VMUzGlBS9vxa183pe9Kiqx9KcnUW6iWDus8QlyfhWCaoDMpzclEsWFUTip80/q7zKc/QVt
5eH1k0BcT9AvNyEh/n/hpULvfZEHlW4p/7QZcj6qkY/JNDyV/GH5Anjc0w37arwxYaFH6nAyDkwf
Wjww1vXzVPFGF8WrT9t2uTWe0TUOLbb7540Kf/NklZWtOehuiRZT70cBF0BoodUgSm9Y11xeLrzr
eUdQzDgXMdCuUmzyxu2yTABhV0UQmuyIiHgwxCeU6z9GulcR5XsS0wq7GhFxNfSOMV6enJdvpRB3
QCwgKGC7hbIfIkAoIg+bBn6HG2djdP1gZy4/BcjYzX6F6IUM7fMQ08LRyLqDJyNpA/lkuaLbvXVk
eSac3/R6H39TFyAgA122ZPzlIh+1ez0io3fOLcOX+ylJmCKAxGHicgWztwuaQyooY5sXEIL3EmBD
kcMjJf5DduepL0H+lG1aNdHpGJWucve7jGvb/FaLogCPKV2GxfzJO6E8CREDJ5o0P948M+vSHqIF
3IGBp9mN8RGok77IabO4BuUSvUC4oDFVIP89CBlv52L2Hbl24Lqd8n4rBgmyPwMhyZfFZ//qgZ3Q
rxAu9TEvGl8W2GjX3X/SNZxoZM6V+1eaZfYmoQwLZufnBjTlSq/xIeflYmRXEYIpMxNV40mSdVkT
WfrD8eanMNX5gCNFPfSXuDi1jy280hZnZSMTQ1RBkoLEsiAl+88TzgqmRBWB9X2HKiGqNzjYtsZP
sIdRENyWN5hijsiXiN9csDf9dtbkjvIZzLzCHT5EMWh9KecTfTNe76m0Io2Wn0NjzKb5/zh4930w
BLg/SbOiHPSafK49hCf+W1nU168+Zulo9TPlGOnGHy7tY/RgcFXh/EnQCcclf0C87wbzrsoslVQI
/5HyJfV3TrwtAS2iIRFQia2dlJkIvG72tnGbTqe/PsOSb+hmJAu6Qmqh5+04qu67BovXW/l29CTw
bp3m2S66av9KYkEFKew4D0QIHqal9Py04JEG4OdoIp9BGbta5/glJuoES9I7VCBt0yJq+2eSOR1b
TPIV5Wa4FeYEsv3mYvB/uBWv2+RB9ss1aL/gkgZ6a30fgn3+Xe+7CtoH8NjpORTzf4nJ7xwtt5RC
1EJ/ieQMvFtdrjYck/DcdsRdZvo8La+HQN8MHmstZ2mTbh7WOB6ZPEmr5r5yknjTirncfk6aFeqr
klqKjf+SDhpmjnJpVXhWSGqe+iFJ3qobYQc69uMo9rCJkEdlGVWrhSAMDq1nRhpwzh1ckFI0GgoV
XMDsJfjkaG/XZER0H9o/imNglilfT+LUaebSKPKqK8b1i3zjxlmKITSntt2Va78UJNLOQ1Sk5Dvw
vg1KgmfhV1Ki/wWblVfUL/uUHM3+SmkOz7yRJ77bDOfNpOYWFh5179iOE9raY95r5yNEr/+a3Yk3
0TaGrM/cd5RMc69c7HuKJhEx9flJ1YCgO2BD30v7efkQWxHfLiBjRvPCn9u3kFHAkp0C7UlOoyLr
lEZFtiNnjc2OE2QuwxU2jb7Lr73i7qbHVFEYk8rT94J8v+kWRpxA260LFhrtcubzCasfGR5ZntLI
Z5xM8v/G3EmC7E+Zi/D349Mj9STQQt4ludse2HREMl0SgzSsdvMEfnLooh12+TUNkKCyC+dFjEOu
nSOjXVQMwSlsRQ+FZHmUL7/91PleTmGs/qr9iiMEfso6HASbJiu8AtyWoxVcZ071XgJ33Ue4yF9z
yzOg9GHdfipx0tKuMhJcx98Z2bGwo85qcJBF4WWeL4n92aNF+vRzYPV5WTGPuUrQHxw1BtKD2Kbm
gOfc4X9lomtU80LOzW4GNEToXKQbO04/mHVKoWAXmPncgIJJaZrR/rraBu+MDebA0MPtrTAd1EmT
QNcstJ1ismGm6GlmKfJTZpxOn3BAhLZfC1FRSTC2G4Z/WHEEjYyN9AcN0flM8atstmYLGXNzP0WV
3y7OAdh5r/yudwVOFP7CwrCaI3XhRK+ovH/d9U+zo0Wt/056HM7vgklK9glM1bzfB1K8DIzOA3NX
GENQm3ThMrXCYWbaaCPFm+VVivO6fOv5f/LD6FrLouUz87fz0dKTCZhqOMjwEOF3l/1k7eXaPUHN
j2/rB5UDpj3kEI9PMb4wAXS54QJSC4B22uCFibokGbWe6Q2hyx3YldqjfmdyNGoUNx/2fDkQ7QeE
dc1OI5ql+N3SvrErISQHuzcyLbiP0UsgIAFmvnu68jml61FgALMVlV6AIP/W2Ot0af6yZnGVLcuw
NMgt1skx3G4uhH66X80BViQGT9RUABWZJQRxZbb01ev1YPNPeL9fT8JU++iFdmldm0GPhRbiMhBk
tM3LGf9yCuEaXY5nYG/6aeuhaFli7A1M1vNwxXec50D6VczTpFVB/8Lbd1eV2obHRaP8nP6//1mB
GSJ/VK+uFzgKgUWQjyROlxsyNCBG/CRN0cPgjeV5rpjsusVEQfg4S8sOkc65lxwP3B6/QWxHAkvx
eZ1CzneU7hmkzpLZpETz0qwvrW5VI8c/W1rYFS18yyMwFX1yWhmSa323PMhceQx60mpoESluTZwP
1DkM/dVmlvAtc4M1XLI8pnpvD2xEDQqtO5LsuR6EwIupUDgmOUDUcbIdDY04u32rG+RTt2r1RhlH
iZWUmcnpUGqGqVmk5leQS17BfAPb/boUszAtU0W/o5wUwrjhoeCKZvGhRQsw3IzMDwmKRHI/qqWX
1Y0g+tnWeZffBcIiZIlGEf/7LSIktXUqZiJoulUQnlhkUcXFrLaAS5/nnksmIO6SnjSKTPQ7r6Sa
f5B18SaO0rt7K4xYjtdpeLQwTKpNE6tYpHnL+HycPF02ZzWDNAjAuRy4BajGi96PXLA0UGLvmgZm
G84HHVtQZOQbfClC+pQ6uW+H3qz0cUZKV/flTNv5m4jaYNIQOqhGshsZSlz+GoBKV2sdNrZNJp2b
FABMghuSq+mYBKWuKmGR9BY4obcsiSpG4u74BmSG3Qtl3fIfR6vWO058ouvwSFwPZZbbD7YD0fDo
N+778eiVLFaVAE/X8WULd9SViSCFyyletUPVtE4wgDup3UvyJpUKNy0JAL783a2HEqPVpDawYrQP
lOcPOz+XNmxYO/gKwaef65NhTZtSl1Hd6iySomBEqiCo8pu5di8ee/fg+pEBCEUqf49qx5/F2dcE
icapRX+sItrKp3TXQk7/z/ciZNWeIiGtX5piWpwDFbIpsWyAFEpCNFK3oFYy6M/UFBLZtwcyhS9a
iWFM/6P2eWQ0V3TzfPfCCSs9SOSbD2ZE4HH8sdklNmnhKUkfkQBhNIcjVwb2mfi/DnKCR6YkLSlC
A41Hte758T5n2dO3hSabXH4D0C79VEdZy4FaDdtYL2gaaL2UB38dlKX6cBPjPZdZgEs7J9QFyK1d
sitRVKNpUK9gbhEzxjtUF9Dl9oAPG5EAXuIQjJCy2CHa+Xr0+wEdEfifdIhCO9xwuP0uDqibaXtx
fbIpCccTERuFr3O/KjqGS4KESTreoKk9OT5fIJRQ4EnqQ7ERvYPnQbJan4Gq7VVG5rLT3wapOYAU
t2divq2dLQtDnISquuUJQNSIk7d49xes76aYQb8vrOGTJfP/FoXC1ba8W5LDebaEVpBzLJtNj+9n
bPM+GlJ274O21vrdTrbK1xGvGE0REFn6PfV3UDsih7ErS3rZ947wxkBdt+ZNJslTpc9BsUbXavJo
IHE0WZvFz0ZC0AKAnyZSKx2W4M0sXsd+idzFG3ZxPqdFT4UrTvxP83wTUsiYVzYNo5HwhSMkrz1j
c6pb2iOZn5BfMs5+YMACy1YdrRsqLUgt4luM1KNaMAmqjcrkA7ib5Sfee+nPZyZIxntPel0FYR22
hlkJ/CVILPQC7iq0bxr4Sp9/W9X8h0bNG2fO1hWxU8wx3/Z7IEhUDAgB4Ta6L/XkSxoSTNNbZ7F0
PP9m0v/bNQn8QgBetPNnyoOzgUsIWT3wQbPF7Zk/vmchRvroyQyBtDkogZdo0zKTLI25vCJgPerP
eH1zlx1qPxhTkkjVu8w+nSGpujfXF+LrFwLFjRcQizZVU1eRMZwh7t/l46FEcRNX8NvpKBOgdvZv
E/0zqqtAdj5YcSWkd9WUvgyNSAI1bB0c+ZUKS6yHsvUBkHSfF0DhkrzvP/whotKfPwdbsPSeb/N6
KuE64SYV72AqcU+ATZtjhoCILdUGsk9dWFMaFiCs1ktOb0FysT1ln163XiGzy/+hpi1Dzb5AQl10
Kv1EzbLhSlCz0n8I1K4jMnAmesZs6xb0PsLxGaIPcQpsloNw/D3D03MEKHN8zqANZRW7URalf6uD
lTPnYubtrkgtQbAg/r+6qFIknL/g1bcBqYEB7pQG3pM1BRetN5uUve52SPhKUaxxSxdgYM2SEcrJ
h2UfF3ma70GDexV4OC46WKpeAx1e5W3lSFKP4BxZ5jApMzeRpnSBzYzVVNuzVcVUYKOi0UnQx2Fm
Umgt5FLHuX5q5jEuxlBuVWuxiqCfcwYwDHFSQa1N3Ar3HyEZsfD+ml9g+AUQHS+jOR1w+uBi7pNb
uplScdcHC0VYgC0u4Yg9Hg+zZiqo0GjOxjAGzGxddbd/ammDsBQCx11x2OBRurEutWxRopNRv9z3
4YwHDD67EIJfiZiyIoQzeoC713hfs5+TN+ClBZWcIEIq/dgI3dWHLiiG7cCoP5xYCAE5K53dPcPZ
cJAKFsE2sI+KYVync5X4TFMEsi8EhAo+OxpOvmqNCIQ0sYh0pqT3i+i30d0UoxBsasNur5H4PYEr
tNji66bt1U/G/PLoVmQX5VnOzyB1Z05QLDZFPlQ1v/RF2pkcs+LBsgyPVtDFlCQpNB6dSVAwQsRW
ii+/7M0vSeYW8RXLVj6jY2IyP7LZEc2fsEAPcFTQCb+vtjlO+RQAVXGpO8z/j4fFDOK4uxzkky7W
kE7nNG9CmqcTQL0eOrLsmVmfUgtmOd+MFfO0kAwIs8SjLtQhuDzqyGnuZCX2I1ni5g3gBqBR0J05
7PkCjakkHoCL7rErU+1yVEgGuXZlPU2/ciATdEYyY0rKOsMV7dkUBsp2AQC30WDHhXkZITiB2klJ
yqO3r9uvP6oLgSDz4UOzgYlnkiY0glq5P3sdlfU410+5nS/2GzF/akhmcqZrEEmdureDbO7ZljhL
OkYShVQZyxwtxGeZ3gtnvXzpsexkqwN2/5qNap0zgYW0BWKQ09PXRYP43jt5CsJClc90z3ei1uN9
wxuH8Mg/MbiYvddd8ozBw43N5OOnQWRcbT0T4D0ZjBkVQbAP9wI9fNK0bfKSTpoesMLKV500r8eY
QwthdCCJLs16j1x8D2KJw/1u46LvARRYcvKEaiT/d5QoLi6TuOQH6kCPlBnRqnsuKBbzWSpREJMT
ZgwxnpOSc1Z6Ww1ayKzhW662+CWjHlC8WQDjJ0KVrRREcNk0wFHwZB2naqJc/PCAZWRbjlCZueOJ
NxznvFalugOeR4ZeXC+rH3LhgjqXXaUygvkbXWE5CNVD370j/dAzVuRcFsTE5OmSxvLRq7FvJgKa
ny1D4jml1tew22qv2KQNwAJ51AfeL89R5RmvX4JKRi3qlXaOZyF4uwB82cCHe0FhW0qQ8dCOJj+U
13D4fYbWLot/TBu+aLQzr7xw2VV5OsMBaib31qaq5Xlpt+mGSkbQzcaHxgaJnr2DS4S6tvFowL7E
J719oCCbXUPVbpIxIbMj9x9Q/AJ5jbOtsm+aUBdiEtjXntOwvkt59bYHVL4KSIirySQ15BL7U9qb
K9vph01GEvuZwBkEJFMl17CEvSEyVy3SgT+0/tISYwmDq44R/ZHIEgdsnxjuxhCCcvGg/INeC2al
k5aB+jd1E4ulIMYuIZ+heqzbtO4u8ejeRVKMInVjik1O8RQ8iCz3iXt/nyVFbpEeqc82eN9ffVWu
JOs0vPh0huwB96I3I/CNKSfBrOr6+uPuw1fccjTgZbs4pC86ycRzXr2prU87uEjAYdPEGFMcogor
P1Q+qivTPx4zjoAExxZESi7KISWAmSG2TMcGkcZnC53+3qTBOotD8XimrCyf8Vx2Aif7C8OJ0hIb
e18QyM2jS0ARHlLUsiLyUFFFf3R84W9yv760l7hMnVqAAWcLUJIoB/AybaMTJM1zuCAycSnD2ZDV
Rw+XsrcXGtUmKngY/teQAaBZn+XcCH0NIHC2GiBByIPX5yW1wUM6XnhmJF1i8WYkJbZ3ZvkLUmju
utRXoXcE0nJcyyHSd/lRvpNtUXBnYMwuLRxyeBhpksos0othgWGFOhpQYND/V+sRif4Mxn62/dZB
8VKBR75V5UYJkUJMQZ4ajsniCgFnGlzqYWDp0sKuWohGUt+3vRaNL3NLSqG9wRF+qGovXN/KyTU+
AvQ9Hozo+g4sZxsIrJJkNPU/Z6cJsyJgMNQ5ZrVKks0mp5QKI5WZjdPQpXs5Q2U9DaVwjCuF+MoE
iqiJNr6SwqaV8XmP9Dur7RMUbtNJOZRA0hZUikPSrK8fN/Dyd+XAIKsXO0xZvIPp4mSgn3Xkzc+P
WjeSmd6o/Klsnt6XfkCKkSWC48iaAbd0vGqPmekOJqZEza2+cFrPCqEVkZGdcRQZpiMqAlm88hSb
FU20hBx0oPoxiVwVKCiI1yhqKMnqBsNEyUaz7YUOL3pRgdR7uzuWzPHf/SIO14jABPIH3hGVuCuB
qCyuA5TlAJpuWEDoMa/IPX5F0UeVJSpr4Z6eOWqicUtoBDOt82Dxvpj5IBe0Xvoh1s5wxWYY9i/9
XU0jFJLX1IT2P7MTVhlGwCEWj/TjsSI5L9po2N+gO8CYjke2Kby7SjxcbcralgBAam2lSFo86WoH
P1tylQ1EPe708/wOypq3lnBJUrcQplEwl5d2pSpZB0/MNf0MzEIK2KBdvCwS0rcjxXOyp5yJbadX
Z2/6lOThFXzHh7WjKdURDIGNXIkdrFZosZF6ljAaeHJ14Xfp5OCiCfqIZ9unTkmXOzW6j0WENEoh
84VpRulxOD3n+jNHUR6FrGdVu1Xk68srakeFRLwXAfPyj5tdIY8k/VyhWfxC4yLKJVVVBgGJl6Ms
eznFDrY7YyOlMOKgItTkHd+N8Vz2WH+p27Zevg57k6HS5U0gf10UL9BodKCr9mmT9u58/gPYbMEB
jRWY2fVSKpPr4WBRsSp1IBUJhr3ZLOWZlUjlWv1metbrjfPYG5rgFGPgAxy4a6Xuv820TfFl8d//
VBfAN+DxM8wwIvnT0VwTf+gCUVPcLieQMaO/eX8/UFjiiDh0MK9fj1JV0eyiwxL2NEWtyDv68FIo
MrVcB0Fn0IdgjznwvSMfxKh7SwwUDbwDh24hlVkRsx+P91R2BVlCq6S9JRHr+ZKtkUcW0XCdQxSN
DgWo4zQHuTaEQlyEipab6O8n8/8YkMYj4KBPlEGJkJ/f6KA5bSnzq1RX0NOQSw3NPMh3zLQXOue7
F47xNdIxEySsplKmBh+1VmRu8tGaWOnffEne0tc6LlB8fqnSdeqHwLwCJW8s+PJH4ZRYm3mkCT9B
lsZAdLnCnngEFr+yZlzwmRMJSOE0FKu1oVyZ8M+epR9GqifKPa8KL6sQjgP3+D8dzeRMR4rkt1kB
4Ft6KcyhPOtAddAIOJL++qOWYkyxzblmcWtc9DpNXcjWR7yPquWy9FwUk9s22b7zH4K6ECcZmC/5
UNsUuVfRTVYiHqSZ0BnmpOe+ni81e3vG/MVuiBGSJPaWQ/CKQGRmpVgXDT7aN+URyT46HdOLtSSH
5AC63FjSs2APqmJQckO78lOR63tfqvC9fV6rIjJdcskVLpG0dN5wd3dvNOnNH2WJgrQCi1f9kHoI
r5fl+unWHHwM2aAgIJQNjRfHb8dY4Nugn/dqgsaXt7W3WUX+HhWliaQoca4AoFbyNBr8u2qo8VxA
icrWvzU2BA1CLWSjO7b7WohDhtmG9+1YM6Bg7/JGL7kp+35xCR9qF9asI9/gOsoibl4cQRPbem2X
sTt8CI5SS+ybc0wJehqHYTGUEgjeiTlFNJ07ngKpcohfA1OZ7fTKMrbaBRMe7V67Zl5Ol4kPonRZ
WAaK1TlvPHh0IaBNBFoEgvFfa2c9/yezxjS4Qw92bA/EsA2SRR3s/z1FYY+V5SJBDmTB/9zNz6XV
W2sc/XKjPbw8RKX5cybsivFpyxCVE/QGliaBzFNKBVPizlLV1ysn5Tx7LrybjsQTiA+ug63c5qCW
x4cuwgdAkcT0EwJObEjn6dXjXCswSZ4qHNnV2dBhZ9iveTbvTTXzwELwSUWY8P1XikvlryLFmCvW
0zQ5V11oY60AAfGfOTvrcRCvyxXKQCIZIuPG+pWJffpDbiRmLEtcm1gDa6vJdk4Ic5UeTLdRORmq
jfqjYKiFgHLig4SjNgSniUiBNgjqYX+7HTziraMgL1E8Sin+0YE2T4Lh2rdc/cCvHDv4qGk7vSjm
cugt3M23cNG3OMF0FVS7eZShnK3xwPoB2gcGhDGT8mP/5O5DG+akfHDX32jeC6Ijl/0PKZ6MtyEY
Trt+xlIVKZFqAZYSO3GMs4k2nIJo341ZxBJzvWb+YZbQh2DM56StdTpHv4cHw+OpDJmYcXZ/nLKF
UoM/IH+sVKYp27/gHRShu5G7JpvOEfsI2qtnlQee7ns3000NgBzTiO4BwXhicwoXeuR6QPABst21
suQd0+MyX8Mb12li7ZaX9LQq/XFIpCoapaV3EKngzVRR+0X0XbKomKnkJlnx3YHEx3wcSEE847X8
qoJLztx//47DDp0UXXO2K4GiztRT0gSrPhs8EZ46FdUnrKepZetQ6WsG2d4RSYVG9C7vnjqUVKMs
f8MMV4fYFXWlgVJ43YcNnc8lFQf/g++bdopobzJLoxFuxlzCerSUESslinkMe+xlRdQ7ON4Zzv1W
xC8vOHGJ3h0AdyKsbEvs4xKKfWVo4UD7GBxtA7J9NOx0h84g6xKJ2kUl13I4X5y9l/pyVB52lBZe
6n3SaXsr5Q2wxiHlLCguVkA3GmHSqvh4V5tW0lVeDUGZIGE4tzFcOlzzW0sIenQOy5MM/Vh08+r7
DKuyrzyhgFIQtWk7Qbk0pCe3Zq52ydj/jj3rstgAnpjG+FeZXoQt7v0tSplBcFxkENhSahrrm/Ut
FzoqDBovDJG7Sy4q8q7h2Posh0xJLyMOsG4DrOPvtEc1Nvvpt6VUHE59gSl77xemuZWbBGz6ucyW
j/Au/HBZw8S6/crS1KNV8KmcNGvH6R4o4bqyE+qCSDrJx/8IZQGkw4i9koFmeFeMXsiJ06tYRn8Q
Mtgb02cbxZQRd6W+pQcbbSUX31SJpV6mt92yKC5Z0cMzoOzdGUwE5pn4PWCheb8xogCMqs1U1ncX
ilSYaKG3jd+7FiLujCb72NqV7cFr7hUGlqiw9A6Pa+O7jTbl3AI4i0Fa3gfQcQ7sduEHGukMFxvv
OtPUmJeo6k348D0sbPa+6Txxym5H6mA7d9/fog35gIQiV/7K59x1bOzgusVAgs/zeA9PzURr1nw1
0d/MqFkTeprmyZhPhDP1hRvZ8NwHsPyOh6qBd64m3fsQKWes6DAoTFF+gSM8F1BP9dBsIk6SCeBI
LDd6U925yvGDaw1z2F7R5VZLxBseLgZSnbPmaldxNGkQYMB84FLAE43yaLFCP1vGbOR3oj4+wQJB
bsGQamg3duHgBUOWFwX+igXJFwz8L6s0QG8hUp7+FzN2nTuwEZvQWEfQ342up4ddnp/8LKU33GBB
KCgq9riaxDemB9jT9AwhjbdSm1QKtse6HEbxANGXYn4eps1oooDuvT9M3+PHUm8FWR1gYed4saDl
gBtiYOX/ZDx3dCZxbUCq15aL1onKNjEpWmZiLNpNWv50iaVD1w7j8UG0yomibeJkFchJ8KIUeu0u
9/xWMm3PFSlOdwgMdUTV7Ag41QRsbMFlkOeSRtupgEJ4RpdhchJcFuehroYweLaRJkaM/uCiaZTd
Qr4Hsxj3MtHYsWGntad1TBpfGUQRTLd93B9DV0gsChthqzTZ7QDz3HZeMoH0YBBT+vQBsREiUIVp
OHlU9+kIEWkhvaHhTpbbTOsTmw9Nan+Np9fd8eiNoCbym19g6oo1+eEVcoLFUnr3IQQrcZhRayKP
VgBjDPdl7pz+t/3PI+lLaLwMKXyxHBtaro3gmGsA7cLzC8ykCcxUhR0Bg31M2spAekeWnGuWkATh
5V398FURY6z9REqaOJj3043nMak1WOInfD+YIKCFXBt8spbJq/FnD3t+5YgdeYtpoaT/8JEofJW1
DguwEi395Vl3ENEuwB01x2OhV7wDnB8rQAIbNT4hFg5Huiy4DyU6qnIJYef16J50x0Pwjyvt6Ss0
9rRRkErIcQqGGw5+LW/ZeUSd5WtuaKuihot9pW1W4VRDAyTpIeXfSG2PXmKqYsgnlwhWpP5xcRqo
Zb6Z/e/PRvjt06uvtHn0gBWRCYtIce0M0KZpNgdwefvm0wTTUjaSn56NLQBOfdyUZyCsC6VoQPpC
d4fCkgPMv4g/YHV2l+E9MYNggE7OaKvFaPuULcOVYd+JwrQaezrWCrVzcFuHvSD5cX36Ya6CLUko
MFXfRyhwn58oGqnTnz1TAAiFeiAiK4GOgaIrRzg54JWLM8jlJYe7BT7TssUeqiAvsVZbAmJfNVQN
if5J95CBiFx7+VGxKrhPaELkNMB493vpMhHnyHccMxaqrItvGUa4xoh6gXPMkNE0J0F6FCkgM2mv
xsXPl5Le1HqGUmWo2pWAhgmmzSu0uYnp7PknMmoNgjPsO2g0zDjgs1XQ7iT6bimGolyqETJC1t8a
j3nu7hVCg2jVB8/OY0RXElSLrxD0ln+7L36UhHCVWvE2JPL4B/Le2zef1CrUmsjnoGoJuCVwAE1O
NCRJMHSNM8NVQVaFz+fu0OeaoEPt+unceAsxwQtY6XsIm5tePirQfiaBMmwOew9s0QiIE3cixO7N
pHqTzwBnVbSJE+oFDeB4aCsAuV4DR77lrrbmlOUhF++5tYlMWK5ElR3PuKbrpFKSvIf/DJT1mo1Q
lhhIsUFmC9nU9mbnK6+ZRop0lQ/UJ01lVWXTBWic1XDcA/vRAyXfjNkwspHEwkd8AxddcsAhbcjZ
r1HplWFGmgyHEr55P4D6fr5DkWcwRzYMTU83CW96mdfrWnzZPnppuZTuqeDIm9xim3iLqKpreSDR
id5uYJf9xcszxp4nevNWhLqjOIWul/dnIwHMySrh934GZOOYq6fBJ4dWEzNCeB6wrsK4GbGUawlA
oQzqoShUZOSjaPPmzqaPInib0wPBgKNtK+RJ2EyaDwZPhyoP4HidTMr9jL5p2UqwLWd5G7ZHq/UP
Y6b524PtwURllBBZT5/xR9Guw8XoxmS+cCpYeqbbxiED7aoC6lmYkBQdToGwbtQu2YrPAwGs2nKe
OIz5f7ZhmeAxyT+T+27MS4AjypQTHKAxOQpgvbVWs1QDTawpdwsKMSBZNfJ7N3B6ak9lzQmhB4uX
ssBqMu1aX+3qPkumrLntHhkRHevvsQb0k30u4hEzvOBPyPsJKu8K66yAz/LFLA6GQZJxwBUGRQ8l
IoOD+ObyRGXuqxZ5YhkDLxQaHQeciNhtpHCz/Jeb0iY82AGlAuiKSvsfnCzejD21VQiCbsqZkUPV
YiqnPquCth0XNKZTvATc04NYTUoUsXrUo5HrDGOq46I67gCKkIU/DtQZNvkVO6s2AG7ffsRSJ8vR
nNXA2FUK+HuQdHO+w6+S0qu8JC7Dtfzehc+qU0a+MsFrw0RGY4V5TtDKVz2z3oAu6xd+NhNH3PPp
dpTjHB7ZyKKiSdOvTC3n5GqXcanFlOrFw7e5Q80DYiUZ5hI+qxfopxjTkAWLk1KwNK01Gz+ixV7c
ZnYcBf6lnC1WnYMZxEtMvuE4yJZNpVAcMVDc9DtLApAd4YvxrTfI718/F+iPouIKB81fj1qwWnOR
l0R/R2My1+2l+bhBqcM0kX02Y1tzKtEYLYYcrVKmxe54wGzXGcYkfoafWESldTgIJ9yM9iaXP8NG
oRLHKW7LAzOlV86Pb24GwyEBzW69o4oNEb8DlTTNHxVSB5f/vppW6Ws++1wWlVyDB8cgblf20bA2
aQ8QynVH/CQEHgEIML2pvBHoM8hYlYCYPxflBk5OkZGN5LfyC/8FoRM5iu/8eLt1sYcyPT1wr0t7
IdtI2DMRNviCTiK5Dre6xZKahCu1nc3Avj+YXPPQ0HIEn22nCM1xYIAkRKMkrriu/rdBalqbjXvk
JgVoISCqsL+5N11xyMJDc/B46MeHRtLpunQNLDeLAyOIuBa0wgxmTv6rcO0kuVz/n5107f/TbsFU
ov13SgI2apdSR1/lOzcPVxmt+j/0bidO9rjO4TVibK0bcduXxYLXYVhzRcATWR6bPpVSvsnHe8TZ
+22UtncQ0Ik9W+1m5ujVdU1LHttaRAcLKs/IVQoabS7t+UphI3Gyf7xk+ATKRxNYZpS+WpyHtPxy
QR+6B5f1vrvUKNENxGmXOivTGATf6xXiK1ocY80TVXhIsgpjcIGe54bV6ukF4MgqHW2oXxXsJwvB
3HHgS6B0HoqaHcS+V0JXM2mO+69T3OmYhytj7SUBEoPxhaEWT7iYvpdGhUhsId6SSI1j1CZGBAxm
+AD3NYd+8J7L0wmXc26m2HSnfusSyuu+dLApXfSBVBOhxyamLawRRXYU8LCLCZnYLDbbQ5H9G2DP
xUTiJ+wqXMuXN+9pCebK9wITZAcqla0xOWlR7N+kCi4qtbW0AOQyLgNA3epQjRbFnpx4I0BzoYzF
46cjPWKuouyL6ZMC+viMePcs9dM5Ch9tnK68dmhn3zbcsrN0nhsgdBD8tO9HCQdxs2UhLSdpAn5Q
v1h95yRMR+dCUOv+qQk5K219cn2cXsujfjmUGUTESGUPd6aXueCzzJBnL+Wp3p5bY4ZyEZzfPbxW
jLxfWFzGARsXakMGkokXgArc5zuh9ljBl26xJ3/ojzrdykj4rjL5a8IwooQlY8C079emzsYLJdV6
JSW4tr1zNdJBvJOFsmWhA21uaZb37BZH3fhkf5Kv4VjE3wk43T+pGvVokADhBc1UDO2m+omNUvQ1
026RqSfyjjhdFlpVpFj8JMRBWw05CkF2PBuRv4bu7oDCHlGq5kQIBH07nV5KiE0IpSfTfSgDae55
iId8n3kMc2/lBxk9UKJxXVZT5PPWCyUi80/2TG8Rb0SoQYECse3punGZnJRM3Dt3Hj6MnpFNCPAu
LnhlBoV8q6+YNr6JaD9slKiMGYrBbPz/yENTocZ7PR+nQ51T9G/AB1Ea6Y9CH4BDelMzKNLxrDA8
FC9iO4AC25QFiw7686iOj3SvAGtvKnx997RD9qUAl2u1FfjtC8kpdSMEDkhuKnpjkVs8MgeCM31j
Qk2MzwHKq2Gj8b/0VdIG6XBVHuaNHDRBKmVnwuEPUfONKecjq58BhvMb7j0gvoOkmG+Gro9Vclli
7WZ/cV8vqduwZrWUAVREt5TC9JszwmnmaBJ+UL33kNJLKg3KXYj7jUb6N6QITMpuH9UFQdzTZqdC
QFjebYBDYqZHEdk1O/sN1f5Rel0XkavFUr9LRuFkW+cR9ZiEBHUDJrYJ53eOZPs02xBHJWbfSoRR
7uShVozgcnRTLQdx8guPbgLHeeEEa0oOuZlWMkhPoP3iHkf1kzUKqieZYKKqn91xdUFMSyTegtXf
1m6e84rmIf6xgytVDBI9DNGvdVX+DNjj20hysAPn6P5bgcSm9biJzC2xw2po3GhDGJuRIeJurycy
ppyEdv+tHTPVkdIwKhg29srb2Egxwd0VBQMERc4eYsoltYv9c369x9TAbXZJv6cIqcskwUYriyZL
Q4XxCNMV4clHTSfUSh8BPhKlv7/Y++1fBmKKlf+FK3y1lrjJeAVspaPvWOAmjZJ7KZlrhJ0edYdM
vsKuZRDqGMg0iVrctiGkL3qlIi94dRUSoP6p3vBN/VnoBJBBtxhT5WmrsoJckTywowfpb5unL7FM
fiWQTXV0NjgFqxTsPuY6H+Wv9pGfYDq9F5AKyuUDJz2WDPkw0KM6tI+EJkk1y+tJqfUlURf0D6Bl
XSmG3U6kvF/gii8DjXj6r4x4SV8aBxfOWkrp4wEwpKfKtp5BaogDSqhgzNvtBOVttzDxDc93pukC
S0UHua6uZ8E8eUp60uidmcrFQpDMaK2tTML2MkCULuQcmoV2ytBf69Wq7wzfRwkzN0am2WFp+F1V
2RQTJj4rUhACzyw7MvYiedSGKZFRaugN2pCxguriyLxJvsVvCw/El8QDJ6LHakX3doUHIJdGQEbt
TDgbEm0RfyXw2sb1xV0dULzwHhMwnJ45do6FPgfVQdWy6bpPIiRfuMhaZNODVDVHOgjnUsmFkAjf
E/VLILfhxhneQDRmwtYf5Z/I4UmlN53liSMMnircr+ykD3YmfDF6ey7OqNHUT0r3kuQqbRgx07Kx
hCegrdyx8nwkgXZM3KoNjozfQQ4zEiUUGR/b5N8yApMR4yo+TsJCRYtE2udlowWaw4xDXePja6HJ
no1QrauHKFFLDtAvZ3RsZiwV7cq5zScg+ZrJJWhnk7RPSHvc6u2XgBfmiep6AbuThjg5vAc9qMT5
AGUKi1GRIjHN3xUf4LwIUd8sgY+eNiW58OBjnGq1TdMBLZrR60tHJO1R9EOOlmAjemfkeY5hXLeG
EijvSQjsMiWGPV2hFyk050g5kv628TxOIpXUBtJTEWOuqdpSrWSUf9OX2IIhQDOTrvIJBI5euu/t
hr2m9HCi++0Js95gVMIDp2xLZ8B9wTmRFuyTfjj80fdqTwaGzzkUYYRJRIda2nBnKyq3r0JLiV84
FX8eapI2RobJuvVaJ9+KD7VXH/NxgU5+nZ0836pFK2Hjttltv62LdNLj6e6/z3tAjNMVu1svgQr/
fOUsqc4n3B8wxiboEPQc5MYM1LMTRxFAjZIJmhOlZ2ce4k3X+0tDJlsp91Bh7LLLCoPO7mZDjkm9
rAI8NmSdzwbKDDqrKiODWUOSlfBJtSb7fYVnecGkiYA28O+AxeSbzLBbhSOrI3+DHJp6E2VATFac
UKy6nTRSx4UuguPEe02BMSOn/XqVLSj11xfGnDnlSbp0L5brG2pklAxrLKLHYw76JpkZJcK45xyQ
vLi98RxHLAcFX9nK6JTXjNj+UI0g110/Wq0hfZwR/cy9566QLIJxpxa3frcmRkxOYK+agJOKcF7V
5hxSs17rcLeYG2QWsTUiCb0oYDpZ+EFTz+GdJsciHh5glBwnTR/cMh2OMY87XIwuyJgdCzu0Oeqd
gPWJTy974BOaCfiXedRthtNvvPZo7L1RaB5FveGKg3GVHlnLJdgXDaKVEMMlv4LOb/zIpWszE7Dq
N5bOkxxICeQ6mgnIyYDTMgKoQ4/Px2INHyctOJWjCPoGjOG8+WQNRNd5uOKMKdlkbUGQ3hC4aHdP
lkjll7qxKwt86R9QXBzaraUxHbhQ0EdOOynwahdfsMFz49c3liUEOHK1YK8weRAngmTAQqFq/68G
O/n36qFQ3rVXFFFosgbfhneYVkJRhPv+N7uA6NMWLlFVn30ZuoL7rQGJ/KUsEqu017J/T8nFWZX2
7RlYiLje7ayPGBrM+L8vkWtUzjgMj5Rj0RbVBB3BBi5/c21SMYn42lmDCwM/7lT/to6k0YfRazu8
F75zD0FFAFtApqLiFUJoQ+oIfgbeFzvTxdRDM0NfJacqXEhVD6M+N7uJ44Sw772vz1bDEto+yuui
+OwJkfoShsNiJJWYVHtUIOztiyQwZStdMttR3yWCO44JE16udhrcK8+t44hjXm9lnIK0nd1KiM04
Q4UcsUZEARDgrLe0quN0/BipD4/vdNToiQpxrB7Wi/uvhygS77XwI6+po+vfY5ypQi+fDdFBiWdC
JdibUKwHLFCopjuOWGS40ffzukLTy07acZDIZpstwR2CcLXOND2ckveelPGcE/8UKiSiJuzzTA2Y
EraXWlavZFAULnaM9xyObW+jb08PZ6H4X4cWcVdHA174SMJOF4pQmt+NyxLywJ3fp6bvsakTptYk
M8RieiVsY3quTiOeujC7awiHynMNz466UCu9pQzn6z+a7ZuMJS+kNftwXvSob1ZueGBTdfvJiWeo
xY6RKM1Ke5pjF6FP0y2BeTsVwz8m/dyZGVWvLBxdBHRDrDrkUX7AL6qFvVaKdCFkD4zuqKRcEAn+
dktpiuFu862B+eXR4OyGKmyXnTq2bRiVewYWrDrmKJh97bX0wXFTxuANJP+MYxZYSKHz491dJKCE
dGmiH+N+tIv/Zwv3pA48QlcE+Ybc5HiX9KZ8kbp3rOJFBqcWJOeeKPLDx/mD7q+8Bd2gk9EFbPxt
FzDhbbPybFND9UsFvqUTyXhjTWYe5ilDsfQJshhrySgPMYRDVhQDmCXqLowZSal/hkVXTBxFQ8UK
S9TbaF/KY2qWgk+M6YXcX2hTAcasrVmgoIrgevfg0MvHO/CaRf+sGWeHYXmbbmgwDpvIl3wtZfGZ
aAKDov9GBBnVstXrk8Ji2i4p6KlhwvbsagcqzgWi66fzOQiRydJpyq6bKwOay2vExxk2HLdKc77J
qMhq1NfbnjHnUpbjWGni/UK2Q+I9kfa4noSNEVoXye9bx8LzHJWTIENKyhFGn0AgIBMguTwZL/IB
wWr3J8fxGRuPLwyMpc6IvgLuMMeZ5eav2LU+w4WpkKaN/8FhMftLaABNegKmJXV2OFKwKvIaho8Y
TeX/wIIQAxjCVj4LXimjYHx4apPWKIPNQ5nwXzxrU+khkajVa9mDn8EOytnxxLaj4wbzDCiQSwMf
9aaWbhBKe5BPtm53FQQekmCYWVN/FPUdiQS8f48bfBZ7ZYMEmT+7QP3bSYl/4YH3xohsQznZZksl
gjuqVVDeb0He6hihTuPqcZtESWuFv8+TRader8ZH/J6DfFCZKA6QN31xCgPK8MXsJHMDd1In+eQJ
W6ChEj5TdQPZpLEHXjDIHSMav3KkOQ8FJpdaWlLcrwosBg5RnZjUaJWVXydggFMRthqVs/n02uBq
NsuwF4fkG85Xfd7v5q5qlfD4oX45xnzZbwHnsm/2je7XVaGeKcTj0yJ8u/d0cFocw5pBuGXfUJAq
qAORtO9GHuzJHlf8sEXQlZlUu/48S8Hfmq/QdxhYc9xcuQEAGlLQ/VWuxbnpaTT5LhV3gXQ3jDaE
+WPClDMc0AzXCOnbhjuyz0soV9enSE3pWVJYnEZX4+wkPI1pyPEjyBTnTIQaW/a2g0Wpc+Dl8ie1
Boosj4CoC/O7g2NezJFzt+i6o93AzgC0QQ/hVBGuFF33k6dHMT3nXjSxcJ2LrOGEcdjQ168cBu2x
kASyAxRn38rPCpGaAcCur/sl83p5zlogH9Ym+PUAb/m5G77jV6JjO7+9U9n9fdXCoOpR247zV8O7
eZddIBrJWP1ez9KoYIgP7f9oVkwL8jq4gfxREroGv3ED+BTZcLLtEj+0lLIDhlTZAhQqbN0+d9aJ
Jgp7u3cW9PD41EGxrJZ3Ny+Q28k3SlPsOtVh5TtNGmPnOzIU7SeN87GLLKgaRsj4c+E9Ujn3lB2b
Y8BgvIwHM0VonMEvBydm3vmvu0v7RAURRXWEJzfPsfwo8uvegXJNUN0g2vQZV93+6fkSGDxrC2ap
FUXUDz9z4i6tXpzBIKOddOgVD5mIhtheqp0rrvpK8yRnJs3FiHOhh8GhcH0jx//mUmLPTlyH9zb8
DswZA1X5ms3aq0TULXoKPBMcjpRRgCF4y24cpKyAttw6Im+ky2whxtYMEfBIcAlkSUC0ZTuFblx7
R+wjQkX2R7mrufmmEYnduyrgyGQfqsoNFrfPPUFp2w9MBO1BF75Tqq55GcJV13Og3SN+3bx10p+a
ns7q4GCczJEt/svw5rMXMvY/WdnOLwF0El9r6cw77qPFAHjM10FeeNigfjVko5wllbjrzMR5hD3/
HwowpYiZjQQPF3t72P6TBDVqkBxWY6Yh7oGign4PGx1Ogp889ZZ2nheKs9Z5JG8m9cANhgFuxumg
AQe8CtUbAepxz92YT9el26IEI9Gvbk+EDifZKIjfr3o0X2lBirk6Ie2QpEkgND1AYTDlMCTRt3wj
7vh+qgEOjwxtpDvQoUMwX34kxHKOfAowGlN5GdTGxegmehICD4hZR5BU4ULcZLXfiFAyye1zIT/m
ai/fuSnyd83zC5ZLoYGYO8n/qFJxEGeu2rX0Rc6uNWa1ggBFpcj/54G2LGz0gEqxq4qgD9fDsQzG
g5Pr2iQGY0vu8pCIOGV7GueVh1ambgkRuYlC53hgIB/DkOVak28SgM0UiB0jpaPsWLU881tvjagL
hLxnQjRu9/ymoexgSVhNPLmRHlY0006qohJJU04xceWTFgUXyRMv2hr35GIMp4tC9RSUCLEz61sC
c9wPMQHsa4WbNOr/JK1aF3tjw7OFAxCAeRFgN6u5/EcmcsgvigAsWFpFXA7WPo/Ui/yOOJWuiQBY
IM56vKsHmqSA4mhjtke1c2voaxIcilFErm5WXp93nfqLY+tyUyc1qXIy02Q92kXjsV4SJ/y1/LqD
1X8K0VAq7kST1gN7iZzv4UNUJ4Isd5oattzPToHLkYbgake/3+DPA9Ry5Za+oCCihCY5jtnWrBW4
+4Enhtf93JQjmONyhLMDAh9zzMJ18nLEurxswPZrE2/+3GSpKwoRElh06tIbiCs7dnHI9mHjAPAW
Nkm6MmSywikzqKGi6hqjA8iXD1mJcW8UsHtBBAycHXtH3t+Ldh/iRprXtgyh1SaA82q8MYUs09go
U99eoAMm2smd+olqMrFzJg4+TyDykDeSxhUvcBRnjFtlSjU73bzAu7INAWWtTMF8pG/KPHlJ+r0e
f/ZplWYNvtfUXOYnwQ9n+ZblYfFGJVF3elm5y12jlnzeaO4RF8B4ZMWfDcH5ugJVocWIdqKVGEyW
JkCZXB5w+ukrQkhI/5GiUKGjfh/9IjGF0wOIxKb4hCJWTf0RLE1tnKuA6vEPTbPTFH+hbibRKNVC
EtIcYsvukDypolUUzhvFMN/+kLFOkz9C6pYrZ7Dd0USVxR/mwSF7cBftw5p3A9wM4Mt7/wqZHWFz
Ad+qEoznmQOzgOKIyPB1q9zlj8L4Dhrm+9zPTiZhYUG28OqGkLgtGgLWtbmX5plYBvIQEHu9fq6v
IuxclGfXvJ3bXDpkn+X+AoqMSpgogcXoVS4CW2AHSaZk5fp5TJ4zzEv3DnmtHVG0loVZH8+t97KS
rFyOXB1kXqTDHShnZeWSQG9B25R7mEis69U+Ziu5Mletxn23MGp1sogP2PsVBoQ7damYCIBlP+2V
J7VMn+o3E2l4IQuO9eJfspzcvPtIMXWD4dBFB2aBpTSSLRoY9f2LTcIK03/07xcy2lZ6adZq4yxw
z7iZLlOfOGW8ftYPKfVaVda8XihV4D5cauZZh381q1EpqybLRdMb+zk1i7YPJijAlG6XXGphZjg/
fwTAa103r7ubxq2gKNezaA42/m4kWG8mwE4ZcsgbtrX1rNr3loDDD95K5TjGX747gzKyJ7lUZXFV
bBk+uNb0QyVTVLoXWcPGlzMc1KW0w/55w7zUrZTRl+rMHXN9Sp5/340nlBuD0TtKzhn+0qNUxOWH
DWnW8yGYCuvuaIwS3sDe8XYjndHLDZeGlBvqKwfhg+MYQwlvNPC5t1X0Z4F1C9s5cIoVv4Vwy7KM
WsVTVDMGZhhgaNozKLVQ4q2XIsPBzV7104a2ErOtW5O3zrKQxTB92Gg4Uv5qrUSfILPsOfY4ssf7
mxt38GemEPnVn76j/xze63gjkeRDluzJkqkWYs7A+x9Svzk81krC5BXyF3ZPBEOwbpjH/lIfLTEq
Q5l5ch4/de9TQpcTXmt+IGHeytmU+VONmb5JdA3kZ0MaOgpix7StT4JM1Ag7Yg2eSWPS3cuaCJo7
38gQXWlD3Owyd2RaHdQD5UrPHu9Otk+oblADc167jFe9H5PejO323CdY77ykZ8JydHFhdW7D/W1j
75C07kfs29O096wy93jzdxM1eflToILLMjCoKhkYoMlZbWGKxpPwEpTdam+2YFRbNklehY6nNd/Z
2nbivCT6hT9Ddt2qtNptcAdUU/uk/568AAReal/0c8peBfBHz6NgJr2lhyV8G4zu7b0ZyISQWdYz
wdPx71nnHEtamOd5F90WBWvBLV3vuil2x4RSqpfu7xqxGx61X1NrxWQLNocI3AemVQxLvu8glWUb
8tjtKAJ8L3eb2M2aGrDVbYsofxcFjxO5hfTC7FNEiO3gPDgWKeVs0Y2OPMN6/b6grJ66KgK+DWQp
UGW42hRlumAc5+6R6mbnoIuZBsTPBBdeu/tYxiHFtnQQ4W9gyytmLQwhRdvnbvJ0Ozbe5lEBjYON
gvL3J9s4DCoJ8uFBskmKhTGmMYEsm6jyk+7+G0GXlvHiFlym66Ejv1By8vg51hkY/YJ5gvVUyhHH
U/CdjAIFLVDkRpAax+SvxdMdf+ciNaZiaMfKORFz3aa7PanWFP9bHqRJBhWUeuaPsFJJCUxjkstn
xzCzQ8s7FG1R/kYhdHsWnh7m3w8EddSlb4MwpYTPxUzygaOhpIZn2bPnL23WhEHEk+yfLhLqXati
xqGds4LTVQ2rlQp0P4XC99CiXAr8TiPkbzkkJXyFz2NJaCXwa/K8Dy1KudZ7jP6bmD+1RWs4dzwB
0ndd+ulB4nfMdzEJ/eTGWFwZMIicWS7J4tjngEfWE5wXEYGR4yAiRwUzkqyHT3iaagRisdq4ZX4s
2KmhjoBIm5k6tJbYRnGNsvkMwH9Z64gdsO5q46mIdHqrwyt1eiishXuyAPP3SkwNr6tRfyItWR+a
lheUcmxSHmGAgMYJ44rnPesIbRfqi54fX2VX9mjGH5eRBPi8hyCed8n8nwmUG8PXSpTX4xRvtJH5
xyYdXeGhV7fkjex/HfIPcUIPOyTVW6M01jW5iwryE3cFx7n32nG1lD2v8UGpUYSc1zyo7j2oaQUF
sdQmLd/fB5wBWVrkc7sKnn6VBFllJAmXWvD0RGMZYqaZ1cCOn2kahvLIKL6POX3t4cDi8W9CQRZD
/2Y8ic+oIN6sQdzGO3e7BW9y4FSjPkICF+i7ZysQBVZV5nH4i80TylO0zlOioa1N3JZ3pdivennU
bWU9RaciJrJXkF3Qr7MlrFTb258fUrNurFFpee+IWFlPYRvkFZbbhasAOSMmFfTzB+bQCFQFAXzT
0o6TH4vSAVrhGzoU9nuaFaDV+Y5PAepaSceTNvPQGrF93fsX7cNdhHldQCs7yJJNCgVrQYthvm2n
wmSJG9offb1HOg0C+YW0wMSNPgDmLRrrqmJndlIl126ryGBKZw25VcGclhHKZhtz0cpkJaxvcZ6T
Q5lwISX5AakGHFd1nCaeuGoClAy+rqBEGSOYLXABziHr4eoRYzjiL6SLRb4JCt4wYTdMe1WXMaDn
0yDwaRoW0ZK9DhgHshxdpUO2WLR7zp3wAIjxlExUm0TXMBlEgcXCl2eNs+e3K+RF2JJQ/GcbuXwU
Zt7JEgpRUM+k2iIZ3OG6ek4y6E4L4LYkjSiaOi5AywDVQSKxKBoAvZonwjynxltIfxm11by4tXdl
OWEe6ev28HtmGoKnVz/4AZnpEqsaJweMNYb2qSHEXhVV/6ISotCvqfHwMX+vuUm7AEllrhqDPASM
MWzZ1lzkcD+UCNSZWpIMQmPVz1zwthj7wTB0xM1vmyVlMYveXgdiLvfVr/ekKRHIRMwn0LMC90ku
TL5gaFVOi/UAgry0+N2m1kgNlvO2IUu5JYCoc7B+ZKyf7dLylyupK7AS5U9LuqSx0WNBpmR+RcZP
kJ9c1Pc+OPKgm8uOn2ZFCnfq58fUqwnvEhoqUA9/yCZpvqzTFStwx3cVB5KUfrKiAwFe45QLgPjm
+jrxrkVqxcUuF+Gkkm3hYxZKSonkezf2ln9TFxPuYFX3PE2FrEqg5062Cx2cgPsi69pCybEiHc8r
w1zqakqXR3WL3g1/HziCN1/oAMPW586uNY/ZYkM8xyel3bfkVSrn+N1AQIqg+/5+qypvhrT9X5/p
y4UPyr3OGG0HMtko0MLfpFQ7YYnBk8FDFiXZb5BAEgfSQY2fJvXUz/qaKF94Mf3/palEcIwcX0s7
B23hu+eO+ojdG9hiu3VN5h87wLSRnPPu0JoAnaJY+9ByDam/yEbzO2WjfSdeI6rcnIJ3aaZHXzN1
nnCD1/YTE++LyYxTXo9XZ4Dvf1XnumFvSXfxIOaBCBjNoIIfmqAGp+3VB72qaCgl3eBIeFzIzLfq
EjSsFgzcHUmqOSR5sp4bwS6r6rycTlVPaiJ/kJt49ndcfA16DPo61lwwlT/fZQFuASz4vbUz2uak
eIFWDaBvdzZB6StPfnlJkDHY9Ghftj3+aV9X/YvB4LO5C3og16pbWMwxlJcYnMfdTriRouS042UZ
W6O7MhjefUTb0BIVGvXeBTkiXxym2Ah9+7qllY7XcA64i/+DWf9isFjdM43+oGmQOEIyimSk49zI
dggCwxHBR71RNf11h3SkyglQPxKbxHgxnvK+ivBbKQI4xxuVxWarjre6QLYQrb3bssvysblmIRdq
TVtTDPjHrGQA7SvXXT9vduyYC1paoAfjKwaNe61VH2cFK9Ru6pFHhTOXXOba0S9ESQI8W6qu5MTW
aI8Du98H7o0s/v27bmrhGdb9ITH/lTlG/umJZ5DM0/lPrBAR4RQ0oT0Z7ga/aDWjU39hkKWY+upI
zEqWcmTfzUmgmH4NdXwHYe0BErUHLY/JUtYyAHFmGzAw1yNxTxl3vc/fQxGJ38TXoe4GnZH132jk
qSzhl8LeE2rvtxebpbKnRFqDGo0KIB2QQhwwr6VxT5KLr+P/SVF9rJu6HYZ6sGWJ59BLE0KAsxB+
CJXJD5oDUVH2Js4/ldy0F8dkyfELn96nKL0qSYXO6exmCaTIG5CZYjugac6fYZvMe2OGzwBN7nGG
guOQN2/JHoSoygYxCUJ18OJh+14rBLXyT1Wj5A6iMsWhx06A27Vxkh4mOJ7WZo6OQvUTfWoj/Rp5
BvZwbj/3wpjQdkyLG7Zc5D3e03RqhACv/H+3dLLDETPOw7qBM3pvBWbRByUVfH56b44MItv2qqHj
3T8CR02hcenVJfoRUFweB81vq/F7530qHmA61H3eNw16zeRKEPYR3aCuz5f65wiEVDtnoRs9Cnsl
eDPGR8BxhhzPSMWgoydUbtMhry2PzzuucJrHT2xg0ivYoYbxfM0W7tg6RFp96k1CP3B01s3rM3YF
uGoUxI9WkuPKXvdOccJMUxtGgyYqZY0zHwshUdqnYOOZZNwLiEeGF3tJvuMWFGZQ3NwcNM6Bf1wX
edQBmoPv0jl5xoHHk8Lgsu2QBM7iTELrjKDfrSdUOB4bpunigdgMoMEQlgEO9DIwObIabKseG77y
CfUOl53SU3Fcpv1rRr/iGzLN3Kieduj1vnqjQfwCTqJOCeE9bo+EfzgeWKg7rgO/ZhnqfmUsaFzv
k0gP4uzBGbM20hc0ztXy4wP9TUdwpxzFwWkNPE6ZqX/FOlm2AsuGXma2s8GKF3u/wyHJMpBZXxY3
7aufiTggYs4pAWmn6NCvgY8vatGidBL7QDMjCPZ6m/Na4fxYJizctS+dL7Py0bYr2v43bxto+Tqq
azY+ztwIteSiyQ3nkFTZBRKRBu/ffVDb2i1anlQVPMTuNj8kFp85tKPFcy700FyLHQdfJYp1AzCH
qTcELBBAEVcamfwx1xkJQtJA+IIR5CPcMRYTMspoh06yAumhMzsr4hSW5x3gi6efaG7e8z8ssBqy
hya1tkHZSSvKZWEAZMQRMoP7Wl+sWI6y0fGC4ekGzjL1ShIAWO58WbR7uvnZ8ZuRjh3kA/W1ZMbF
C8sKE8LiPwmS5CKROTmOoqjGWLmFqDmbLwAfskslVynIhnTBxmZckvYewiefO0sY3pULVz6uI3Lv
1bjC6HGN0oF/3BVcZDqbHBfDcn687EYfOwyS+8vs5NG4tnlrUDryKrHruGcFzhRDwEnnKmQgWydG
njt8y5vesNQ/9vqt9sctf2dncVhEfH1yTlbXSqQtEFUdBTiRPIv8xDnXnu1lcTu9VUEhdiie3Zzh
smo8HKoDQk/wjoIvZ0famtor+wSvpCm4599LU1QsPcFfZ6eOR9eN1atFlpXbbaO8zN3BUuWcQbn7
FI8geAZOhNxpj8p31KdhC/6cH4DML2wkJGMlflYEEuMKcyoXRQy1UJJppXvrCgs3KoG9jWryibes
WfWVuV6UOvG8z/iVDnOxEAlraFDUBMZAZulGTgB19dOpat5BhNeY3cl9VqGSOsZ6H1B8AU1wa2YL
+EHRHVlsieSoeaQi2WaB2EYABFdAgpso1w1YxJjlF5JV8AeKLw/w/wI4ykHWYiHXQs5rfL1QxT2T
BbKGuCqW8e+nuC6ut5G2Q1WKkbXStjVvWklcyZtavKNA+VjHR3bifUZV+KG9Bzdb5CBHsdK7+1hM
sC/W/A0VXgN1LmotPF+Undt+QitLvS7e/wEJ9Rg4WLCQqmviZ3nXibebtOxTPcU2mxpcl11aOKHz
G4/wrulfdxAyuMcNMQGD0JaWI7dg7Wb/eh2t0kpO4p3m0I/dDYsCyw9WO7hhjubbC1HUSIp4TuUd
mgbHSkCeeTDHZIYVsipEnO4aw5ksFLqPYDGAdRn7kJtd4t0F+m9KvNntNrW40e4eMQFttjntcHMc
EnDMBsp22Yc6dsTw7XKqivEOtW5YSwfl8oE3WAEGaC8mW6aRZTeRO9fag9v4XnltCx7J5hZJK7qu
q2Z0PZ+pjLP1EwO0qIHDV4oYkkbziuJRtRd0WSM8kKenkx0nM3d4rViMaVYpQCshQ32pnnDlhiZ5
v86UXHrqM0m5gMaIKDibTBhPaBvqVJQfBTfREME2HVurukRzkTMEPNPkm7zKq6jsfpo2f+JslRl0
wbZKg0NK1WMgjtWKHD40MiA3Rx6cIolW5YJq67nvplEDCHoMuZR0IG89fb/Q1vb5cbjGH6yRtUMk
tLfS3FyuGzBzv3tfg3zFycZ2fu+eG5L0MjurUed2z9k3/l0wj250MKQ39roK6QfFgXRh2kL5tHiJ
ADywZyRcenFuoXg7rXxUVlLkQUqWUMlh/je4h67ZPxnsACyCIjZiZQ5HCOvK+KlhcMlpZ9v66KmG
mHYzaa+c/csaot3z1XiQzGDf5NBhdZ794kFLoT5ScykBR93hDDxxZnvhBxIjQpDDFm136+Fl7Cm8
izj4FDUQXarNkRFEouxQmPvFxWpeH5kAXbtgUXlKJpOqr7amqSNz4ZWxCYEF6GiXgh6ODG0wj+sJ
rGT/Xn5ok7PcIkyaSTXUztF92eniy7DFDTn0UJYbyP7/5+Em5jFf+wHyln5mOMP/aJFvLI+apOqO
ukauYL6/naplqV1yukHXqX6L/ruS/FAZ362Lj5PRzbeKTUdDgk5h0GissZ1iyfLF9rZzvN21hh2u
ELQdDB18rvNea/qnTnimUurAWymPBaoZquXWCYTHQuc6j9abs79krMdbZRRIcIARuMfndUDpotx+
huA2mTk2hDIEh0VrcGw2OB9lWJ2GVUrUWKKkGvu7cZ9JkoOrtKtJ/QhBUN4/cdc55mQa/Hnhly8s
NSiKP64i3fIuL/nA9gmxtQj9Q7zJ3VMTNL8vPyfZ9T21vU4Gqty4PK/kjGCI65qMn23SYZkrjM/L
dp53rKRdd917pouVbL7yxrIVvUnc2WajM0ZkXMHYCXk6vWbn5KXZmyNDvxjTTwvNZp0qUrEC0goW
zfmy5oawPODg0E8UEH4HA7TU6OCYiq646DBRbK5isVZffDNRAGBXjYNcLxcTjdM/mZhCkOF13sn2
F+gzwfeeQ0aRRfUwDXZv7+LjRAHSIxn+FejgWY0UQBSMQ6/ilzUkSG6jp5gMPPHAJAVgni+duvol
FPUM0e92guUUTDx9yYTxyEbVvNCs3lxAh6h3Q65Ftd6EMabyeOXn1pm+mFj3TLXrmj7vgz0Z4FfF
cjHYecj9SriB9pye0zA2ny3Z169COBdD15x00mnAf6kfFdgLTs/yYlMjT9RaBy8vuRz6ml6zaW93
5NVehnCUEOCtaAicrCfQ9MpLUtAB4B8muIuTtd1Hd2QHtJVqzBSWHsEv8g63XHFSYs7FdVhAsQme
AylqO3u73EnOje1GHGQhhzXPqqui0QSPT4hJDYy1jVAePNmBgEDPqhOQbZGA/u2JxLhNX5bfknrM
mHV9yR/ewBBbIPNny3S1qWwxsMgTjWUXLVSYhdSqi0U8dZgAXsfn0fRj09cMjM668b6h5QJptIAy
QNI2SGOHAjZLXnaEnIng0uVhMsOBm4OiIkRlNl1y8+8cXOdM+/sZdBpjaBfdWhyasQO56Uq3/zU1
A8aJ0UC0dbBIjCrcp8u1L5rAZ82v9SsiZAYZ/P2+SAGDxFX0/5F+byJSv0EexSHHF831468pE2mJ
JXwqve19NqZhsA5g2zSggc7b5RIWGK3SRRiRx/8wXnSsndnmTwfWkXf9rAUWgJKS3uryz8a8m1bD
6G8f3iah64+8BK2wxnWFmbuueyq5KjnTXEreZWl6RKA29kQxM6hPaIifSMEzxRL2sigHjHwmCvTE
k3UDtj58pmPV5vEcTxUAFKuhf2TPlkf0xWCy+nyQs042vjf3eK/U9GwipRh0zLyiUC0Zqn5eh0lg
EWVMBLgl7ylFlFi/gQ4ajH7zpRst60QXzEp6QN0XARiZtSBJshgRVyhfmOPWzoHnxXFSiCnb0R26
Py5Ywu5BNNWYbaaBemKmr+34a0HhhxIiizlZWHzJgzYuh7puQ7y6ipA0Xcl14H4up6vxDf1sECcU
VwpXrtXl5F16EIGY0jWS42gisGpaTuyy6z+AsBcv5NghvGK7nZn3eVPSG9VmjcGpS63rUUjGIs1x
yyDgjoVwxG5eUiqPhMs9i+jSRK23G7K4/+r1/0ib1+grI3C093ehhth0/U/Ul+4Pyn3gtFkeUsPe
z2akBqT5gy+A8+vtFiN5QpqvJhDvw1eDTtjoDfvSvVCQtRUX6VQoaNyUI/2O+/CpXUW775vDsO9p
SsSrvWbB7hfPYa+f7qVa6jtT0TpN/cC0c+t/KoKFiy0CraxvVcUp4Wb6zlWmFO9dtxvK/bCtJ330
9uwQYNkgQRBqs44zg8PK3s7bcl+rVU79zWKCTlf5nOeohV2ABHjxMdfzxMor8gwCo3lCkcjt+80d
vaPbdPcjfDYIuetTPRgEoK3Pz+LJUHfJ/7DjWgTqLfBj09KPt7cwxbINa1SMIwpCioZRXvpenOf7
YMcOiNPU3Pyg1zp+IF+2+hq+Vrln2wYAms1wzNuXF/UPqb9WRlgpk9YpmUnn4Uw5LGhmhqS414oC
pDF/+b5mZCoKigLyEh/80YMY4XaOYW22nG5EgzfMkQ2j66XNVn2LAeouOpnTmkXBmorNZv40eI8R
nrAB3A6GzQ/p9ORtyU1FBGjpEWqMjrDiHwdYpDLw3KOFq5lAqFH0QvcQlEsoCXE58W312bSiL/0q
JQruhm88qnDck0iWIJ3MZ4WL7crIWRg/QKDHw6egX73kZrmyanSYuP7nF7rBYD16CTfnsndbQgUl
qfohNJEvHvfjyUUjZmkCiAEkAlUUagVqRYdQh55fYG0HWnxko+gVVChizEzfPMR/KNC2SXVavN4h
HBoBOAAwguXKmnvimmwtb7SLv5/p6IupNXc0mcRshui5H7dJAHREeGQI/IJYZi2JWnR6sf590EUB
x234QEf1qteolj956YOGjqQqGQz4OH6bpVZ/1iklrz4y3FJyJMc5irBMFQAdOEKopFcvFaPzaiiH
dAImGYlgmm9/eWego0+JQfMLc2i5kH4HBVKtnI7Z8+LAuKrodizZozlegNrvh9RYT9EUGaglt3N8
EhMHU9raMelOnEMESEQGwXGqeukffp9Xpo+keLAnygl+/ftARGBwMlYAE5Rzu9OJixfZTDTkhNSh
ZcQWQZ06O9yKVziafC440O7U2Kvd0iJKN4HOhGy2nJ31lK3ZbYek8y2Rsd0YCzfeBpG1L+tD4WWN
5pWRaKH2V16WUK8l7fBe9jL5ZMnS+xVSh9KhQdSUp56RfZhEqdCQOlddkVckRbBw4fnWSwxiK9vS
geUhDM5v5ApvtFNez4uKWTu4Ze9c6IABclcBfA4JJLXOAIJHFZX4KOGcTD24HIYFpWKTJDQTf8zY
wc4g+5lpWFR3V7uYeJt4YBfvZMgD5xdVyCgLsPbA9dlKk/yzw5/gnIlOs1MVl7fVTNQSShyvshcM
FDHFZJBac3/PZnIpo74CA3UHdCXmB4PeabsYGoO/v3eBvoi6fN2dylZA1Tew2OMCqZv/XzdKC22t
nm1wZatocmT6lblWzuK+Zb8EWwtBFKjv4e6SIzFAuYHDZroNp8WhMuMbEciOBRJdoIrjPIjjyAFZ
4f9AwOwzjouR4Pp8LrjeN3/aoci6Cv2LVTHubTSTjipqx7HvdKJWvqDtdX4wJ2dzFtsB5iJpFLtS
EpaxF38pUDvx9steeNisjc35hIOVqu1jnZaZ8DqA8HKCpMaT1csT6IBGFX6pZq87Jomi2QcgVa4J
IhctUbNOysfy9R2dJsjOcVu0/Bm6g21i4u4F/lzidhSaibbkS6uK8FohtUd+4EEjh/HtlAPRvSri
my5jYoFKpkxx/nbtDxeMepHQSOjZNLCn4YCv6DG02QggZY0YHvWwitmQDVYgg7+RXY6lMwSOPsYr
K1IVRjT+rjqI4a0wh4dV0yc9khI16vPq1IeMsYLHk1JkufVhfdxfrt5hw4KyeaBhLdboxlnvPlZg
U/47li/NZBrvsc26+H3uNcqD2PVb1mVbnJ1NlHxWtQhse7ELFrFqz0lf4Fg09SlF8AWF7hY7R+wE
YZNE3xjmH5Y7OxwPKwOL2yaZGjXsGLw3aTvd2I4i6f/vxd73yayqH1e3/7Vuk8xNqYAaYN/m5E21
RlNJ1QgGww3XEKXW+t9lBZstdU18TK8eq8gqkH5k9Bfprq4owjfCvbHneZOIEWTYiJwkvnEFkWSe
o1LdUXEH6uSQaEk9eOtwPY4Ps3WQ+FijXLtydzWPRuSgHR2CobGENB1nwxbS7UmzKhZBR96QQrt8
hd7+PjS8ZgKlQLeWS+mWwLSrm0BUwqyEZk8wwNEzzVwiuTD6xbJMH38QY2zRzyaLX7WXE+ngYqfO
MsMmWQZoZJVII/7TCdui4p+zn0L8njJk7A8vv4ycWpCoJgUeT4xmz8H+XlXTIKJiowFvIaSkWSXU
tLHq3mZp0hK/LqmKMyXBpBZAtgzhNvcQkZ2tJcFkJB/1lYPrf2xaH3CMwTOXx5Ns6Jgqy5WzNiVy
HwzKMBtjNWYENi8FYGKWFPJuwJi2t52swfNyGMrL8FxP6XJutoAOcQ2tdKzwmV0w6gGgmDUflOqk
fasaXO0peMrDSQSAIz995TC+OoxCAQ4zLmcFmEIZQ6b4wfKqwF/bLSx4+JEwrEAdr7ymanN9q8HX
0PXNpHmOvvKBSp8VrBZJHyAezNqI6a/3vnR4jiTzPinP7n9BH06SFHCSKIc2fl9ErAZll86NxRb/
j/FcRveVClzMbjFqNtpYhZKqSBxZmMMCnksttTw5jePGPWwYoXlRJlRSIBgz/4gzF0acHFn8tqY1
xI4i1k3Jf8bBjZC1AFV8PsORuNBMLJUg+G1SEnlXvVhFGxL3XXtIQvxNEzA8v6z79WJyBZj8ceOV
XbWnWTnzoeGEE3/37vqF9JAv8wJtL0HXXquyS+Wumngj2MlPMo0UHy0nyRTCt3kaRD60/O03GIh3
+I7LGJU2QGea5YV2+RpzF1ZAiIjqNfm9QgBQAh4RVM/i3sG5SxduREzYWagJYDiPaGGe0wTzF1Ym
ARqbAvvsqBlSu7S0HG5wHUOfrklxXUuMyQPnRx0MnXyYxznVY/BkHStYai17hZU/9vDNfUHO8mv9
X6fyXnzw7oD7Fk/UXSO/5EmL0rIh85IiCkNfu8G1q/QevJ2oV1pbbbZkdBXRRgs8WEzkP0f4+zcG
s4TTd8JzJAL3jVYRTiwZW9BpnmX7BEksDfai+YmP6oOMVGzSjSRa7q8RoknTbW0xtV296EV7GMsB
pdUPIi+SgSOM6QLe7KUWAZzdsJCBfRVZYOar32EKGeQ3OHFXT+h5fKT60D0wSNWdY2GbnvMz//m7
yWp0HXlkrGVM4GjNujAxNjIHVmykFPWaTrJN7/zRKYoZIjl26SP6UjAuIdneIviFELmQAyk5ArvI
nsyvxzum9SnSt4Um7Ycpvjt9UKg6Y/xwdCJzOM4Uhot+xKD2W+SIJn1Tk4dOTw92bGkMpittsf1+
W/lSMfmalWsbgOS3pPoJx1Ek/mJnPaevf8D6P33nss0EWACdBtzWZuO9FWN/dteTJVju+DTAOFws
bR7Ab4Do9m+9WYL+B/IbrKVbtGXKxWs3piuBDZigP0GAwzV5zzf41ok6cXfGOhFl7wd/AP/+0g3m
tkDIziPoOr9C3GvoCt4yaM6QNvEQHFHOlzzMotZQHXdDAn1EmemprP0HT3fo1IQrJ/zl/hv5cBOF
Bw+p5j8gcRLgrrlsmsFTPSVR+uwWolUdx3rHzTlHDrZY3WjHJN351Mjep0lOVVqXRz+WhZa/2hvq
7DmW/qHXGB5SmagyuspuBvl+1hqyJZXTKnEuM+fPZaEOlJk0CanFjeTnXP2mrXM3Qr4k/a8D6fon
NouOQ7Bcnnatmzs0w11r44Q1PODFk6WQ6JpOkoEhwaK8diYqMwcMCqaQl7gRqrhxMqPIdfqMpuEv
a9Ut8vCVvrh/bVNG+YbCykcCRbjGJasS6e8fgLd2YmP5PaREASPlVWwSNgBSuextBBANH7Z8R26e
EeF+RCHLYdJ12be/OA4v+kswMcJKGyBtm/FSH7pNLkTnKp/+QoPN/8yBIEHoA1Nc4WmQCe5+GwX4
DxnVVQANTjP7TzWuw7Dg/wZ7kDzoLBwwZzvxeLRAqCaZ+3f0EPLTa/ubz+liPBC/QNs88+DV+GRn
plPJ8nxabHBDl69QfRZ0PsY4w3keI+mgDvpZ4hRwQUXOXALwj8HiiS7OAMqyE9RR2ExvwzVkwtAg
ah7cvcXgZE5DQbCKqJa1uBoBXw/aA9Eqzy5K4Ex5/IFJJTC7lkfBcb+COWmEtq4ZsRqoLAEHm5hi
20MnIXjAJPJdWvpmbKwL375ALEDIH0WALbqRX+ZbB29ya0jsQCKzwgzMnl076tjU+EhomeNN6lF8
Q+pySYuy5I1TTrlfDBNesTx8o8R+gDHQwc/2rENAUwawJ95ls1sNgt8lK0kzb0IcfOA3NAAhFVnz
J/6C0uQnpUpTFGdJlrgE5lHsqOSOff8NYwD/IF5WaqamXm1AQ865o4WM7APnjFfqSH56No1SZ5YC
8fz/5RGXcBfe+QvjfS/bnTTwT2BPEyv/753qyRe/BtUtK+E2eQ8pKOoPSaNcLYu4fHffINRUlEdI
t4HRiO9jt48qNVpThZNPyN93QhGa3WKouip/XkSh6DMt29BGvuzB91qqOVPkLdi8uqbUKI/dLIyV
m9CKxM9mYlN+Pkch//BnAoPLLQL4gtfLQeuTWAe8fmA6DKJzYffCeUXmQlNUTUwVSUpptewkrDkw
Lg5ersDoTY1SGVP7KPv2njSO13LWZ/EtQwZQI2guM3XNsD1JPn/Z/pG/obxt6zYQZhXlJEcf3+P2
bljlTU3j6ElMEGzY8vOMaGsGge7DbeWZbhp47V2ceIS0e2Azue2myh51CBIYz+Nj9he3drSqriib
I9hlHN++8vFdUCyWbu8q0d7jh6/J3lUOKCgLnrkIkZjXMC26nifsdBQNPvi5f/4mlB0Wc6hSoJnu
mfBkJRQo8a3MYrFOQVHK3ymMPYwkDvcjd8+4VpEQ7P7u9asde2UBIeEFRYCRQfdc+m4movudFn+x
AQfPxILXi+PxKvL9Lr13GFNhxkAUuTgKCIY04rgMsH+heg4FZ3JxZttpoPUSCJjTS2tmthomFdna
EVKhVvT9NaMMMvLZjU34cY+LTjr/veC0I30DJ436Ks9ECdXMAN5IucE83ZqKXesYAM+ffo6AQpw3
1CDXO6eRp/WpLGUMkDR2Z52BIUB8JQeS77xFUootag2dyHuOrKCZmycS0L3IQYdvAPpY8urg+euz
F8kt8B9FxZDsmCP/rW061TL7EI1ywDvUXEE6hrmVAxBu95kCI4BqFZGJ5EcN0KQEMdIvFnHPf+Wk
+Kaf9g5f6pl9dTpPbXQ3dsz+ZTkyAg44O7BcbHt6j8NLCm8ZoL0j9v16w3OPDUN/SPdFW/yXNOm+
9Z5oW+QzpUAJGSD0AJQB2K4SOd79kut0cJrQ7sw//YaHfKPdrUHawJGypReX9tHst3oliKXWquoG
FnYhTSFMaxSWsxIAtHg1EuAqBKFfLlIZPcqGjVrbb0REPiThimKtcyPmH55OPyvjsg/mLvAQqLC5
vFwHkzrE+AJBWHG0Y2xrnMamP3F+qdmD3cYJYyXPfJOiy5SllpDA7g2fzOb1MMJES0c/wBuQclR9
aUlig6yWjLekkIOruPYCQ//cH+gZR+NhBBDT2YI9+WtxOKvDmksCY5YvueRZYyWKa1s7FgthqQvm
qzRDb7ood6pjN3tl9tfOm1Jv+amxPQHqMyMwoWbwHUYLPtJEe5FRGu+iy117wvGyVsZZdbYe679U
0Aai4nrJcW6D7E8hN1CVDl83pnDFxEdPgwgYLkxrcaz2b17j744K6R2ndVC0JUgkzyvoFXhXQrVC
7kyf28XNXnk7ZirB/ULZXIfKv5NgA8dEz4m082X8NOqxVuKEwPrltg7gM19z5yKwenkQz2+eA4un
fvgYw3Yjv/WZAr9LtIw93dR3k+uF8HFDbk+u39hcxP7gEi7EzsH0rhCTwr0u4uhU9P3sOahtuxcP
2gOfWfY13zAEtDu6a4BZL5SYAI7EeV6DQA9FvNjJ+5qjKk3n1UDPb6FAS5yYCn3cqeLkMlTatdEi
UyEIt+HuGxbhpFFE8bp9cFYq5j/7sMuqzC2IF6X1uDeAocgPFg7m264aFfdMCItPa8/MCSLydgNY
+q7VudJWN5i6j7t1gdh66q+8ce9uwZFA9IkzqgiVMZXr9awvQgpZEA71ZsV7OxxjZ2qVtB5oT3lB
lKJgne5q4OPF2UC9lppxFH5qMqw53dNRaVYjlpqnPlHQ1ruKYlF8R1eryKAaI0o0vz7mYhiJvlMT
XhcpVixQUDgi8i3ZaRHA+ItV7NZYjPDXObIQ0Adoe2Q/pT9yrRnWvHEr4JIkPsDPiejptGa6VjdZ
2lofRv8anVD077q8cMyL0pste4QsbCmBB+fdeTif7ARe1lHfoiTDHqxP0pdlvnyGaRAEN65ge5ZP
qr5jAZKJ9t2/ABBalRUwvNbmyU4pG0hi1qVsRB5JBBnm7QLrLJ4rEe2baN1uczu5/+GYSa63amDm
oJUSFEfe4wIC7UfBL89EfDYWx+lp8hPmUkBRlHWhckrWM4H1nW40JXXXcrU9em+4xzJKiuuUH1Th
JNl8H9REyRNqhy15csa7SSgCYAI5V1wAnS9faFsdGKHzxRbfVbj5isq37RES6Yq6xZ/o2Xt0KBI+
BDVwtap9FOz/8qwcX90nX1+4DSIz2qnucWt6IAMapA2pz5KL9u4C/O00YDhZY+d1zg1cPxKVNfIV
AwxLKWaZFEapsWcI5+kLfH5qTxkYAEAg8RSHHoc3ThvpowZQQeq6kWPPlKa4dFTKQQ6fbVlZFm7N
zefNxH2B0Uz+dtz015yAGlo8D8+QbLpihJswB2HjAzcWKAhyyvX0thmXXwjdp3ueV9KK0c6sew1+
NgDhoIrfx9DwiDvZKj6q0wCl2NAB8nbxq/6BM/yJ5I9HxJj917D/6+HKAkpQv/pORjFBsMtUSGUQ
YFqgDKdBd9A5d5VOmkBa38BzbTFmhZ1BACJ4I+Vw2WHAUn5Qq/DBY//zSdllrMzGobyN9dkt0rjx
HojyhJCVb6FJ977RCPjjR9cFOLEniS+SJ03VZmbUGv8VJZbzQHaNXx48EAskatz8oRQAtv4OkJ5W
xMcSKMyuzHlo7Co1kMCo+nSWJIBmv8i2tssu4vkbz7mzBVeI4qEY4bw//jJ4lTbUqmI27/NtlaGL
VUZARhhOyHykhLLYw7C+wdT8YCapKnKWyBFa+86KHQfhiuAjWAiRJl7kEmJzGFB417hg9qHSYvPi
p2N9DK0Y1vSENvdwBYe4MsyNXXdUYqA4WwuWOwtB5COnTud787npBWYoNk+32UQ72DhszZGf0+kG
22tkiBPz66ty+mlKQm4RT2uFobFsTCUo1Qucj8LeTftp7sxORo0p2qNI86d7+OLYLZJi1kKxmqBp
DkqpTk34NbKB1B1r0WKp99G5Uodn3hrdQK35xcEUHlsg5LCSNHSQ0L9E4+zE/aiH2dtlUKTxsnvX
M1ATNZv1TqYvmy010y3e999em0zYSvdZrrkyg8DWSf8e9Nsxn7vFgfQGQlHLshLaXW3CtAwJTTgk
abTCPgmrrebPeLpDgdHefSvzTBLH8rGnmqpFSPoIi/nuCmatUFJwomjuz3Gqi2uV5MOU2Y2uwwBd
5s3hpokDu9X+zzaE4y+Rm3RpGL71Je+5sp87XbPiLbw0ivqf3p4z1H68xGcvsAOl0eLu383rNGoH
tFv9i0wJKGDo4nD9+P3Fe0a2wcVFC4VwQeq5hcmqMKBohZBrPdzmQB5EFAxc2Ej0ce+RTJrgrNlM
gthtfiX4kqhZwl0uz4+JMILUp3SwDUhowOK7955ySx8ofBltvPgEfh57VtwCuzYbFH9hA7XrnbmE
s3nFbB3uFaJ2o0oQH6Q9S56o1huw13XqBPaLe0h9AT7fNoGqj5hVXDp1FkTOVRA6hKqLMY8j8pBd
ycTYdOyDOwvViGWThgrpkFXpqnI/HXmX+N9wb3IZy0OioY+NId4m8W+LJ7fk2H0FKoZRbiQy63A2
egFAfw6lilGVOmhvQWEv8i4Tiga56phEfIE4rl9d1qi8WvYemh/RtK4yvoQwx9KXfYUk6qOMr6Fo
7+gsfJhdqa8JSDA9sxuHjuuKQ+HW/HvakXb0r6NGtpZFWp1lSnFITbbXrZ8BosnkgNfDBbrUe59Q
jv7QygX93138seVTvtdrKvqg5oEvI1kAKhFtX3DRW+pZ8E5Ae3yf2ApWXOl+2xKIX6YvjXjqML9b
P094Ns/jbpo8N6jgze5qF5W8bU7C4+qD5e6ZPKOSl/Zuc1ub0D1SBTwGijizQXohzRnq7ywc4ex0
K+bbkcPFdDFUfhkp2tJ5VSOdr3PKsKvauUuMtqLwQphspRUudRTY9MDyKcXC18nQS+tyAvhvqrfI
r0tX/jaNkdiHnodZkrBb00c0r22hb5Rkf+ezIg2Xw/cLmL6orYGhRFia9x47kgG6KzEO2zyjLiCE
gdLkHp6cw3IMk+uHDmN1XCA7DU1GtVXXvXHJCUhmk9cR0Wh8InCnLUnTNBIYhvyd1r3S7xf9fANf
LSQCOjlflsjHBZvMSw473CUZF3LsXmRGZqn8mydRI6vY3LwRQoC+QXfl+uw8yqO5tLZJS6Yu54oM
KR5eQg7PvaEkjoagjhxZeopv/yzkYWL/pBPDuf3iUVphgTa8UIuz017EZToqVzQj7rhC2QXa/kQm
iW7ZyXpCN4mAsQsEdR/A7sdlkrvWf80OyM38U3KgVxr8DIhkIL57s9Er6MhAxFtb3L1S7/JE+7qo
wAxsuId942Vl1r3FKTAC5uOFqW0o/OIdQrvFHDkcScziU1sYP5VPLvg0ztWdzoSXrQ5etsn5GQqB
j5B8Ge02VkIDAClUyC1lcCB5fb8O0x0rei06ovHGOYY5OC4J5hDJvNkXJOQZowaSLw1yTCu2TX8/
KfT20IdMm2TymkcGE9BZLEHZsHMSTWNQGSswrMLDW7c+PxeLTfpUrUvv22NuK/TVggMy2TjoxzOe
o16ZQ0uul+Mc797fbJGMYgZqu2/gbVlILmRLOgYOqOGKgxUSSPs2Ewp1OwuqP43cZcAmInl79trX
s/10+K4qU9O4m5wbinqkgJG51bR41CKyJ2kqKdg565hSpWK1mmpD+mMXYSbZHN32rshtZxV1bq01
lPjb9AXFSywA/pSjfl9l6l9c5tlHU+BXsMwfqv0p9OSY/UfOoo0KKBeY/wz6qVwddtytCoCtJiDI
E07sGp54W9wc0k7JWiIHgdj7r4AYp2/FLS24NXlfzU/CHLJxJksH8nG397N+/lrwtsfiMD4z/GwV
akWrLju1UYfnIMauem3lSwdv9YekbzVNT8bRN7+5qo9ewZYyUdQWGdfLmaeYhMDn5HP92XdtCHGO
d6QBlnNUsXVIIjWGOTTKlwwzR3A0DV0tEGOpuVU0sXle9X/xrsGsRdGgDfpsFz43C5V4F2RoLr10
9zApPmrtVfMonO1Tj0lu11TOpZFRdLUtoxlL6fhyKxLikelZij0VNaU85xmOayipUQJymQ73kQNC
fJahex4KZ7FPTtJGWAJZA82jnKMBeUqyXIAqKcp7LrCb+O8eNVYs32z/pvBXe2PA0WIcsU3nmIEx
Xq8rGfroLxp3GUp+RX4sq2JOFpCvqvP413GgnHaFscnX+BUWss4PWJ2EuwuFQRuofpHpaOlFPyCx
3MVvjO4rLFRkR0W4WKGHnBSlwCmU9qvJE+ZaOFwlnZ/ET9S232CLhTmBi9ZPhxqlBwDnQOegKLJ2
jGpT6b3R4B75iTBas7TcIyc1Y13yrkeKNzDz0a0OBvDi96WyUaelUPnYa30lzuyJI7iYBaKdSNr8
JtLuIGWeGybUjqH8oYWg0V/TifaaSMrW5kd5wJFipjIeAQJ2cG4rWe4n5iZD7OYty2y56p0aV0aB
BkGLpphQuhqzt/w+v3pa5EAio8XVakL4L3BNnDPaP+XIAQPS4H4m4BiNfBzcK247td4vt77zIieW
HSHxSpV1wTOUbJ5e8ac/6+Hh/D1gtpKX7XwkHa6RRsnAIrEBILpJXZjKyzevVsqZuEkH5ZRgEffr
UqwCXaqbuyxlbzGf7hlJA2LBSHP4Eaa/1yxYzAQ9a4NcChDhiLhxkphiKDzwA3o3gjntp7slVOcB
yl1UX44SrYgofR6SZ74SqVf50ltVFQ/M+ynClsf4R1sw1oGwkle/79zbPWkfKrK1NtJnKBXz/mXO
tvi8L3V6+xKMX+Ch+6BQV6JHNhcE/xJvMltYUS22bBL4y08exZ0JIJ8DuzUcwgN7KD4hCsT3cE4Z
6k2rvvbvs65BEf3gjybGGbvwiItcQ0QLJGlvMGW5pQKeO11lHR7XkqQeJqCn0a24NLz41RVB9LB8
CcW9CxO370k3wuuWwmbwqlBpp+VFnrUEKjaSdwVZMBUCCSmfw2rZXTWxB6vAhmzZxoG76oTvUf+7
vUQ2YupFXiZf5VUHKM9uunw87b6fe4D4RSt+xldB6EJesqZ+tcQ9VcIDU/xrcDL+bepk1AnAvZr/
XcwgS610DdzjnCWaIR2AgCQPPiXC2GUO7LzzKcygY6kaLWLr0BVgdnemxs/OKKpDynSZDyTzYBRV
DccIizPq1us7UR9nT/u2jOWKd3x9HRok6lMcQmJAgJL4roGpX8wujVHX/yfOCsz1xqDTMkHlolYa
JUFgiq0axyqW4FDsZC273EW+hLFq0IjYPuh1/o1AOEuNQluPDJTDKclMAPpsfvHNIflnuh+ci3An
B4fwzzLa/7CWdodbzCiCQ6V+Ldmd1wUHBlEWnYaZpI+ZZy8jXihw81OrW83iwWj8FCMkexBpbGYG
NPcUtty+F8isqDy5jN14BN3NalZ/65TewFHlPPhLNXbBYtJbu0B5cwIgJU9KxfzRrqCaUVzvnxUA
DxHdhfc8j7GzIsP1CJp+SjlwVrSMaCuMdyRGhI1CokWR+3WGAER38FptwHbH3SWcJ5yhX1v/LvYj
DDRJlRbJtz8hgwcqS2fD6T0fGF0yhF/qSZ0qCsSb6QWGGXKrxynT2asXuFBAwks8yGlipr/CxQ+3
8oCLghTdO2ovAkcYBZ7TlZ7YHGUPuu4fzGYp2m15RjSKWmfy5LytStPi07gSkYOB+zDtZ5rkZUkW
MtE9wfldi9x4IXMg7tmoMYJTlsuCJZcpWyls9b7bmXUiSo3rGXV1b3sLCp0a88cKAbtbK2X8D8jF
PCpyQskVWfiIxH5j7kj8AICoPgVqW25Gp8+itYGp9A09FsmG+5WsVah89zCtb/XOlZ3ZKoSm7Bz2
zhS4zmgAP46GcbpkAwgm6c8vWpf9HuQ+dh17icBzcRyJJW4t5Lf12EvTh2DBFEE3vW8O09ewZlCc
D144Q3s9iTsUpDaEp6Cd76YUEAz8jUIBMOl4MLhiCuNJT5ThuNov2OQlJ9FR28weIOu8nrUhPh7g
fkmoYDA5mnGaEJUKJpQvr0U9RZUcg5E4jSXVD/ICOg2u5u4mkUZ4C5JN427f9YNAZzlMl9dhNLkR
o8DUHPSopvoFe4sHNL6X1sQwRkzOFveIFmJpnW8FWJTa2xuGK++Vm0b1fMnD+JrRxknYjjqyxTHk
5pMR02/Zev/K3hzMrXaWgktwyU3UgURGl+UcIw1N9wKCCqX7DGwT8iqdvy6h4j7tOCq0xMRAUKOt
xPx9vd8JACpmQBxtm3RQ+ILHh9q+JYFtP+cgx6F9LbAS+da3mL9tYirA/l4Ahh2DEK6YaK4vsKic
2BwiNwAmQnlRjXRCcbyrJEXg239Vud8JsmTgkXL8EeWnnRM6GGBHKtJsTbKmzmWVX/K2nNlqTIlS
rxbJX+F5D8G36/OE8iIhz3SE6Que+JfiaSUTFoqwluFn82+sWKKhHiasVWdC3xlDIrhX1OaTF98n
UR3vgzt2hQbvs64R5t+I7oFhDJXhAchwJVFXP782DeOgEEoK7voTq9E3vehzFveRvHMTh9VTeFQu
4Q4k2N8mYvZXn2WnGhkVma4zs8Fm+EXQoiFHSRRWdL36spzDhMUauwZrkNheDTAo0yN28c/O0HT2
EHi39QBxDTJTMfN6BRROA4OxvT51WRnnnFLJbfN4F846vje4b5Hwqc9//8jcmJ2lJBti83XmiC3N
7QHsR/0pfNqeKYOgCz5g3WQyMS4wUmNkKbGXZ+pzKDQjaH669VupBixtANNYwPcfwvOA2u1/agpJ
NMji8qmGxWZsyV6o82s2yxgUItQL1XviSh1cx1vuCEoCQ46W+9nCXhueib1cC5cxAvlG7KmwDbyW
QWf8OMZeppQpNb2QukTSSU7dSoVYHUwmB0vuESXrDzc/H2zmdWwon3lE70u+apkxhf6+IoT+azr8
4eOh+H2pxSu/vi70Uc8CdYYRjtLg6746G0+j68ESnBv4/M9bAsjc5gph2CEOzQewn22iG5fvrp/i
5RzFO5JU1dhYL3pPJr75kNrxHAeUj5eNNwKIlyY8WJj63ejG91nYfyGt7690JyNAXTWGzsLykFIJ
hhqt8WUHnk1ECgT1ER3isQKo5zonUB/aJL11z/Te8DbIwfKfrdVcGz2HbEPvm/LDPfIxxUzwkPoO
dDcvY5wI/AmkdkSQrl1m+HtUy7ca/zWdWEgMewoLtvpAkUaqJ98+CffObMri3kATy8N9x9HLtVDw
gyR/0BOrzljAwM3K6sX3tJP9gBK1NzQis/8JFEfKc002LCQQqICxQtxJONxNE2G38vKnF4cvRh/g
iNumRRPvndZZntp06EUZzTdBQonvG3Kmrdml4iCcY04AsVB3gxfuRYdBTqvGTtYwEEvL/ofdZiVB
vLJbesnwS8VgpVaDWZGAWTF7N/xtchsggwgawm2bIGBMA4NT7J78adXeB9tn5m7NXVCr/4CzEaPz
JcjM6/ynIXSSwCYkVXY/lQDpRbNq3ZgrPos8jj7KH+IhZigjQZ5sc3plBSCrWg0DWbpeIwy9qVee
wBky3aTH5ev81thMenJ5Ho5+B73bEvfMfrgkbvii46sC6VRwrRYhqNT/sxt4oWoFJ9+VuVLl1cOX
FEsznlWqaU3tMEJd+lVIN8NPNDkWusUgGqeF5H/ImYBSJ5xMuuJtvfnoET+6CUE+BHJs169yVeyg
kn4QFsKntLCRRgoVLov/J+Xfdvzu6Tpn9sI97hqq3LnBO1UsbdZMtxlWQvzNU+1heo21Zw8cglid
x92+zD/gFJLCC2cp2Mj+pCS9+mtT/YVgKQ4G908ziwgeNShtCTIeGJAYcXB8b/QD/qSEPH/5r0Hw
MpXp+XjpHGup57Nu8yHknqiNXDoOiTQg76oj+hRk8ErXaGc+Hji3tNZmRcbFmcQPxAgc0GKlHhYi
Cd+88cK1n8Woin+zI1j/DBqXcNd1qGRIZM8mQ8ZmcVI5qjwnSkdyWAk7P/Umoqka2nNp9WrKsz3W
AtSk2Y+n3ZfwJhQfSt73IyHBVLMnzoOCV7CWLeU8maVY6weWEAZpJWwJ+UlR6xpryG66KGTZlVHI
OZ3F0iCzAriiq/q/rq1bZ2XNo821QUzzGm5YRu3dFo3j7t3PdUzgP6sjgSA/t0dJovPgwduMePJE
+XQsuDrTZcdFtDGwBxpJL/h19mmdM2euiGyxDm4BNesVGPq/k85n8c2G/rs0oBmJlk2V8nhSJk1A
mBfgyTcirNiO87hiuQuNQOmudiL6GZpM1OKcgNp+qOHczAYYDG1cTGiOk5nDiPMyGMXeb45+ChIU
tqkbheFH7ll1n7Zt9MarscKrUStiDKCqHX3oESvQCO+BKid+HXil/lNOYuUOMfHzH/UhBA95nsgu
9QKA71589Kyy7bccPHVrCHoLDWj/G/FQ2ncPSbQEP/YqrCgmI79oE0ecNiLakeEW6qVcJMT4mRFQ
8cZes+NLhlMYAzIe9uZSSC5TqWkhOe15h+uKi7Lj9z9hlOsSWuy/RmYXVXvksm2I5lyM53LV1V3b
5jgi3/pmyVf1FNldwHgMM8Te6DYSUvOOIBGSbgq1MDQVnOjD0rdgFKKJiB+8HXTw8yQLZCXeBuh9
dpU7N7Zr74svCDi3ATkkBW2a5ZwEEXEljOAIc/8z8IKwm55Mp7IXk/4ynYCjcn4xFPghyxb+HAhA
RuyaPNpN8vMzT8NTkrJ8xXXxU23LDi8zwgS3i9og3J1FVOgVIEu4as3y6ZTchbGDgxZqzQc3Hz5T
r8pUe0dES527e1p0r/qpVogHmFovgp5SDsQk2tU/vKiagn3LhNwZMkWSRqoIYbHR4m7/rXWwFFLK
UID7ipM8EkfKbwEJIJc8x6PJfxOwNQeImWYci2KIx6xKMFSJF7PAPM17YPPWLHlt2hVRiqwvU4ym
NU7myqQaOC63ynvnn+HHshhdfYVYCeVURVt+QcHOC+pZjab1YmDBZrKJHoPUKPC3Q8Fsy1D9wYVQ
yxBrnQuYR/bsWSLv/b6rjjTFurlGTW1sFta+yPMWUDTc7yMdnA+S4NqnFjJyENvXvioucPC/L1+p
KmUs6Niq+gst08BVwHDrmUZYFqZSKp3RkMxDR45pIrNIr8aYp7UwwiGMvpBcKRTXV+kuHutcjZ8Z
t0flt2R52VbO4LMjBdoXpfiHPrxSn8df3yD0Z81xc/4n2jGelAslDoLVDp6WIgs1867nVcmkLB5k
S0Eda5p4ZoOoTSCUmohWhqKaTuDBPPTiTbd3d69FDXmpABmKPLtOQq7zuHrnOsDUMaWGPsx0S1Zx
s7Onc9quDEtYWGgt4qh5F3BXh0kmPwnkCN7ILLivsZ5gKSGN2fUWcaWabPiQk1Ulsnb4xcQCKp15
5Xbp/rA0LkRFHTaquqjCOFkUkY9B3OQu6hq8dTpvtMPZfRaprGs4RirLSi3/lc+tv4RIxOD8muE1
dMqzZ1JdNDFR4FhfQ2raSmePEqdxrm1wbtGy8F6tfWW/j/2vFcvbj0rXxaBijj+F7Njh33e+sciH
yqpXZm0yHCuyhZAbAypUL5CGvG0X7hsRHYbEKazt4rNSA/1BbRSAIjGca9TfEKSSx+ca4MJc4rgY
5eJteraTIGmR9cPtk9Z/UiTZzGtI4jMvpr0ienv/vHAi9yoIm2u+1IfoJbDV8Om06z3/fVhaIjg9
PpXumw4z+Gl0Xf5CIF7MITQh+unGOuuN7808OnnVUrZ6mHS7Cjr7/HJf3ZIF8K5lvbDWQ7RJDSFJ
TwhYfN05Dhs0Ntxr8ZNR12q4Du2Pggh+f71bhqHI23eQWG0+YF7MRQWqtMdWVuf1a0vJzoDro79X
TWP38xgzEyt/JQKnvEWARUPLZZMSDOHk5i55u3y2BcCKHt+PK37vVg+xTmDima4BLfIM0Gk6BmYX
I2jsQfEIcv0u8FJa+FU1BpefK6UscfuDu+zjQ6d2oVQVMiNjCb2pYSa9M7gj4YCNRQLWjNU/D1P5
S+UIR+9sq2lw0jHNHCu3SLQZwGrfIsKFBO08EdduQRuxOESZFRau0tu2vfgY3u9akJs4NTt3rQyI
65QEn09qLDrvJCF0wAsvSyGjFqoysYp4VjExGMX7MXYe6PrSZmdNbMDQ3zs711NjGjuYok2uqpj9
NDOTHzQV8CzGWQm3496D8vHhKB8muZh0XSU7KzaZ27cBworJj1sEc5gWUQm2LC18xrwj4CWyai3l
KaW4B475N/gjk9jaRFPcLujwFj4lZpTBRf47My0QfMyETseWZEKGUaDTR5ekagk5CBA0dQp4dh6G
BXtBPzv2reFAGATAfxGhaahZKax+uh6pPYL2vMO6bH9Z2Cbj2uJRha3tTS6I6DyKIW2rOahMvnnA
CcJrUlUA8dL3b84kBzh3gYwC6i67rC6ukpW9gTKiWFQvWljwpmnq+4fKz30xJDe8dZzcMgRRgT4k
CFG2PDYDFTZQus3P8TZmwLuey3LVAGwGKBHNHPuM0sFgM6RVS/uG9IbjmuhhT+LqWLQqEvfUxzJP
zuGOB8kIyo0EaPNCEHJQDNSIkdPFLFFr87IUVuoLM5DH6b22nMC6KRqXY1Fwcs6UHzGFpLhhkuTN
uSzQtWe0/JZBeASouI/LlzpATYeoYC7yuKzXJ+O+6QkO7ZJvqsCdvxMZMm1A9/iFfp4glh4j1oUg
oFxo4bzR1WjveyOAOrlX67MIryuWdKIMsUqM+oNuxZUbQ439DJH41CMyUa19+mpHcot8XHY+H0dF
xMxFvugtDmDTDa6i3a5X8urM4I0pr0/73cSqVVRAOi0MhDk8XWJFH1hNgw0TmB6eLQL7h6ez2+uH
gaJbO675Z1JgZzncsE0WQ9jbLypwGX0cOrTz1JowIyMSnSmSZvzgNMAHzPQNu6wY3KeXC1cy3fPL
yYnI2cKTYbAyiYtHL44XiE/UpW+IYAM3HCQ8GMWkzc9U5AHGbvgzLmNdEjE4rT8kjAcmspmsEQ+x
JmRu+7kcz/MqgSjpjMwjS1o5WAeNuMoeYvEndFUH1+ogV1edBC+Wo4IL/sMnCJ0t4G2BYfFT53Kp
JsnGTY0SMI/K5UAk6ukr/H8hYHcT3rCy5nL0cmpak8zaHUIfbPOjoFcZbgBQ7Jfs8yNuWA2SIRfE
QDM1nrUpY50CHXoNTXiWfULuMFUc2gFHlg5BcaAH0ffuuouDKoeOMScTXlnBEsEPCHhjo9xAHnhK
rqp43HIEcdmboxcLTPCYBcD8SiOnG3wsdam5EgfUCDJ8DAGWLgO92F09hggVUUhH3tngEwxqxnWw
42hWm1LRJW3DoJydx8HlOzH9cptJkZ6BEhFipj1HIbGTZ/k/ikCpQ46cEnyyurYUOgeFK5RhQc8v
7mebSDo9KYUrEuScZFawl+hiDL2VIlAtLwpDincOBOz5SSmUniM9tKwFDuAVCnvRmnzpQaHNvlYN
4zVIo+yxIIM9FiaRAXG6NdRpx/jjPRa9+lPUmpAutwgIxWz5enX8ls0rD5IaMICPbfIwJJrFjgpy
JUkmhCRAbJlzX8WaGJpjmEgDuLeT9u6LKD+BI/EwhC2NBwitj+s0+wRj5bVpef2yMed6mqzJM5QU
9ePa5XsrBRalRSeFHX1i3bqSTGMvBZw0UEBBoBlS/Q2cDYaL2dWpsiwHdQsxIvYwdusbJb7NJjrI
K7LzdFg/+IkTaxjf4w94a+3jXCyliT3xDUJ6hQFd0bzxrECqA7Zj69drsARMypVLceUJecZh40KJ
e02pVM12VFLNZo4u0gPfLOA91aWhou4isLHuHb9B7uFApyJCE1EXPM+kFUik+phbxpD38O9j39do
Gd1It0D1xrvg8bZHovrns/YqWUwudxjTk5+84s+SRDnQPqx+/Fxrwyfz91wwFFf9abDqjxPsiW5e
xs9R3SS8Q4BXabAwxM0Ej4u4ByDlaDRXNdBhmPlzi50N73JwymB8RJ5u7HWAxtRM45dAgqwub2qi
pbTFLRgIA6D8ojQkV3iygCZ1yRpj9pupteU8+B3jY0eoB/oI4aSBQ8EIbkejW4V79i+KKNSPKuup
8k1+NRPVBRzvskMn809E4VW3HExxrh7YavUw9yREcHei7o7M2JVTwDXM9lgSELwjdnPaKMyhBhZI
Fp9jE3XPEWgPnOcv66/c9GMpXGLVcWkCF3ZBHQQY26/H0qs9aJARbFRLFah0pggefK6sgem6z/zy
FmrRvhQpAH/BtT6oWhI2wbHuF8K9xB3Z4c8lYp2iSWLR//bdqUZXD5T1r/V5HtFbIuDhk97ryCvh
6EIiCbotSh+XKTCiRHgx5QRH6d0U8xfCIYfPnwmDBEJcRc9ZPWBVKl/lxVLdHQSNigm3lfkMscjj
ETlzbi5XQS4AaMPNhH7nkoGqE/bRrmXUxYPHOdxQo4U/p1oDn7YivxMychfWw8sJ7kc82X6fAW48
J/aJ3V1cnZUKAnJEfamDjUPVmNYFYHxeZ1BMMfWagqRabryMTWMj9ejMuGo0i3fe8e4s0BttgFT4
GirHvworWzsCBiy24UVGuowFG+pEiJGgPCCVQaxVitPJquplDsBVtlxlhb5A7F0CHXKwruRR9xJb
3Hkx7/lDf7YV2WraLYp4LZe+I0NRrfazXGjqr71xQqJWN6HZ5xC17N4o++Jarbe+AFC29xwRFbYx
F0NL3dCX0+4mDZXuhYtNKfCOt1RoH1XDoKBGyl/YyC9kL3k2JANx113Z7oYTXwLAEVStA8Mep5w/
ClDd8E1cGYDdV7dsRgSvM8xPuZQbyHCNXT5T5yu9QvJc4wIc7oz+/EF1JKZAINBMtteU1u1jsTG6
23n+wYlQtaXVN/ViyImcRCvfDVj1tBGEopBL6/3cCFVeoFr5bKcaLOXBj2yEAuspqTc96tuJK1on
bN7phuULOEB/MfgPsIrNEN7m+D00WxyhWuOSBllQN9X8giUhpx1/n+J13jghwB4MoeVCME0KzPgZ
b5aMozTc41ehkQJCFeM16w6OWJxpgV2AWWrkxsGGjUQYQ3rQ5XdGTymWxHFV9otiEcYCBZ+8d0FG
eqfIZF85/DcefAJGSAfPu4NTGt/b4So+8Eu/+thWijHU2j42Vx936AznJoABqH5N55HKx+9xq7Gi
mAACipqWaNjnGsJItfqv9ddB/UuAeGQcLGFlHegWTe72CkmbE1BHSAH6Rr1KCd3vSXYav+ppwkmf
dk5US1L5xjWqyL0aaq2HIEC1Jw1lRdA5/yqjH8WxT+Xh8uam6OYAeRQy+1mhv+8IEOKs4c/EdNgQ
S3WW0G2IqoI0gxGwnRc/x8lpx+Ta+fZA7zY9AZGijf5FW33WAKyacMgdPQXK19x2YsBhM1ovx/OR
nrlE0Trx7ObQQkj/Se0AgSvTqP1KCk/3qu+7DE6ls9Cj29Bi4Ly5qKtVklIAAYh0UPP8KMmFyyrN
53eiPzx4Ui7xKdrCsZHScIRppPG+adN/6LscJ6LV1BlKbbPEkNt9SIPvIfjXEmQRwrrcqQSjzVhf
mBQeaiFB74bMf1wYswDteE14esW7W7TPhimtrGLxCBAk4/HBH/KKi0CL88a6vLkSPvFSmBXi9nsf
GauvAJqaNXiWld9T8TpgQnJsQgqjcTJvJxrPVuZnRRtlKhJFo/PqY887XXs9VLrYgdUmyJibEZwT
UUQldBjJ86ewre4oviZH8TsZy3z6GE9CIGipoKhZIubeGQOFJJYmknuVERvMusy4oFYIULo6JB9+
TM5UDWNao2zutAvxnCffJQ0dYjZ0jN8HwIxsIyZ43ZHqSzsblP7/WWBbpc/c+31gPO/WY/vNXceN
qJBfiN2d7y3vf5lZgYZtWH0SKzfExLJ52raGTRpnh7AtIpBquSZjVkKcLqhtaiFa5BritC1zgDGn
k+RzbOaSsd2W8onHqxmdvtoA4nPUVFG9j5J+3+3g/zM8OZQ9kqCrLlGmhbxK9lM8UJV08z1aXRzk
i5984u/epqSlsTc2T3qVlMlYUR7UGAit11GLFQQnUauZINqhMdEvq+Cm8+F5jpznL8Qx+H1EWQcv
jfnCPKfHtvvRV5I2wT2IavzShTfftciz95BJ2PsuhQRC/9clqBublxkaOqM96bigtDzGpJn3438S
ZSc8YspW60Lmis4w/G5F2Ci5pM2baXgZUFt2j9epfP5j9tYoEhSD+YtXtX7W1OOuo1CWvi5/dPa1
fzaNeGQVcSFrBmx3Ropg2dim6DkY1+XowlikfYUvIRAKV+FZ3Tq8HMx7VD7ps9HqllfU4RWJeTNg
6gV/AxBHVGm0DqelGxJ0uDx04gmkDY5uftyXvDhLWCXE9X/cBtz2u22BwJqDjE8J9mJzUiIqrs5v
IPlnKAdcIODFgjtv1GB8IwkzwGeAOeRheDWtWbluuHKc9k7C5RWoxTkZiKcspSuA85mYAG+lqlEg
7tQAtfm1NPcAXeRbQPIP69+Qx2tVLXoIp9CxNHzDLBl6yZJmFNjJSE8mHP8x3Bv9yuocx/vpdaFQ
TZQ/6m55z4f13f5VbBTlX+8mBY8qFLoiVqb5N9G0rCB9XzFZsTnia8b0QO0UZtTeLMjfu/A+DsGz
OR1Pu9O4PpEzV5aQKDsPiEfdFjxeZLQLn+ZvUGrLC+cdKUSigz4rQXb2MOB5l8U7Vcbisz4LDNPS
brl3gVEmd4R0UHh2A3oDjRSGLjbtqBcjST98GmcP4v/HS/MJP9ZLmYK8DjwJWQJuMI9ClQcRjgZ0
wyuZ3YEPhbdORB+BpGOwX0o0v1T40cPFvc4RHuBT/laaicFysUmanOq6moDyNbuFZpqp+WSa5qz9
DXA0aKsdBz1uogPzbAL5YITEDGWrOPeS4+6yFT8yK+AfE9jlQcK7AMS1QtzSYRCg51MUe6gGMemH
wpehyvLmwdoZc9/1VmaBpYgBfbNieTwO/zW+3i5LC8xYKNCM0BHwe98PgMez1ikYBjLyLU5GgpPj
o7XeUATYCGo+Ul4sPzRfJgf495s4HgoT1boC6ixfTxkMYJCtEFsN6R8vfuzBo4pHx54Y1zmz7MxD
gF7lniK2vG4MgL66O7tXaos9KF7JMShf3EsT4QYK/ueVcrV7L2KvmkivzQklP72Acpbf98l/8e0s
vXEBioqTw76IBg3gxdvrzwxy0TmacxubNB+DerCBW0Oh4AcrgpVZ4tgXQKX+bV+fi4Rg7YTNAXV0
3WwvPonF6SoF76KAcpjPGTOoTTEDrJ9cpjj7zTjSii807/if5H+5mgRl/EGaFyBolV3C29tfdfRc
PsnnlqAhOZmCcrZUR2Ao0eJlCiqT02fLtS3HovNDJBVP0HKpb4XAzlc8f0a3s2E8EV2sJOQuA+xE
itZvvOKB2gMII9Ty9f4/o6rU5Dn6XJu+dOkQ/LfqgqWOxvgdSD9j/1Ssa9JXUUHIKQrJ3y8/URCl
sFEG1tih5iTwFMUV7ZvLdn2JPONjZroHuKLFREQWRnn5Om16rBLQR1Iyd6j6i6LjCuwkANKvkXi/
dU2ivFpxPjDZf3U0tQtiEZ7AcfZaXiGIgm3G/jQORlzSZBDObDc2Zr9s0pAWnXGduJRC1QkHKTJm
TXqR22DyqzGpyf+tn96xFBldBOm1y+dxJd+IhCYvYvrzt/brM4YSuVkxdZRqcb4YzuwRhYqLRBRK
JWYQL7xFwjDsLTwiW79mKCwPtE1PYtthAWRf/UsymqWBVXivZvgdfiNEzItepWhbkxNkilTqo/Ap
IyOmO2CRw7PUUK1R4TheNto1zJQeTcBO3xZYUYj3BR9+/k2jYX+AO05+LXNh1MMUs+b8JC3nCdHc
BzQsMsMHDkmdUxlVT+KuRMwR7L9eYlu+wEgcHAIyrusdZPcCEyaYTeTJ5SKoSFMMhl2OE3Er7/Q3
ym2yt2/lZjsxkDTiSoqsE2K2LxfE9kIb5zWYz0DFWYJ2e6rqbBvhbTUMPczIkV/c8/FgC7UelrkI
BHyv5u319MW6v6WOWW5bYVxxW2H35rDRE8BZrK7DsrGi/aPBTaSN7sUNt06VYMfsbpiiSE1hfglc
HSLEnvb1IwXdBxljZ0Q9QKNIMhCH/oSKXoCUnj4O4kEMWj1X/qPvxmdH3WS35DPUbd6L1TWpgRf+
R+M2kLhvi/jJomQYxrx4L/3uZVEVr3WFGKyH5cIgx4mlFxm+uxs//0cafk4M8SaUkxJOMBgkUfQi
jEOTmvdp480wyd4edaaR2aQA97t58+HdcYGwMdav1aWTaO+U6QEP4isTBW73iiKL2nj9wN24QJ7N
dWlV3iXfFVDR3oH47aFm0Z6XE+0KGDrhgzlQg7d9sTWDQ/TUP53FmLe232iCb40l2tI/GJSfv5h2
Bk4xi50LrUU4vjhAPUzfBqSQlLmHBfO0vLYCilQibAkRdijDQR23Pv7TrfIisso7dP1+f9N4f2E3
0Yw17TqeDw0hJiBxJc8SzJf31AxQcqMZcMdtqpLqIFZWLxQzTBmtW12/cGe0ciLo4/ZNPlD/hEbh
RIb7v+qVDsK0h+2WDzjIA1rIDssN8GG26zKLNvPEY/yN5HbXG9XeuOgI/WgRYDCtnOGDGHzlttvQ
UGthwOti8BkpqIGheXE74Bm8rAoVIxcdxm/A3pPdvcNJZftk/UisKsD95aCWz4MmaWdJMgb0Iaqj
FtbQYw11R0EW51ZZxR9AZzejhaQETstABPaVOc3vrz6FDMISTYFH9aquGmiH3KGI3xfbRZbahoxu
DUoPJeyWhDvi9eo7GbpD4sZX6HbFh2eTOuuDMBUlp05xOKsq8rN7/ICLH75KHHdAkMJYtVOk4fuu
QROB6aLzhsTc69ust7cMgG5Ne8Zn9onTxp+LSUUMJt7ArYzPglU1yRevnZWEVa1TAFhvORANuZv+
P5HoTph6D6sV7jqlRTqhCkfQ/oKjDiyjGVRYVBLNlMUc2UqXM2eE/Ec88CTVfGjKfb9jAe6oze5q
sfvgux3ca+SYwDVYUBb1usrRZaHG77JFwiwgKBQceV40NbqKaZd5LPkhbU8cnoSG8S3cFMPGUqdh
BALG9MBdqJgEUTII+gTzMF9qFdabs1Ahk7KNLTDhk25NQ6RZ5gIlAfZoM28EzDH/sjBbczvtVjhU
NtbFkOJxisNSP2sZlkvTU5kRs8ngAUshQp/CLa0JKW/DlVKCzpmDgEtruddyjoV2PZ6ATvtSxOd/
RYz9RO3Qi8bDdHeo0lRLT9e2xQwr5XJs21wWcKzJzedPK1hgD3UhJlTD79AF4JiL0SagAmC+vCFF
Sn1iwClIFuoOnTfBsyhRhEuvDkxLc/iPm3xqeX64eOnP95cFc+LMo7OjAQB046sXqXo7Prk/wJjb
MHxpvRG00eUdzPUL+6vwxNGNao/Q9TiDWe2TcAxJkZi3bwqRfH2WXOBsZ7ogFWrrXKLBeN7KJgGP
ejh/EZFndYM6z8s/V/64kGv6PrIMFX6kZfeIXzAySnw9t8g5hLWRbwl4UDwVcFJL+luOolCFtEwi
WmX/r8kW3UIXUkUTFR2jMhLrbbXFXkoyy6zXekLozU+M7i9/ilMgaWZk3yYYtmPg66aNburEUIWN
ZCCbxJDs2NOrIFcze8nOHK3Nidq4W7l3wthNxiNx87H09uq1RAP/Jai3F3ZuzFuiYQFrOH5lRu+z
Fty6FXx6J/sd4faGhqPOyms2XV67eVGHr4iAnDgq8/g8FLYQLqZf8rvXLYzR9i7TbsrcTbDNL7KP
qGsZO6OFJOpOg53m5sgX8MXY+9/ItytR22JKOnT/iB/zaaMaibiPkktnZ/c64dHmf0NeKSF2lDgx
usdIx4IJoJeFrm20Rr5yLY6Qor/qH0b6oeW4lQ3BjX1w7QBuqVQNgallKvFQJgDpoc+nu6kR0XFq
Xt0rarsLHUPQnCHCGvJwCUcnkPUzqBoJgtz07noOuykBNsZMUgMumeCi9FZTlhA2406Ivh24CF/n
/NKY5y5vcIUdpYSwARV8WD3P0g/vTP9ApWFCUHhSB9EM9QXZa5JpjolVjVYBW0KT8KF7hLGOBUlJ
SzNajgRE42RApZeyRi2rxbTlEhgeAKsSo4PxLtk2GpzcxL0PWe/w1A3ot+4byboU3y3oPIWTsQ6l
AtdBx3EO0N76CtdyzOco6v7h8qE/rY8RjsZeJFb2tSoA7O1RrbYJfRBrzzvXnjv2JCosASyESIVy
cc8bz0mcMk589aSgx8feimy8Xt1hPkrrY0ekZ7Bkpq7iaARJIro7lnBUpnv8aWVGoaQJLA7RWgBW
cnhFNQnrworc3gY6rux7W2sUa/Ce5epFt2DZHqo6D+C5R36+scuZXhGZK/fZoWquFqUrm0iAWpvP
15Xe5vhXUNttVFVMXO3I1PKQLzWuhoMOh8cv/i7jYPSLMO3cb14XRZW1d9iBEYKkMUgJWodr6ypO
mZiEbNCl0EQur3aAtjDrQZyJirs+HCthc9L3LL6mgS4+VLF8fZnyw1XX4QhN4vOSqt8aj2bJmmk/
6TW3YmY/Z/wZMiE61ra1/br3p0YCw4GSRiubXbmVvkcQKbMOaYB6UOAj55QRGqZvaBJHlsyBbp4q
L+Tj+eXYtU75ZXIUEzluLUi/ufohTfdXNQ+9HzBGGDuICubqgX8GssGPFxDRFE4CEv4OcXT9ODfu
ZBVOCa7Duba8bal1LeAYqSW69kcDazHHj19wBsrgKtRu3B/whhqTHixMyomIkzrhOVVgawRgFQFQ
M5GLdf0ZaopHSTp1MD9vsTy4QZB/eu1KWU0+Wy0FJEjdFDIiHZDApkgGQZuIG7NmRoNQFA77Lg9U
67HP/P98yld3uoc/z7kKRjfrLgnc7DYdmWaTOUsu8OLdbCyURros8xesSvxolxp2I13tSXZu0306
emncF7bDOELmqajg+pz/oPF6c2OamgUoCUNyP8killZ01IrRCTUNezdSnZK1yt6epm1m1+Ke/mwd
vPpheMjBfGaG3m3Ai3EOY6SwFYQS3Jjgxt8UwTzNgliwYdDkgan2MRv9gFhcKgS1w/L/8rSpQYwE
uJdAD9ILrH5lw2g5jDlSoxEgyZFW3QCSZGGVxgMzJC4/o+CC0pEbnStnAjE6CcnVErClnYdnJXn1
7mQ+EXoq/XbWoEFqSksH53yDSSkzJ31bxv/hSB/nRCrRQjuEOUNsvBBeryWyk+cOGYLh7/GcB6rh
km/v+Q6RE58K6W0NQKOfscumS4gyi8T7Z7jNALMMSw8PTRUe90bOKYYqwl6jrS6LspmN0uUm0sn+
X1EAx0xiLNZR0sdQL+GbSjTzMdiJEC/Z1qPORHUpcN3CotxtoSips0XNXvT8G9jmXaJN2J4g+66L
6L7bJmaeGSS+mRORDWzhYfcx/jQzovGcEIe81+IciBKgdXESUzT5vFjmZcrYP8lTR9f1+wqROK1/
p1HszDy0+CSM3CqKRVd06dkh2YKWC7OqENWlQ3KCZDD0kTrAE1keUQreWnMiZjgSF98k82ZSSyZw
YKDo6nRt8UjTSvp3CpM0Xf6xnwrQHpmPgnhNTFA09XXeA+9Q576xkg0JyTNJWFX4m4xMgibu5GRX
TBcMpO5fi6Ir50G/dG9fIUfTvwrDiuKgrZW/lUETZZuWyFeBgrFJ2H4uTx0szSP7mPls1ie4y+qN
3JYwMUu9zXcmsBF5X1QmYMBXEUQd7V02gOoR+sq6mirHGYh21ncvpSFlwW3fP6XKYYewXFqdhr8J
wJMlmcoiIcDqu/gR1AthEsZcIXbqwhssJRy/0xuKnIGztQt6Iw+Rjv+uZLcWTc0XSTXHmoKA98Y5
v/5GshLkU5Phy9gd+EInXPNCIk87yInsijijEOVFYdXqyKMZoy9/i1LPVxymQRJKDeYtz/fA1IbE
i7VDcKRJB2C1W55fkMoMqT9uzxUgyza/6kZcbPJ7BLhI/NGYj5A9bmHlfRD2nC+f0z1ysGcJDG/J
pbVAR3eAumCzP1f/AgaAkkM9feEpM1xzQMGWomoA2L3xmJFoByj9jENeRHpkkzjtoxSpcXmW0aaZ
Q5UIgqAGVb0Vs3KIh7iL4xdtIujuLEEI3iT47umiFzWNgUO4DFJPz4O7jAtDJRcUR7av4k2AUcWN
1ylhKz41r8uACELQ5v9VqPLi3V+U+1KZuW0gQoiTOuH9GoZJgVwPG46Os2KhKoYg21vqLi4Ki4Fk
ECQ5ngupxcJFQwWmUjUqbZWgId2BrtNU4z9PSM0RAUuTgtxMtfFM+tBXG7xD+kqnlvdeiSJa/Rc4
CTk6eJjIvHWQBRVpLcu1Jm4xm2lYDDw6a4ZPd4fqgZSj7qZM3tBHvzPwnzRERbDwYBy9lukY2t5t
3O6BCJeRzChfrCHm2UmbD7pArtzI5fO6eiXBCRWby3dpIQwEUR+1jqueQxHBkd77c3qLQE3wF7Bb
EUlL/QQMiBCsaqEkjo/w4bgeONV3BHNHXjGe2C1zFr75qg7BcmNgOqyhK+TY0BSEeLq26MkheJmE
P94tUpYkfZlPF+R7Btw8DGoXvavhTK/AY1KRNuDFYY4wpTxsH2F3ENZCTBHqJYO8RxA0bbTnPhZj
Jx+gQKbEC8CvcgyItvjnVNeVyaMXZkQam/bi2RyTa09Nm3p81mZMISv4r0wOpSJ4bD3Ug9kGkx3Q
QJSEzDp4PP2DdEQB+Ofi8sZJlPwbGPiIpF32Qy8jydvfK4KOfyoAsMWv+M9zwv5NSmkQr6Xl50Qn
ZZkpYLPDZp+ALcdKFcyR2MG52OiGd79nFMPfyEYVb0LZnSEJXCqva9ohVCx4MO4d/MK0eBKsPiWc
UppD7rO2TGDXUsf8m+2ZfzLhrxDkhDfNgSESLGJrxkz+ngf9R9xhE9iV3WNuhqwWXtsBVuz6NLtT
FPmUeUEZCQJPstTUwpMsGt5rikxpj4e6YmHbV1Wmz7bf3c3sVTdX3Kj/ZOo952nD4UBymnrglkOv
n3k2WWEb4mSvFPkquQ4XVCMV0ZmXnTmyklr9rBSHo5x5Cb9/8gU3HpxYrDhJdINAJvel4crMhwrh
mNtmqvcVcB2lIyKrJO5UQ2ZyDs8rQG5bMXrIn+Lx0aAakIxAEJlGi4ECj0Yx1lRAfMvVKKlBmWhK
gDgVoKPWBY/eKIvm7VY0f0Bw8v3gjbphJwOKp2godvFNPkLHI7TZZymVSUeOVh2j7ejDHczvqL+W
txmhNu9SQ8T5snOuGIbIPDjeIpZvfywP9CBl8KIFqMVAI9JVv2DTqBOYYTH5967ALTek96WGeGmO
5clBDQnfr9O4lSWeLZWunORCHejpzz2/w3NaWK1DJ2t0fgZCV1G5YTnesZYM9rD6DZOy2JflALkW
bpsVCtcce3YR4jNL1A3f9M6lRJUSD4xTyEGhbdndH6hzL6u4H1Ct5u0IsBYvvE7LOintAS3vAOLf
wQMyAnD2nwhZ6WVQZ9SXDE0tUbR55IuhVqZgbN+WGe9WRL4mib3XN8It+pJdaWOjww/IaQ/Wnaq5
ZD3vX/+VCZnlALub5TbyfCLHMmNCAflniRQfA4QEH7W5SYuEFHiww7Yim+ATym67ue57FqFgUm/R
UAeuJn7w02BomSFj7AW7xAOnBZrTu5kcWun9+TVnmR66NdMemLhKA7rOc51D6utuWWYuTAZ2M3zp
qv/dwH+uSz9jJ/8MJW3xIcdYcFDfBkzCd6xMtNh8PG1peYDvTuy5p1Yo6r4eWGhECBYyHyYN9eEs
GGzQ0JLEY5AonYQ51fqkk83smh9faV7Dshq4YLGZgzKaETBr2W6xlOC6JrCRXrkP1IeNoorNlLeu
xP1n5YIfheR3zM7n3twQQ2+5UPjjQSyyvsT4sg9pJwBcPmknuREaXKUz7sjN3mHGcxK/CUBE4OGF
CeL5HenaenFNdoVc0fGGOqDMumenXf2HnIKxhNB0IT4D2LcOybE2hzxo4AAH7iIz2rTC/nWh4wuA
/qw0YqOwmOZTytChFM6FDhgX0I0v7ZlzxQs5dTPThR5INKoTNXJOrwYpStXkbxvT3PpuyWvaVVy+
R2SgySb1tp0CbdY5Pkd/4JASvGiET4Q+0jPr+3gG8NTDQG/AbZxbDAESgdH19CG7fzqUHmApvGLj
vRgyydWiRr+ReTFgjB5yoESpk8n3kad10TCv5VNpTTWgyXvU4ClJHYsN+8x7IZrcRtQRY27PBTIZ
cTFEP8frGGs8tWgA3htbtOpRzIqHjrBCwlBTZ61lUlrePNf/2RvEIg9Q2P+tgBqEP8WMZmS552k9
QCKnKWdx4ihhH119lhVdNlVEMIX6UzXkJWdF2xoyecUIM2ZkMENIuBp7HgjGhNT1gQyCBDr93YWO
vGZgb5H0khnCzF0U+IW0TlYOqKn3GvFBw2Q9rF+qGbQKjrWBfChB95jJzgUuWT45vTbesyGYr1DI
AHm65q3HFy8PIzCSeS/ontCv8UbB/qM0KEJm1ul7/v5ASnfzCWayQgMXa+vNeYEifcZeYStMl8Qx
LrtQKxOJ6tngMlyWq0XM/d+0ZXJHxzYF59DX396Gu6s5Gnz3Wxjo3j05Iklj+nXh5qubZTijAMcI
JsMiykO3UHWAvnDZLqGYryK7jJjxUtAHLcouvrcszqa8qRXA/462joHu//lZeJ72HRpxN0q6LTey
8sYxRue3lxaJKsxImBbC3sI5w/mV+X3+mKolHmelhCZ0zjKiumh9E1YMlsMkCpw8QQpFpOkXBUQ4
avrfkaJXLcKVxVAtcwD1cUOhH6QdhWeZFK2pHXUxGYa6erTb3wlAP/ViGN4Dc5q8s30oDHC69YF1
XIKRqQPD6dzSeYBkQuAY/+J7F+/k/UpxpssllFXRAiL6EeJdFaSCWoSpejuDN0xz+7pttWlzwbmZ
6S081JgL3DX1ZwhSBa+jLATuFVO0o6dlsH4IGRj8Yk3okpShpa+3PQfzwnNMMdn/HxA/I+ZZRK3j
r6uyEJUYe74qJErqXWWVWXmwpbVq9EpPy4I2r7O4xox9xNXQt/y/qJtbv8Nuza5PKgFZkydznGRb
JsH+e5U9Yx+qOf2PcW8iHdRGJYs8GrXTf0JSBQn/3LbQ1+E69bTUOqcpldLPCfho6envNBZ3m9W8
WTAU1cqKeZhXp3OjrDlkAyT3qY6186ouCNYJla+hVgsHFySV3aEHtWtnzuBgt/XPMgwBGnFzoaNh
GVp2yJo9O9wbe7ciDyTg0cktjWH6S3stXjou5DfDQEp32tZY+kTE954P6fMsKIE4gvSLbWTUBqNP
EMjtPXeej9QwE23WBpUkgOxQ+sTUQgWaVZL0+LPxM+ZJI8jdA+FBW4z6V1ITG/WzmGN4EqMHGHPu
0orf5Jpxm35hdfLwzRgliSFLHMNfpaavFbX9UJWkGkNDfhJCk3rB8/ukojWSDJT/55JpxNXQH0ZJ
gYg2oHCtm18/GOQoE50k4G6OzzMbiKCmqPnlKayTOZglIlzdDRvggoiGvPT/QMFHGkV0ctig6156
xHJtTDNqhT5yX9SEWmlMxqZ272duZA77DpAPmki+4zq/dhPu8n3VjkKAAWffc8Yic7D+WQWFUQEV
E7oXB5+SfhnRRgPj0CbB1NpbXOkQR7CrYjaWTJ1MoHTdYcvAKOgudSOs2ti9NqkavYlqdkIa8eOf
gtwSxAgTyPnDGqNiPGc1O9DJ2CB2s7obhnDm4tGB5sO9KV2OshN77Bg1uTYBqecD5Y4gJQx1KWA3
wXNtQlCxk0RSeC12+PDdtieLU7B4z1wSdCYa7LpTRoPG78ghx1FLlwHiSUcT68YdSeTBgY3e580V
oHOkFJXuPnI+EkaGWPoEIe4KE7eVV3Qn2jP/o//zKQ9T/KaXA7B2fX0PUC2rd4ScklV7hNJiqaX1
MPg+LI2j1/YznvAVX/0J4Wg/+BgrQwvuYVEByeQB8VO4HV3BFZXdB3Bs34bXu9cEX1SRUDqCL9bu
QRNZw90KHol8Ik7cyta9fZY4EA08doeq3ZGMk5KCFC8lw1bCkrwaqLQxfKY73lqwoH4WPcO8LF9t
dMnKmXFCF4zEiK3PA/iuo0K1BFKBCWGTzd1EVyQAopX3JTYjJqyiYCKRRWqjcbwgGd5vpz/Uoyra
EhHe98fOCY80S41j8nYSdCH0RzQ2ADiJwnSdzygTTjojrpf0rEvF7m+73RjLiipsQDCUypWCBC1R
hz4SIHQNLxI5ZUyj7So2XT/TsCJvNTxANvpDz3Uhv6pT+wJNS51eYoI5K3nd/8FmPT0oQZynOgZ5
SkKGeAoqhl0+sdkBtDZJ8KLxXD3FqkGzq4pR6b7Y3rjQOtq73ADwfDBzIlMFUawTV5ZBNcO4qXz0
O3a2M5yOuKPbR/ioeTySyqcA976GuLTDgOcxLFYJUX/Fk5QIlk/jPGCzLOu1x9oorMqVMDvWIt6x
sRdZvBM4lyS8tj62n33eI1mea/0S69H1ZdnKZ1N2GMBLtP6gj7exae83MGfCziD+nUm59XfZ/CY3
TeQUBAQraaMwQI2BAJScSeA9uFkh9qurnT5SYolAa2p1WAsjcEIVElvx2prr9KxTrA8fO4u82vkM
oiG9us1gkCCposgOYVPxdsBGCWywRWcJOk9X5WkUb436XZvTJAAHRfn+yrmlG0/3tlzs63Shd7r1
fdmydPZM7E7TvRdsGdQrPmXGbXmJ7VWBqyZsEbTeJ93fmJoISjJ9XtHuUE7Hpwd7hSuMk/+FfLTB
KmuA25EsHIEUZLB9SecKdiuW23N82lCnyclsKJDj0y8qEPprn/yFhn2uMFscKOk5Dpx3GCRiaKkP
O3lTxWEob4khHOCp1ONIiSf1OCgUzwU5yppSM1bs0UtWl+Fai4ZZcnt9c00s6qNMZK1mLWjxH9OV
LlU6SwLurL/Yr1MDNThnMmB9CIO1PxWWo39YFn9NQJ6K238BrPANoIG0by31o3hA3imz8darbroL
uCFth/T/1NZAEzgG8eUTVKEbTPZ/v+PD7925YNmPYdTkLJEiRRz3Mci9KOh0UyGiQt1g0Yy5K4LF
IC319PmJ/yTHFTbozidyCPE1NmX0SZWQI7QHW27kQJjGaj0M8Krar72GKz3NsntlpxBIF1VDHmNx
14scg9V5bEgjOWR6Ip5fsphJxfOvmDUnPOKjZR0ThaJHxcIhkxNdvMhhf3DJ2Tbevrw+37V5JIiw
Ev2xzFK4Yx9mPpBiahq9FJgpImGJFMnfHD0tTwWmrOAJzWr0MRfdnjDmYMOEJqQL+EKcJ7ZkJKpI
Jj9wu7l7q0OLJGSsXjW3c2IMU2S46/jYGrgxlFPl979/BA9M1dVdTARen6wvQOAuCPCxUf6kpH2I
ejTQ+a2ARTd0GUZ4tV0mgiYLlVDNAieIc6O75+LTBzvHFfDkI2e0zg3IxvEHZ/IIiX7ekFInGkdw
/dMO0CamKQUhl4Xis9A2dnLiS7rOaL8oWDI/9aCilHTqL/J7nBqNKJBfETQ80Q2/CNA7Nu7i2z0M
SI38ZYsm3Thk4Y6TS0v5/GcFfhXX43KufW+AsJe3zl9H5zrn0Qf/iR73L1jcPilcWcqGBLNTA3Le
96SiA3dNlPHFjbBYoPpqbvvHQ1y6Dtq7Gt+j5ENs6My5efzAKBa8saYt+h2dGtiC2tUf3DlS8yfz
X9o3vtdqkET3dNSfRGSetccX3r2C0RRyNK9QwGFXIyH5JCfeBX4EacXjmeqs/WgJ1sBGo1JYQtVv
SoojvdYRZklQmAcu2+8U8j78Be+XADMWvXQjhA+kBBP6q8OP43WB2LkFuxdeEKBHIGOiuy0ut+X7
otIVgAhK/KElL/duB9CUHYGG4vLJGNkGU6GV6T2YJ+AyaCJCCzlU0qrUeR59X7gx3OnkMbyTovfS
QjohKeRe3K3hlomVS9h8zOux58SH7CSQ8zs3isqZrigkoIhj4LOAeUfOHXAQTeimJGndTtZJqze2
2eM5TOxBnl7rwegfOLlDOsuRXoWuOo+KBHuYKGTW9pSUe/QEWNFHbrMO8uamqc2J7S0Pz1OxMCH2
qbZOLIubRUO0Ug0yC2nyrEIBJnvfGFep155Y5bs0d/yGEHYBZUmDHtmvVGuT8Du+QugnLtOO82Pl
07vDIRO/jy6NDTou/Entr5recpa3ZYeVwgcRoykPqAhFKxQCN5fJ+vWHhlnsbIGwwCte3pJcURdZ
+eGhzQvaBQgA/2FvmMSah7b/h64cmaiGWlMnLxpyB98WFLYc3t6vRKO/jAj4H+3S69zBlU0D47Fv
AR26ZFIQOZdFSmyh0DGNGPHJvIV9fG3wF3Aj1l6w4jw7Zjnrub48TitO/eHUFllMDzbHmjDSxTXr
1KV873fhhijcG0owSwvpvaDczYaCg6qLZmh3YhtIQfd9MAHFROYjn4hBWR2NxRKLaNz6ZZrTA9uq
mVKo2Xs1IFbizlKaNR24s2NCaJ0KYUrmrTrFPerM2KdSlg8GyhAoXzBsxs6Y8GR90gIyccoQ21JP
h9D/UYn/LjTPL7W+Q1wbYWmtsZiXTG50jFYm7nilQdPPbD4htz0j7pvit/uQGWjprK9g6tWL0O5p
aKqudYQSk8WMAV5tnivtsrW4FKBoVsB5oACei5rfw46colKXRbRjZH5LPnVVlRity39ZinPnqXGU
XOnWYFuJfigd259lWPAfTEi66OsKMGh3jFktJvQ+Xyl4Yp2k5HAmuLIwD+dsvA/u4qzahlqR1z8X
FrrX3Onzx676NWc095ZIxr05vkpUorJSagaRhPBUfiFG0wNJHgroLfK2IdlYTTCOBMwA0VeKmgzC
TaXdyk7cRrXXPNV6UpX0kMIshIT6M2urwkoVlZHovTnxfaRxKX3SloNR5zNnLNKjSyN0ezPE5MvW
pCPJOMp9lRMB6F+S84i320mo7BAiM+iVHAbx7UCjyDJppWzZny36JAG4vMKzF9ItIrPhBWokUUQ+
LcEoeqclIW5pdmBKTT9mzoK/kXiwNdHkojbm+HEeH4SOIBeS+cl6fqoNcfWyft+oP0fZ/NbSRA74
00f/eA9KZo1xwPNlZsZNbpvtmblP1QTXKm6jOOnR9xfh9VUyjckkd7E+LQTVPpVbK3dFqAAETtiB
hmpg25FcaF89j+x0JrIRa7TfwOWKL2K0scB+REuVeEMciXvK2hhjtGrVi74d1HrQIB2j8ERg5EjO
4IT9ldApplcOZd0LCjs89IORMKtjwY/ew1GeRQZs9uOQaV4PgcL/HeC5SzA4+8SLHystidO2DVBN
rt+fWsq6AzgRzJ4b/aJpBZvyTfjOpzq9deAVz/m2if0W0WVS4XA7vlmDC/STjQ+lzzAgfshAEHXT
EAhaffTuLf8E6zGRN1dP0Yxou7n89qWowAMgUtqe0CMvq6VssT0nM4t3xADVMqpYJ77Ozb49OMd2
S7nWthMj+ZtQC4ih45bubE5uO0JyOP4qYU9vWAkRJwZWNlppoNK6Sq5+fDksNpcaINnk9WrCLJt9
/tZ+q//649aYGqtfOXHNTu12jG84Eicfu3iN5+ogzK/B0an2LzI8aZdIFNigiqvAdD4pc2Coy5Pz
dxo0aA1DN8K64TBJybDNB1SpieJtsHfQ69TTaQqko20v/ejUo16iD6+JLgLV87HFUXVJ0zWX/gwv
Ef5MYizJbOkCER80uCAOKm+nayE1foq2y/ShH9+sQ3wo4veeFtRNbW7aOvIPUW6mW+SJTaLKyj1B
JBKb1Fp5xNoX5M0hewfEFm9h216OkMRMXuOf11icDWmYnMFUMRRSsIgHClcIQzEc14h0JSmSSFL+
Z0nD6lkpHLHeysM7E5W4KTwGLskg/jcDjhESDYJABzAP0vCeZer4Bkd19XWA38LsLPUluMcwe8Ih
LFclJkdbK7bWUMvI0i0m/59O+1uDAHXWNa5b0tpeAPNp+r3FlBl9+adiKblFErPSYa77lIz4aLIg
0yuTqY8H4Gs93YYmaYYB7cIquNxOU8hbPArwdd7rlhZrmkUC/NakM5ueJjeWqHVZl98sehceKxpk
izyOPa1pokd31lk2Sv+ZaWHyukbVLPq2JqTdXtfkWz0St9fj0lRH6WS6+EuM4SCHjl8ht2N6/hJM
4MFjSPk5YNXMJA4oLxF7d3EgQlH3oMroshZPS0BdNER0xVDHlp55u4jOKpL5laEOaQ8qE8slaqXT
YRkEPqL6HfrB3tGfAQdovIGSE2NgD7/vZrRzWHHZp/hGdqiWS+o5lDoZMc1hggwykEAHgT/PmRw+
NKpW8SVjlUeQHpfzJmZTe6vfrrSS/9KCXg5UounBFlVWZahJJ0EiDBJvt8O4f4bMa0ZjkQC11lCQ
yf0/4dv3jrEFk2rUMtIJ6KYZDY13SMhiwGn3qQy3U1FyvjpXXgKZsDpr3Dxg07EsTm4dWf3J87ZL
yA9/HWp+Ze7L6fxeFfMGcpk5t2B2LbMluFFPxmpUx0Zm4qHgFzJyGBm0/0fiQZx/bW31ZEVuJyVW
laNRA424z3D+Hed7td5ZC9Vsybc7FIG8gz6gjgJ/A3bKDADvf/By8nYxKMZhr/xVFDpiOPbFnwf4
ENiTxMwQ3Kiu0KN+l2Ixt2kO0x8Fe9vu6KUk4ZkGi+Nf4cMqtDBkXbeygz/FyI50kipbHiJfLqRM
Tn0MQEz9x92CgX7NEJsycP1s+2U94a+YdwB/HdtwgH4K+QEp37eE8GbtQIOawkwKjVlZ+pS4RA6Z
ASB6c6txEK/+a1/PYXT9naeUoJ4wfxaFDvh/v3XK/ngpX6llt97TkHe+DHNN5Srmeg3mRO6u7Hl/
U/as6yN/M11zgV5hhYA9Q+mLTHWRCm1R6r8N+/a8taoMmcEtZkJ5Im1IHBcCVffJ5d34ox5QOd8e
0m1KIbNn4lqhgH+4wcfVZtUHg45tMTsqfeMf2RCV2N6rQlYeKwtX+GNkMjO6oprPjGQksG/pazw8
hVAXThIMrwdJNGorCNARb7WmTktZ8fUvR1a6DZZIoqIak96ztXs8rG+MeyWve6Sb4Rr/G5hDaOei
g/24cndYxjJFO0ewCDequ3puAeTx2RacLWhsPzXGECqlj167r41OeztlcD0Luw+oqwbY36Z9x3cb
Ib0SU5JZe43YxPpSQtsVGlRhnyc6VQAtEdx1wzHPCJTIWJXYyyBTynncuwQhbRup8xs5MnROQM2O
LBbNw1EW/9NpUF8rF4nOykPq97SgXl+66E3NUlWNiOD3JT0hi47iJ9nEg8XLxyr6g099EvWfo3Yb
Uu0//dY7uK/PvQofkUUljtEs/K6qjlXBsUTke8xyPLN5eJk1+pPanmEr2eAh6yChNaswQNSmO5Jr
OXF/VZ3qAcRHxsvfJNRtBx1ReHeRRITSc4G8VDo9QGDonK72OTdxLlgC/ZVAlJ1zbMpdUi039bIK
fM85t8MifjI1YFA7Hso350uRJbdvuUm4y1nxMV2TCiCCbnrKPox2MQMVMn973hIiSzPInPtCagsb
udg9ivtEXql0CXMlg5uZzoUYb4V0KF1FmNeKglCAuA9Peooc1rBUl5G8ALm0Jcwb3FcNK/meERAc
naK8uJ7L1+g9DPnh0VVuXcewY2eOA7I3ao6UGcg7x8QTwYnbKZzZl8kmLmyPyGJ4Yyya4uYTGgXl
H8r+02cpuRTL4TXqjLeniKesjGMFeXo926vQcSBNLVFsgBZDXYOGKeHrGmS8MpfW1aNqBJihNvYZ
cyM1Z9PJ1mD0oqEWIaKTrVLBTKbxKNWedl2FA8DKhdolanklQHMrrV6aBg1J2iD64XAAtmCJjni5
2Akd8jyLxTHCX7cDxwp94Iv07B/2KIPd+MG9KszjfR9S11aawgDWDAseGJ3wCvsO/xDtXGjseLyP
58c+wgGbf71IS9iQvQMjbWNqJm36RcPo8hsSgmAAuHmW1TY9bUwlF+qzHuPeS5vQELY6rpmdNJmj
zli9+I81LIAzCI8HqQFDyKHbGo1rW7245QKGsm1G65rVRUDlUSxN7K75grK797aT45SLCBZiwOJU
JcRsk+OuBEKC84yL2K+B2H4vwMkzQsktkhYLW4+OXy/hP+hYhCYZVDsUmg4ghYEEGCPk6fhZLY+n
76AlRkK7fi5Bt/Iu/QKMIsCDjx6aT/UUnMHVIpyQNbpAPs+Pngb2QUX0jC8DH8bHs3XUuvKdeEFG
qIicMqeqbvNcK5dLZRhZlQpiLsTyx1OheDZWPKDsXX4MTowZspOHwdWhZ/jfXPOqleSCfLOV2S1b
mvYJNycOaaHNwwxHE0ohpsLhX033i5bHr2yV5MA8bNssTM13dJHJdwm9LFn8KGvhGp4ZaRvuxNs4
ye4GzwyAbULzapSZcAUbYDcIpbzL/vRR3c6jitFIOFZWi5VBK0vQRxdlc0JlZcOQkOxybTm2tjSu
sxv2HVGgd3ZrW0Cgu1O2mpfIMHFW7vJaUMxtSBbC4JSVUYwmphg148sYWUH34RjJwBrtVCMMR5F0
I38KGQy3bNmwIh4kFf13NM6gTcMRmd1k/6lCSbh7CydFGDf731yZ3Bvy2cpMDXPAfnRDyr55NNQt
z7cK69Qs97pTx77/eQ6KMAe9P2eO6D2yMAc8vPjgF0w/l8Lk30hoUHg103CCKJBu5797Ft3818yS
l6L6EB9A1C4egoekJ86TAhJlzXKTDhUsWbmT+GeH/cARKo7jI7IIN6DBBAJEBingpQoHWs8tddX7
TKl98cdM6EckhhSgGwf7mYMvU02GZtQhC27lZiLnpboBpMkaTcpg6NGtjSv1tYAcCIrBDmHAufP5
mRpuIW5b8o4uw+dJysSqnTAKZOjwhvYnj5gVw3MZS30b7bqYyW4BbDCIwAPSergiCZWEcJlDsv2P
KZpkw5hwWUsNkdgUxoYnopAiEQDZt+umK7r2OpGJQzofVA/jwkDm2EbTXFOw4sIrvbBAQlunO5c+
NCnZZVN/Svz5GQtIuYqPJ8Chvm9thdzvDDx6mVBnP9SOQPQvIgUkcBFUO86P9bxwKrmGsyZZ6u2Y
97y6dGYn/WXpywRS6jfABX7alx6BLUMLDsMa+ZCFPpDKhpzTOEMoC7BE6QmEwyc/OiFs1Cp2YsWi
i75trbp7BG1jczijJpOu8tNYPQ4DrwJQ9gFbsm8bWH1RpqbAsW2dSHzhOKTnT8qmrvfUIYAealca
v0kHt+ru6AkTatboByife5oR6LMaPtGnZ947xCJ0CS2BtVglXqTVdY+AaW1Mx0P1gDCu2VgvmnMf
+XFaJ2bDSr69XM0GPp65ggU4M10GfouuK8cJrNM8jptXAwm3aL2lpTi5hTELr6QL06oci4MLMbSo
Dna/TL9+hFjZUoryUv2DSRwUFjqdApXPU818iMPjRRCkp1ZzU7PFDMYbSIbWCqEHVcs8NUN/Yae1
CHvDxHJUzyMW7QdZViNhesbGrNnAuboT9oUQEeI6u+UB2iArdyUHdfquGsOfWNl7k9k/hKUv/5Zb
QJG++/o63TaBtjod3sJIq0D2MqMK8rQ7DljR3BtOWQVTqI8QBh8s3O/JZbRZtTT+SzkuzH7ZVMGe
KoFw4kbC4arj+AteM3cv092LIDrwf3M/AvTOaE146bqQEY392s0WTyjf+DmHu0jj+adsU7ssFH4Y
DjQeRVvs4tATfoR9a4Ln2OHOGVA9Re8MzhwT8X1aO2+wncKX34SchmQYmKW5JLPd2pK+ggexav38
zjsJhYOCOurUss6Klb+7jeV4z5ZZHHGaFoeHHV+ktCMH/59Dyin0/jpDPvuBOUhxt+w571BBhRk2
tef6ed7XcXOOP0V6Np/K3v7oRLcEFYnKXyeNOGDrHru4Dm0kqw1d9xl5bhzWgeVjOWDUbxlhSQrr
u0Xyy2SQpYwEqss/aJzNqnNIlOL9wsBiQZFgLNvVBUldeO+maahoFGi9Z9p/RaAIVmpW8fZzvbxR
u6PpdjSvH2Vn+0okznUO0hn4jLIrfRRk958ZvfasiZU3mHzCzVwA0RkJjOiFN18xbR5/CKUrBVVj
QT7+AU70/M1gHTvc2bVYUMzfSj5+3eKGTFqNnD9t0NzeYR64dlcDnnTbbzMrG5x8au5gUn9nIqTp
dEJ7NZlVcylQBMoGXKxxOHNr8hLACPX5VW99gJieJqgilnBI5kM9NyXkyHZkBymtImrQQ/hjbW4N
CPTURg47lLhkDs+EomzTm/KgyZWhUsCToM6N//xBROVnwwVQcyLIC2FKATcIj1nXNw7JLGp8Idxj
C7XJza1chAYfUqv7Qq0t5dkZOze3nccbLiwmTG1LDNAj3isxF6lJXGDea+eDxD/rooqMTevQuhm7
6UcxobyePMVqVgoGOV1nkW61v6IfupcM5XobjcMmUJOTiWajnps5+qLqRc5N04fjH2NcAmKAA+Qc
tEiMpbTOxmq6iDk4jxTu2+cIQtJ+1kdjFkMRS4ENx56S8xyOKiPf75J+y7FhfIe8r58/BbRrSqw8
4DtfiW55DoGZTlXJoTAWX8GZvZWEjFUO7rWT8uDcOj/P1z6PORzcktt93lOKOoYtQEkyFGKVS14z
MVaN//o0AzRE5cyiq7HO4l8ZgOgxRGlhIEcmloDS0FiC14m9g2ezw93RMndASZl7CsvFBUm8lV0O
lOdUvoFgESxseOuCovbWbEnK6C3p4VTBLDUkqN1UQPDMRjU0+CKRDK8oRTsGQiTXPSjf19kOodos
+JTnOLWR0DpYN6dbatnbHeywIlLfq37yEhJJFhn/0dOhbQfeXPpVcYZIgXswbpIGaYIGa3cJvD/Y
02XPiZLV27FrsOaEE43+oHCU5zgrdzcdiSuvEb+AZiHeWn4Bri4kmd0LqvJT8U1/pKoYOCMe2P54
NzC479M1aN02BcFG5Rq3mLTXrz2Ir8bNlG4w5JQ6WoVvipOBWQ0WcQfQMRmNMssyK8SWX8VZf/rl
eFB786wtXYEkWapLp54xPqeXVgmOOI7Gv/q1l6f/5eaRZS9bRdd24KIv959LtDGe2b8s5rEU2U86
PTXmSQpTr8GqAb1F8s93prQ3ScTI756NO9MyVvMMBVlJ2M4kDXO+HSiY+3b5yM9kEpDVcw0W2MeK
kiqPGrtLLq2xb7fgF6pntAI6SubaeYQDrhun1dwIDpQgiQBeIRjUf9F4M/rstnfMtr3kfoxNSjhE
Wiodv2dbgsebh9yUXzgFurr9gytavbVN/dUUO0QJJWiGdwO57HnsPATTB46bFCgtUqXfEWBFRe2Y
2iEPll1Q9axV3igfTG39lVUl6OAAYfz0bz4CsXVWToA4lKWkVjKHehaNz179KfwAweUo/nZVCRXA
9Qb/ZDoM/V90+3VoknSSyNvC1dLWVK3jpSJfLbQzIRT58Rt6pkmj1cs/6C+a7yGSlO3WNFFJc2u8
KvtqyqyJL0KLm5darlhaXpD84Z2cYyV30QHi7dC8c+wHNEUInMrKe/4dQlEthoujHol+iTYaTZ2c
Z6PptB6n25C91PWJC2FnDy2E3QrmLdOpij3aFpMVTTJMFh6MEK7hzhl9nJvrvx5NtyrhzLtcIdx5
pmf6jiDu+XNa22Kuol7PdlFBu2a4eeMjMRSRF6fNpVyZBxwOgb08lvaO0t+Iq+MKw7j9l30irmpa
Klg3wks4h9S9khneUT53Tw5QQNYTWo/lYP5AagY1EbeRtXzL7CwAhC5lLEdYr/B/7GhosF0vG5lE
JVSgpLDUiJGu5fwHiMD+4qCGOkjdBun/4DnjUP4oARm7GO4TH61RNl3WL3IteHbAFW+HucQIDg2n
HZ1Oqm8aiIBOi/pOQRpkGEhifnT8bXh0Yhi8wDcg/lfLu1ktiboElLHNEo7tghT2BDjgCxxfJj2x
fVYXIBz65+ZObd3x6Jhv5RhPNCRKRDkdqFSspMUbunhHt/dExan8KHodJMkDVRb9yJ6MUZNYd520
MykkwOfjWFOuIezWATkg0cb8vHPS2bvZc/YAYcZ7n5XXhpKVBpu3xaSNSbL/pNWDRYOik+kCDtEl
ewtJVxyA6bf/EnsMMmwKnKbtlPBgs13ncrI0CVWxC2St0ocuzT4AFNiHTKPntOLbzRt7v5WNBhpT
LrSL0/mooMxYIXkZupg0oZiVjj/yhhjb3rOpBW4AOd0Upc8Ew3okAN3XynP7xYoKsmxJxUxZyrz0
Gxis1EIE+HBj0kPYqty+Fh1BDlnertpWbxVwQj4c4aMN5bSgS4297oSDSECLKazs5MLg8M0DwyGW
6Z1Xqrstwl0A8T0fm8hDpva9Ew7TUBcwjG8P9I0SAXKXYdLaJYAx71eDL9OVo8Uqwmln892PXnQa
OEq+prMATNzUbWErzxo1xneBXCdbvzEZnybXcfYXzh4yaIWMSuGL/TVgH70ItpMrh3Gfpthi7eSe
14KSMReCY/mgdA+EgMuaMfLjb0J3lLD9I8TU5/0Z63pW99VYdLYr1GGfPX9qUC1t1F542MjQMtUL
Y06wpKtuSczC2QmwpCB1r2eIfkyib/3oljSilEkxvuvWzY/6IyM6UDQfHr4rN3E0boHK/ShSKEGM
63Sej+dajSjtU8IOQJBg17ayMo6LUNFI6nQzl1o1lBwCv2ZU7qm4UP4nRnSXTe9eD4JAQk37NSZg
kBbxJEPUKkMnd0SI4Od1AWat+jnJtfZ6oQmZQVI6z7G1k70FGi+RbpOT8q3NPj74+lvphKFIc+6+
eSG9FVnJwT5Kas0KfdMgLA3AN/z06a3VNXPqfcdStOwT6aeHX2lrh4DerTFlBBgbGXuqS22w04Qm
k63++sbrwbZFNBMv8R8/DxDBn8sWoC1KE9kLUWNlElKyHPTkS4pgwoDGb4j3YYKxTOCiff4Uae0D
6VvQJ4D2PS6fhgsJ7KcPwvIfBpQcHNosIpmJ7+UbS2nh6bPIypH8j8mmwpNXNwlZ+Y58znnNfhWQ
Lou36mOZIu9H/1HlLIocBdbkDpIOWw9N/71dKXt8Q7teh5Hjy3sn676NwHLqcURMV+k+IJRD9/ii
vqGD5cP8Whu0T2d3/XEMfa6L8N0MgpqaSKQhPC7tBDBPD6uVL0gOLAbGFdMbVv9ZZp2nadiWRP+m
AeIkMbkDWTBNES4XBFeCtuNtMkp8uDNyTt3JgA8vUX4cOnXtWrrdUrJlQ7AoqNgzL8mYeiOmKu3i
5KZzhY/iOntWMq0srXTwmaiX+06UQgcUfJeblfR6Um1g2/uS4Aw6fLYLtLYSK3zrm5fKobazUgJs
YoZwKLUXNrTfz+0e6mPj6FtOmMjKpZtiA3LNxT6+R+CAKS9kDmEtVy+1MqGVGehYSg/A9io0zToT
QBcyQlCxvQKzQpaduRmd8l6e9aJH2G5a+qq8zruIArAeBRJDSytfBZI7c/JFD+x3b2zSy3J1+ucO
hS7XPHyu9Kj5RuT7arDUy5vZvnQ8cD8M5GY4JFOoj2hWw9Cx1zRWRSgmoyoHrGrnH0jmpLE4oWtP
7SxhBozwqdSsMAzGURLyL+bW7/kRL/sEHGX+PBEPxVdabhJUw2+xbgnXGtk0wBG9aCJoB+tJbiow
7MCfL8QwNfZZQPc1zcgu6Nn8/vee1rPXR6j/O6/rlQvNB0WWj3qcDPzCzNdHea9GLc3I1wywlFEL
HvqhesIOd7RO+UQCNvxC5kH0I061v1ANOFxg3xfekDrHMqnIrwEGwsFkyrQK27lr3s/ZqsNorme2
+q0V5HmE7mu2O5bXxliLoN5YSLCmHKOYWyFB1fQYML1T6qg4gulotl0N/dNOsncOVSIM2MSRsOBL
OpG0TTrpiDhvFWzz6chglEvJB8pVC9Vm+6iHh/xTt5jRIL+zWWDkEPTctMT+ZsJSctsiAQ8sVty5
hLNeXxZhFX9ThevlJocXvfAHTARtLMOAWwWiRojFZPUyV9Hv+uZey+xf2/SuoT9S0Dvgo6URuAxA
JpY9jk0ATcyvLVD2dZgjsmJ6Iwxu0x5Ec5MDTuqHyiYDcEQvGBGZukuAdtx8g95SHJh96w0ghWgm
KyzPEAQfLBIpE7gRsiDBpdQrEK/TOU8/IGzuKEOKviiaJMvD0n+GxGTDhxu49Cv5hfPWnMuTLWHA
oKKs73KAIP98HrdE4UeDr19F1gu3ajfSxxe++Rj6OpX6w7mi5kmc9K2MF/4ruMu1uwgzdsKkcMOD
iKMC3m6Cnc9hi9S+/iiFpjAoB3AyvmPdXm13mc7jVKMa3S8CCXqnXknmV2x+JILN4G0c5RogNBhD
QOYbnFycQ4GdXSUqlLJ8qgQnymovF5DyJ+jhmdZuYqD3ojMWof5dne5WwTj9GE2ffF2YpDVLWtkm
h7AaqgF32OjFQ3ZJlATBdAU0CExi06pc/yQi+oH7wu6ROcONdPvT3zSJ5eQqM+7o7P7rh44ZUswY
Kh4Ed4zOfOD37oTy3++29FSem2tHDOUowhRJkyvGPzQ1zWc+eCBBEZWfth1AqIluap84CFWJFPHs
jLGuXaP6RCCvJFF2Jbb3b819+vX4USpZB9lVhueaBj/Pw9f47q6X+Ex4Zng/ZZ9ZRPTDiu0QgPOe
NwOoBP4awNXZdAdcNTydoK0vAICLRP3FoKM/99QaxrzzPCD+jLSDkuS6gf7totnltl44EFny+ApI
yB+hY++pkctgY2B7Nt2JfvOyg8jWeWkEs5wvvcYPtw5e823THX5BIeS41+9c4wNrkKadFBTmEs1A
yjt1RgtqPIrOiNL68n5EkPbBf89BEj6eNvErtYr0DLFWQXuXnQ/WO3dE/CJlCUsqOwhsQrC9JszP
HPfNMbEFAkUGznedqyjPZ0jrj6W57pB8LhRdC0slPHnSwgBVm3UjbsRp/w6RcIvJuLquje1iteLV
F4rzMyJ2mlyxDKG+TZpkfZLcqSAL27APY7hc7uwn4NJkX6z1NPLx7RK79TthU1sWnw9LPY7IcZKz
sNFd7XbyXZXTNUZQl2gkL1LwFGlXyZ5e+ttt8gZrjG47bYeQLkvzPPiohTw38GWEYWN/aQgRX8vC
gn6zMzCYe2QXzHxrugJp0/7nWlv75ycsfb1j6RC/unkMVJup3Zup4X7yKH+K/QNJILPL9iF52dG3
Y9lky0u90xS9hExfKisIaj+N1BTwEneo8Bh9fu+lVlNeIvAFiAqQim7gvnPcwRJ3durVQcuX4vi1
H8Kq7He7vMCJZq31wr4ZhljLp145BonXme9apO8psJmLbe2G3PKYEUmTL9c/cmyoHQGxcy1Z7kDx
DgpyIKbMoen6+js/K6aDAkhcNVZDpcf3NYE0CQaAOCQiQw//rmndUKlXX7UGJcBjQRbOA4+6zs00
jsEIHnZvuyZZhMEggOf8UQf0mxOLBOVlamdPBAldOmTtpv3aT8h59z+1A7i7CNNSy/bLvf7HCb1+
/jROQ4xAGE33eHqx38XQBnmAx9I6Yby8Es5Uf4OAw5phzvWH87VhIq30/23Rki6meMIJkCS7fSf9
0OiEOvyw2Vjzs5/iFxa1O3VKQeuwh3N4n2kPW7SW/snZJ2LXzVFry15raJAJsJNUlUpMH0lW++A+
IqBMrQ6z6GoTbnnj1MVmIp5FD6PkrFnwRZpnii291/cd6o+CwK6jrEBsiyZIvu2vHIRhzVwgufli
kpJWJKBnS/xAF0GGMQpceNufkGhzCs2ukwofE552LPlpDI/8N730WxMChW+tDVuaM6zQoFR9cgc0
VemEML7z4PqL4iaHsIuNDncLMHBegIzLzJnjPuJOsPGRoxAuKJp5gIXKZTs0nuAVgiyF3yGisJTE
wzUq6DXqZ5Mdfy3tH/7sPDnB/BlM9xJTWh4i3OM5AgRSuvvteLNN13CsivGIQRD2n25WhB+4ayQV
F4nutCnwdcFhlGelkViFr1Afo/Oc/jo2jKp7rPWLRBhyuivgPKPtQ6Au2x4pXngghZ5eejq+zuZv
VtYlk7W8aHynRjADgD1r+dXg7r/VWkIq/XVgYULV57N0E9aN52cMEHHe//KmgJcgks8kgkI2ssMP
R0mtgpRoHGFUapOk+vFvFy5hf182ysdmyQLEWX78s0M6bS2q0Dd381bEdLakgr+IaRicuoQkGzkW
9+3Na9M0TWTkmR8SYXezevzb46mxDYFT255IsSXLEIc3EJNP9pDEJeS0zRvCSrx9DbltCtJexyPW
GvW1u5ksWoSeZjhLBp2bFmenn7Yi3dDVzoA/JTvfoawBi7gFkSqJIhyoMVQgfCADt7evCRUH8RcL
KwZTiHCYUrCU51Cg5iVMEYWDCHpzzK4HfZbzyrrkBoaTuMcYI7RG3Jo5mZxnR3cpqLTMZeOndEs9
Xwh4TwbyT3Ff3WTBKaZrxBBx/e5XpK0bkVt0+0KRTpJb8KLV1LmrqsuDm+oBzdbMboeetpLxlAZm
6ZLUiviKiayxTFyU6Ygw9nFh1iuY888BVOTIXjbpo0RMC9hGy0ocp3tm7JrtJlF1Ro4aLmSjkm/D
QGcaED8MWcpJpCj+VOuZVFeO7XzPY4ZWi7CAuLMCMsl96bwb4glg7jBJXuIPde5bxeoKr2pYtsw+
QcjehnDtxY30S9iOauusJG5jXQKhvBqo7g6H4buQNvTb64mZvvoU9+eaHWVnRe2RHO9AyGyY4ue8
/AEciZ2kGqEE8iHRAS4/7h5i79MbkAWwQQWOXZCURwaX/WcxvfX2VwPjQ1qAx8t8E/eThyi3NhNp
vQP76kmGlDYqkuIFOexnLWdSTMtlWRjurrhEpe1/qgtXAZCdmDd75Bx7B05XiXT2YpqnaR7/2SBq
lQfHVQMakOeAgHYgRngkGZeNFeD0Mu46F28tIGw3N2VZLOxQDTybbyxrX+r01jB6WP7rOqp9eh6K
VBkupZA8O5IJ8YwhBfP6KKMXWI0nTpcnMRb9HkYupsxHY+//YLbOLzmVvyjNKxoQGoTcA7D3Enls
HdFkRWgKxv0qwacx6i8bWpAfm5oWDaDzHSr2dEG6IZCvftBjQGg4FogQ/HuVzdsKDV+yjnDPaGZ9
8HwdbE0bgtxOtz+JBYR+anQKXivVjsb/lV2rSsjyI+4yZRxZNG0pFUqtoGnaU3DBAGFs+GLExjTD
JTnFYj4lGS3jFO7DSfzO0vAii5LJJQ0aPMAec6FPKvtTa/DA7zisRAya83GUQn3W2xynaS3TqJlK
tdywvNJ45yt7Zhy2X+GXT+MRttILCr8iqwizbeXEdmQmoKRBPtpmMdtPtKZNXiWDht+mmTHL9cC/
hfAS2G2xwUoj3m1w6S6Xk1cFgikk4jrU3+7hI6jONj1ZbP1QO5CytIy5gjgZYz209EQQOKqeFB5H
pRgVjjNvPex+/40Cu+dvkQY9lgWiu4SDarWq8ZOTcJWD77YFHZEP/m+eWMe93rf1GCNokMu1BZWU
f018wbhv3DS3oLQmqrJwwmL9dsZl2o/DP3XPfeGEi8X9KcQWJ7rt3XuYJ9SJJu453I0MiOcQ/vg/
Oo6bt1IWVtbfo7iR3/S2+Dpe7kukJ4IRsHZvs4TWhlsId+60QVQRvERa0v0ceQCu0m9yhooHG8pK
LJ4kUTy/bnQ+0/eeai8VTrL1BVx6PMAG73MR3NLyudxukcLgIyqT/Qg5m9f5V6b0wIuMcg8j1YRV
8noSf7gU3m72u/gnreFvWsyZURIrB0PR6ZAVPZK2o8AQMQH5XDyC1fNfVyeEEMrs7kfsYXvEqyRL
SI6TkS/EPy4BlR81SJvZVG+9MZPuNq+/xC+9TRdFFZBurxGhl7Dx5zA208P4psU/q0h2XJVBGPf/
e5vn3XrTXBWdHVK6yJR3z52iIVMwHtMHCAUef25bmCq42qPBlCkH2PR1YDh/uTEFMU77tP23ZY46
aVz1E4/Aavwk+bgw/TMpC31JcwZGykMQ0xqgjCBRAJdMJR4gC4PVj8Evfasj8ZyjPRMKtReAuuGe
FCBWhhvjV3lw4G0It1khoMR2Hr316+fxVFUFPmzB7Vh4e77e3q4/uSPsDLzWAhz1jUaUKGsvXO+S
rMPfb+pI1/yZlR4P5S82DN+4wXepyqsGgPHB9pJ7O785u7csMWgbAtkNhml2ScVsJIvmBWplXq1l
XbArxAmWnhGI0gwGVis2dp7448CkcH4rAqjjIXJGSkIFbwK+5qDj7Dl2GCDf9mtkNujDYuxxXU5F
cVN0nKBMBsdsg6njy4Va0DDnwwgJH9UuQpdZLYZnCmQc4N4nTvEnpR/H/7cs5HlLPD0cKTF86Aqy
sW6JCfNQwruC83M0jjO6KnjS5Upx+t5OC76frX4VXwFC875DxXOb1yFlIemMLt376gGHEIdCRK8A
h7SuIlcvnohk90idsQzmZpitJvlxR8eLERIp1DIiQDyAZTt4usviChSGZxgrOLm6b/Usg36XqxL5
IiCbmuI5Aa+fqApHuNsBNjNaSyTq15QfakM2i6E+Dvmo6dHUdsTP7MPOMGr/MHFxzE5ngnhKUSjY
geMBd4Wr2GyWrSMMvnKuKYlsXvjMmLeMPwVvUuO7LhUxI9Jyb0UK4tNRN0DO17oD+wf7RFgjGlnl
YjUcILDG/4pMUa19UN8Ma/zfgDm5NVAMfuNtnaDH5sKPdAStvCOAICuF6tSgPm6ztiYGUtMObCfA
wB6+2HbxDESWmfzOvkHUjllUVF3aoz/EXHx7s9FjarQIt8SHOiFuG7tC15STQa/ncut8Q6W0uCU1
fpJwSDd8TtWjk23B9gvAg1wIDuRYZ5fLZsnQcAZJAbOwitijAARKRrzx1ELw0Zb4AwUlQqjpLnUJ
F5zhdSsQF3sLcZMDB5fjhEPe8AfMe7Cxj2tOlMpsE+ceu/+ylcFGKr99KQx7WaH58MQAX3g7z9DM
7O7acX0V+aaAyV0Rybxg2kWqGpVn2W+5f9tlR8OPPyVlnVBjdls2q6SNK2TDwGfSdUsOIMPuRzmv
vx/gnUF47fY1Oic73ad9jl81/Bsie8ltpi/s5wVmzDbOmWgz6yf4hiYXhKlZDXMrF9l8MXRoS1th
SUgzBVmxHMBHuCHTvPKE6NKxroJTZxqWBfvwGfGI/r2Nnu1IKH8q4eA2AY2tzH5NeUVCfz7wF9p2
XsXNayBJ7HPBhYZe2lMkPJPnXCzUfBJqBxGJMZw00T/ujdCRAH8MAyyc+znd8JxSYJhJnNSYSS0n
uh6ewnG8htp+LE3miCy3L7/yWgeOCaZntwLuikCTYb9xIFsdUgGKuXHY+q0Jp8vvcr/Ma0tlheS1
qXhX0yewl4X4b+6yppqQX3Jix+/IlyAZ1wskGWdqOm0d97UIBCY38wndaYZEVVUujbkQ4+ilfv4N
HhSjz0UcHY86kyHE6SJyHm9hWTzlybqln9nq62k9LWqIhCdXyBRxEzBG/k1If+2oUOifI1kGJMm2
piQnbMtGETxz/INOqJUiLSF48EFiMji39hnxzqurp1hGFMiAc6P7bkyaMEe28cJxBZEQvBtM5Lt6
5p6k+FZJUnfw9MHq2+Y9/R47kTHSYDDBRLhHIQ1lLp+7axaFm19AkufPQwddXufEIEuHUfiqu0W2
5Eh6SpWOABjf8ypxgoBMEpqie7B3PNX2Hw13sNMZ90Er6dQ1C9kBcoIxwlX6z+Gy7hAdWUio5EwW
ZRoi8SNuM1gq3iWFZIxEDX1wOtq2FH0vA/YALGXGU33Au4aZW6Ui3qTmWHqX8kA7MbC2vQu2pgzM
zAGv1VIm8kIHvVBZ9ItHISNUxA2eygMipeKd+Fbb9dyQG/HkpoOCDMybMovTPduzlu2MeKaSlYz6
k4ACDqQcHSWt39A2NdMgqEdzsbT0jMl9OPJPyU+RT0QYTJTYGwod0B5QsFwSvntaFDA2eztuUCMg
8IwWvee7oHZ1cgPkI4G5k3OJlqtF3Ukdwf+ijIvUvzO2QNZ72f/mrLPlqdPKhrZToWsSp8Ec1hK9
XlLImM3gzJwXTE9nxd2fGHISd3oWrInRa75L5aXtG9uFTdojzP0WkyKmb82McOT9VgbPOotpX/ZL
cW70/7nHhFzHS89eSAilJmXrhcN2akatxByWLo98B4sENsd72Q7bHQMKQWSZbuHHC5tIMyQ6iz32
y6LejA9qZMmp9fl8SdDzJDjTXqxvv5UaxB34hLizg9JiIOFzmtgFTn8+vWPOfuP3LoHE5mofJEUs
+PXdAtOG5avFU4JF8OdHAar5y8xvMnp6mEaQ4ZKhvDNIVN7wA7pwyxCpv743j6ElOiSwS+xbvzWT
02iKC1cGcYGmR26G/sXtn1cHpaqsgMCI2NTS8soYr6lJX76E9+GstmUM+cMyrTgUcz+JWRl22TbM
66/A1/CW0NMP8HVHC1r459LVF2XtnYhPE13nmeDmGkrWI3T9Dj+T18hreSyg15nyPfNxjIw0e2Sp
uNX2GzW8m/oMfIR09re42QPvnyGC88MqZ7oZnHe2pQbZptq1CGS5R3zfD11VgLjbnHwXdBC43VTc
S+IFyoLzdUZ1C70Q+2q2sMfZUuBX8tHR40GWlOo1Yz0irzw2cWX3y82uL4znDvnC4aUG/JsSoSoy
tUiPCCFltDxGskcqH3W/Dktmwse7WJlfTN/6b9HN73JLoE0Fnd5yvRrWUZgP4kywku8M6MHpdeQj
H/843JD1d9eyIfkk7wdtIxg+Lh+WaI4LasjpdNooDJHc2k3b2yPfgxtsPcHJWtZ6K12p4LMGUuiX
kF0b51C0VYfJGDyYi59WkVyQyo+8IQaiV7rdVrqLZgLWyLu05jrDdH1FN04/6gyDtWokDO1vM6yC
M52y9Aw5WwArcBn10MWKs8xUIrXKVk4Pz25GPCV0P/TfEnyDIvyNkaEZmd0X4WGhl+Fiw7FScg/J
OMMPC/3RWVDmzvx8dC42XPQSRzQASwmSo/1u0rf2O7qPDY3dXVR1DMBX1ForciAwajCUxxBqCNNO
dSLlD5lgvbc51sNpZdbk5IcVpXP8PyKTj5qlb3JxylLiHyZIkm6H5OzHgvO9Wi6QnA1xLJ4JcbAt
+G5v3CbNbxh5SWAtA6/n7TdHXD+aAJCVSkSwcblBqvoQ7/0Cgr/vCOzJbWfrhLYdmJXrbEAkrPdu
WP7S94WJ151vaFeaO5r+IAOOzV33wp+JfeLLiChYnZASD/RAjYXk5oW/YIuRb4Y+Xp/ibz8DwbgJ
4vMEOIgTH42H61n9rQaX4ZoOBbtgB9cX89bWBhw/feWavL4YV8fwI7YUapkW8Z+Qvf4UauBoJhDI
VoavAsowXGLirPzw/PPCu8POhVzWP2PkMnx3AC2QTYvCjRwl1j/4PtEBKkK87/PZeTgvya39t10o
sTt0e94OC9e6o/D6U5wnrS6wlsELOXZUvkhIECqWhbQIoK4f2slv5lidRbCfbRVFHFeH6Zo+F/K/
Kk3V/bMRx95UQnmYr2BgwRJAfbMQRWAcmM6dEqLIEcSlxuz48WCj1jCQWd1g+Y0hCebL8qQUs3tg
ZuVcoHK9PGKf73hKj7mID7TBcPAL9/1EeuZN7O7m5Ajagr0VghYRpDbjR5kxC3I03I06tgvm8FkN
Fib5KelkM1kaVnvsVTTUCqjBkubVyu2ajmoogoXg3xAdMIOkBXLh9il9Rp6ZWG8D0F7FujLnFClq
hxwVFBG0npXzIMEYo+3GxByVVigSboATdxaYCwJ0MubtIhs32b5ww/YI9zuL0wJmOOvczxg/P2Cs
VZbYib8trsXp9jqwWuQXhYnv8BGiV/x4k52VutThIQoz62TRpdWyMSKGqop6LYqUWEl1IyGH/n8s
VWG8P5TdisWt/p3objg9LZuHNy0mG/3vLLpPyeiLu5HIcxhdPyAProIppI2mO99xBMiHjrgHOhAZ
HlGo/Uaf0zHpx0iiY1Unwh4VgLDKIqqa9MaeZ4ah8Qb6UUlHpCNnabVDyvwM1EbwPdfF1qfFHg1p
6Zgy7qBmNeJ4bRC3Dnb9/eAfU4ZR+MYOZg7Y5nnpb5x0fXoep1Fz3p3xIPR5sw87y7byfhh6g63U
PkjC60iQgDY0R0GobuaphwP7dLRl0FjkYQXVVA2xYAlPkkDs3eUa0RuSQ1pe973O5tKO/cTLpwH1
4M+3AQDaTmDrg16kkqfPiqR1nv5kwNsM7ntPOP6Ghv/zdOo8jlfRIpxoPgJZIZ3NtJFdyXc/bfbS
iYs6fWclehKSl6IvbRh9LDDiD2sUPycFyfsJxYyHBz2H/bD6l0+gmCvJ+F3bn/xGGvlfto9iWX3y
Z9Fo2CUws6Ke1pqUOhstXq7Ok8HoDIxolMbN26LhLbAeb+pVmxPD6YsYaP7WQjWFTLw9OJ0miJ/v
8qNEGEhWDV3SqnXLqAcBi6rOSySb4AKRPQKKKbB7jNhK422jj3ZIoTgWNGnGH2gXd52+wy6ZxIxL
yU2MpfRhvPokah6mH9BxlHeXx/xg7yw1Jh2FGZYZ58zovHc3PSqpFv+FxhsXC7Rk3iUX4vkRtU8D
s+9vBD/tuS9TsDN+teDmA0/4Px3J5YDa5Jy0EvxzcvST6Y3mKNTrd7PXXBZr2MsvUFiMvyf0Dkef
NsO8gALmrIKGztPVViMziBDArcamNtfynkkZsN7MoyzvXi0Mrsuq19PlQ1lyrmlwVaNlIxNAr+3K
hlAsgNSwVDJvq0x9XMBE/B1vQGMso5LuqZAy469kmVNm+TEu5M8B/bukTlk/mMHCpTQJs2GUpeqN
NYaM3YQ+0hcPKEcr2rIQKv0Fhvn51Nr9PaR3JerUHIOcOq7VBfyle5a0haH6Qb1Uf87gHc6ddigx
TpxXIVLr1mK7ZE6HJXu4FRb4rjEbZNladlLaFe+sNeAtz7RYEuRpycCgCGfGvU26TLalzvOPmNyO
fr09EYgGwCY4Jd7nAn0KMWGe/Y45inMVZB8RsfMvgAstsWQsX6c4DLdBEmnNozlzUZEoH2AKOj+I
CJQw4CQRkQ7/w0nEtRwNkvn6GxQ3tHM/HUhtzt31IX7x2/PLMPDeaXRtbsnCsSNnAmgai55ojaFH
kxuhkTIeuGyKDLtMrr4ovtFaaSRssJ69JUNM9JLBoCa2rSAJ2tLhQj+fJGonPGVcWjDbhd+cdds+
ggp8KaCIAH+CZsUgQaJiAjGYM214w0QkUkWN+fFKsNrwp3bjAIAvV/xvBeAg+7e0Fn2AGU9gEd0l
6kcf2MgI3/XDYnNmBO0Ida70U0VIie964Hiuoyx7TMybbN8vig9o+4jmOkYszJXDrWqVufr2UtvW
0dYepGcP6BM1mpBtuGTUi31C9lt42u8RW47bOvQDWm+6H+6WatXZzYLqr67T3FT/t03nuKWBESrh
+QNubGsqRjqlKlXd+yFwXTU5P/14NFLDNk45lk4AGst/wGPVtesXMw9UIbHsYneP7t+OyCPCF1Hc
6lEx+S49TEZn3OnsIlxCUixM6nSGLPFisLWMFZ95718ny+OgAp/7UAMOr/2mjMlLGLCMovVZzqHw
MAvd8zOw/tnwLa27YqZ0TVlPcfwyDOGzMsL9m/OGcziX++hBkCGDLhCJTw/yyv5D81BImwtekeU6
y6VGqeML3M4o3pWetd+2Tlek9J25f9WUoOz7fFalXlSzRV2/KaWuVreL9bT6fH09Bh2vNYW8tP1k
x3eYGxmxSfsHXzFUNAnrgf5ikh3pVG75+pjrOG2dt+Rx19Ip0CWQulPQmk6PNPC1JbaF9pV+IZVx
bjpKalXtG4FMXl54GnFLkmCCVOZ/fTPOkb5ditomvdI3ntsn7n/+ID3pQasPmxepJNkFD8QN6aMf
6OhaLLZKdVHq2LDDAaHuFD8zGufyYiMneyV5DogvKLkOWj0pWxr44Jg8SExsfpp5Af2NObzmCfI7
9jIIe1tCwlr5FDc7WFFAUINoiDmNOUeOsh/75kahZclq/cZ5Rb0ZyJjvxxEZzJIQ+x05t8SyWYPi
QLL6oN4LwNLK+tELMXVvCR+vbUHj7658JQ3HLLdLlkl8oKy5asAs0fU79eGTiyKcpqdFgZHxWRFh
mYxjhwMPcq96j2o0+x9r2Tnx6lz4RNEK+RbGkeZaIeyirk8nasaSnqG5atQ52meVc57rf4bwn/mk
Z7NHRJlfBoMapbON4DZ/NA5u7L6++XLWLlw0gJVTLlFo8twUkyUgep8Qefjx3+SBNKS8m3ezrea6
qDOPexziWovRhClOXU5AXbbcOlSyobL5UptT1lcIWfmfZYT8pLjhoezoOqjICd+6dwD8s2KaJ8XR
/cGHrJSKTMrsh88g/daWqRNHvKez02ahUcNsz6U8PnBKPyIlc8e78jk2peI3xAmSMBmZUe9/Xu0k
tj3AeeuUFwkOskfJz6wmhRMDnRxBbWlVPjfwTVzeW0t/HQ3Rg02SVTO7CmOOcxdxs4TWk5WN9ltn
aW8Ot9y83TCqiIexRVoGLmXE9vVZqQ0RnE4MTF7YfeLJb0z13SaHKVQk2p91HVOCvGHWRsBfGqv4
uidBJjQFy+xEZjPMketTCo0Lo2WEviYER7y4jZlZZwg8+ouxey6mYcO9zZXTsFFxPBGXHsY4xNLV
5SdT9+wdqMSXUGMzP4CZna5tTr1105LZuAr/9vKg73FgTMkcknlrLa2OZA5ppbm2DOQJtFlPJ86+
5rnIW6qPqGo2kT2WaGVDhNpoagem8aEf1MGeHOvUYv8il5rNTTOZmsPPFDlWutlLdm8u5BPrrnJZ
l7k259CA2Iaevd7DR9jbVtSaNQVXUQCK9BuKTciV2b/d/8vfZEOASDcw3oJ0rp/sv0n3KkoXDgMe
+oOO8gb5+Mf4H+HQJotD3LT/X8RHu29f/DNeta3iNqqR1TFO9WfRRyTlBCR0xYpZVJjJwI1xMzPF
RwXocFI8yX//DSHHVk5iqUtragQ6CEYKZAQWW5wHZ4e/Flm233iWPJsAWxdLoIxZ8Sw5kP+5XX5H
nwVkiNPsJhCkY/LkTlZGpQd0JzX4vNYXzeNTPxuk1aSnFuDt58vt55Doi472HrKxktYfXbfuUqEJ
7d7Ei7JcvqYC/EaqflGvHQVuJqAJUEtrXTasEhIG0ryOfWpMqoWNiqHw4gXpqOR5WHL5uvXjjg9W
Fr/lCG3e95yrAgeK+n8S+7EHYc0opwO62Od99hGcoaMHgQXCbdSHqxFixUSnovjqJ05dfe49crMn
CjcxmAIzakFPkfQwRYoLblYG1IW7OqOJZL8LWvPRaC2D/MIRwOPQLEE9yPDhrTgTJN/oTYt+M/da
UiUOqEbnoMFNPePEoIw0cHsGahvJc4nPIgsxa/kTma28L5zSTmSWONm2uN+CTRhfB3/Jia34gyYW
Rdz3uPnxvFy9vxut9wAh0nPooZakLOsnxKfn0PsXovJxr3ElNy8hgn+7mG0nL2vuommQvtoJrDvW
kkUK4qCeUfevq8DeaDHS/d/CtxiIL1pGR075z5hX0F5z4UZHnypIfoMFIy9KeZDSlrnTKjE3mede
/lRy8OwRY+CQxXD5Jybr/9yfP2vl3i8NHncUQXPXBcFb2q6qB6aY3r+qmpct59WZ0r3w+d+D82LR
JgJ5plR5puEag6qHh+Mx9N87U6VeDS5i7PXcTjApgRG3VI5FAZkNin5GkSrfVBnX0MeT/0ESsaW4
p2v9os7X2SNRcIPUYS3uljsAquQHNQvuZG3Cn7Ik4uEdja/hl5SwiMS6Igzk5Hk0bs4yQBb/wguA
SpvCCoEZ5aHdkAjqUD8oEf2NMNeaYL63tTR8XDu9rzPSuf9n+/Aa4EjZTOJ42m3Pu589j4goKuAk
VY/u0EEEBPSup6EgEyXJNXJEdZdmtJzv5ZDr/MdpZZP7HkIn+FGz10a07b4NOhzgaqMIGUnsvxZn
k/YkTDBaCpSLE4W9gTsABSEcV4SMrUaPY1QdZ6+pyw+8n6bq+6Mvg8i2CgGSP0GwuRMsSVuIFsuy
q18JfMeq96GbiHAAfCE3wCI8BbiZOnM1iCUkg/u6Us6UM0eat+2/+xhT/aLvTCr6qGAaJuWqxxdJ
VJ7vWA8/ZYPj5nbAMwgtUVeQmK/iBMesZbzahkGALEw282F0JDXGZwdqtFoh4W+XCgWJcJiznfe5
7u02whkR82/ONVlafsdYhLJ68T36ivJ+3rFYtuIcyxrQbX2tL1N6EHl1XjuRHHlXZsyW5jMaLOnK
bcRbRM3lSu68PvsytyI5k/4xkaw2SNqDVQkYWEms80mEYJvhGQNLNOWsqA/drQn+UtnpElECt32q
mAYLJTEgKH0Ajq5Z4XhmhtzLNNhA581sdfr7nAxH0NEhGbiA6q/nY9yPQszE3dxtqM1TviuOWXFb
ZzQ9pWvD77HF4ruH1rmC176UgpW9HOFLzlTzy2l4bHcDo0pn+mITdTFRvz4itcKNVEJJuU1xYPFm
+Tsd0UghsASg4GF5xiInjRtreeK+g98n7NvM0BA4f+6xjMoQABw+LMcNB6uSGxZP6YuXYQb4mLMk
EItEGbVxVGb6o2jTAQvJ7+hGLyp3UHanwkYwwcfkq8zGbRJ/qksYKaSHfP1v+vWRTYsfeh/v03BY
PGnTlYnrZDM+iTQnyCBMAM/Sg+EpuknzD1+4kaLuJHwfzDOEeBNHmoSJ8sCT1hkuneilxLk3I71S
pQ51QESlX8r83OKB1pnQl5qYXgo4V1zDhoqr5ErFRSZhHcP3prsD9Jx4et/1WcVGb1B/wcnYTY1I
9gruHsGycZ65V7rNTeZJm87yzhaVE0Q1/kzsWbYBu40blLP8b0IiZQKGi75j/dm9iCnLPIKO6F7l
4MA1dStbtDfR4YriwR2l8LkQAE3Ui/xspVct40PFuesu+dAciFEZ5s+mbIK05/fqmjSA0C5idiyf
xHY75oCYok3HA2kNKTfIOTCs69GY+1+k9rKmG78YOMDPCOoGfOU6Stuu//kvCphggH5dKmCAPyKv
k87ucIlAtJoj1cMAJnllSwkz04QUQoJXXs5F5oSUWbKKtC6YgAG4tSVCYYmEgThIKx6Ojh/pQN/x
2zSyCPvPzgGuAcnDbQ4HFwC0BeKMtiZ4DqJTcaT+we2Y7kli3XnUPDbXAbvvUhq0RGHl348Y5ia6
I2qN+WGie7E3Sqq2457cKiF4+mEt7KiERhBbraiobcWHXq4RMYlpq4r6LCHc02ErVKe3WVO4rE5u
STl06G0qsLA219/xPQ+7KNzJtYB1iM+KVBdB1lfMc0V63fV2dfjPdxUhyMEt0/KgkoSAETLJBwky
TtB+Svy4cUnjkcZrhickNsKXD5XxBCH9ax+difuaX/WQbu2bj3sawTiHNtSMfoEqt2I23LCixRCk
+1VqBvwt1owS99iwmq1VtFTshE+TqYZh3brIjAvtH/gtzPsTnrqx8AbXOU+ISoN2HC51QpXCnhbG
WAipuZqeIuzjH6q72F5fjvWYTBOZWG2MBhr7y3AkHtM3aWDB+NFK0mh7RZ28PJ1QPNmUdhFVfn05
GgnydkULEzwnhRY6OAiGXNoO1YCfmlsaWamNY8xd77II5zacKEZT2UFB+8MI22juMXv559qLMovG
08QhIstXJUV6solWbb8BNqhgAm+uNNAkiUi40ATz7VmlOh90/DDvqCYNAVTbGTZEdFwUhFYZOwLO
wtE/M78tvF0KTTqnDIAjCzc+bpAy/I2LRKVohwQ52mNArNhGa/GwC8F+Hw5GMhhOB0iCVa776f2R
GpsFv5IFC9YUTV6g06xHq1jPaTvvUG9IfSLgwi+RutWnC7Dd8tXQH5FXpcQTTd7c/EPoTZMbzUKS
G81ueRfQ4ocu0QSIuB8WNJ8S0UpUARhZueFiPojX+rSyqI2ZoQKal/QbhjfMDLP/0paIkj6CYHaw
9OSeeuuWp8VKmH88i9fBj2V0oJZhizFlUmjFbUnY+XqLa7l2moLz7+NLQRJJKL6IUifhU1orvfMN
A9Q9i8s6QorNdXlgr15yjFlZ/2crJ9S3QQ7LntvuQPWusB6FWcIe8oDSkYFDjIciKHp+BA5vBz7m
xQedS3Ati+elsDstUaOTCQJzJuUppdtTmQcykDI305VI7QYxgjrHe9JjqdCwqaBKoh8UQ0haHHPg
sJow8KCluFw18uYLIND8jnqeX5E/6fG+t2jGjHNnFXBHS1DshQHgqXfLg5+MllPeBlN+FhyXNlOh
Imq4IJ5hYCYf8Iy0Pye+ix4dkUVPVm7hJMogvwbic8kwDF1Tfs4xUKtodDlPDYwPXyYSLcjGdWZR
VwoTcX+hkNDHQF+rBluFBPo6zKEL9YQ0Ec51PtwddKPgLP9v1favxh4cVN2QcNq9yDqHMZJv51ZY
Yjz8hEbqDgBXi+w9vs+TJjYzTjNv4KLbVmf4O8w0e36xvlHtDGiK4Cd7XgLOzZT3DSoNQn8xnWIf
5esaiwRI6N+srbrKoVidQIGMRBqRNNIV9O+c7OnodNxm+rUobBMmHflSNILKj/hT2NyFiZ7JMf9g
nEX/MW0BM3qzCpYb7MMPGiOw90ny6twj0EyOSgtLh+fFI7037U7AI/eOs/JAky4Y1quSV5QbnYyu
zdPaghbS0TpAjE1TcGI1B4fh2E3TncLg0MRc16ImarU9fPH52JDw7clx1hLYXuTBlDqbstYNO+pN
ZSwt0Pqx3cVvYiOZI7aMjf4sxhhZkDucUQfi9E4yMwiwBcm1iTNsdPtaPQFgbmVWMNJnow8Usiel
2YH+X3Edjlhd7P0xrSfWxJMegoixq3Dzke22bmIIsLIEFUmuLQTsMCPPQxWUH4fz0j616OEMq1ZQ
vdLuWUH27wSGIr99I+t1bimWb33UHeN7Pp3hNJltJFYr5YiCCXh9tjCcQKiOPg01mJoT1NAQqyA9
3XRsvmZTpezybD7TP5QB7pUGp4Cf4BxkuEZc0hthv13WtWRUkGO+vJD0GxKzSLtTD6bIjI2BJQT7
nYk7FZqLPRKieZTeA1sbZnfw41Chd7FOMwhJuNMJm1Lkmemcxl/bQsEwljfBSlILR2QtdjsfSakp
0KQoISgNddlCyErEAx3YPbUvezazwzwaybI1UHzB072dACQGlrqku3E3kLYhKvKysYJhaqbQAEBK
XI1MFOOFB2j751GNTQVBJe6YC2cXxQ560qInVyukAekeTNc7bKWZtvcamsh/PVCueoSxXsjrLlFL
cBT+OfQlpsPryI6Jfk4jDKU+BKZmyGGBFLcH3YQC5y/A5uUVccskzh2GI+36OuqfsmfvpRY4EBCA
QyqsaOrsAmLHBjSGg0pX7MRn/T8RRPDf63k4+ZhKq6G4Sl0I0mQitiMcoiXijC4WUc3PlbsnBsq/
Nl0mwC8Fkkh+HJvqHPyu75+X9OGYlvv1+K431Dh8oKixpzlbAONlcDBzjoR/UA3pr1lAu4WPWmBS
N7u4F24Q5lSHEK6nv3KqIN71AyS/YEhJll67ptzS5Y2ui7gST4EeBzX/XQSoz/6EP8np9ATuSb9j
/MzKIUKXh79wN0wp6C0xO8G0hZv4LoDvtUK5aONSHIK9K2QhQ4e+uAUDO6XfXJAPisrmeuxZWRgF
Qym8kRjYqxS2a0axqHOfQKasENnZJXfL2FsabijYQwATSjGISE5uemdYZVB4YC+gYz0+yWxjx0ua
+GrE+VTn24hk+zqG6hqahd5c1YxNWkiCEK+jBRsSDLNEGmNIBshcPZ4jbwp9QMLym9cWo186gQ0a
PWjTaDyrefuSDu8gNmkqF2GLFg8qQBD1XtfQ7cDGH2d8R8WDK4fzFa5G+4vj5np+iaDQJJUmt786
SqF6VzR/ehgZ2JpoTmqjMySipcNABSkoeXYw+YEdNnKSmNKeacFYVFS0iEfKnMRPo+E/eKVoJ8UM
Ubj8G7Ba7JdKcuUsVyT7W3amTjdLsDjyhXzN10189RVEldrGI3KB8BAtpvBHJSWmerTKPOCMmsPU
wjrcRZQW5vsuSuBwalMcF/b4UnM5Ig9J77cCHSwmFZ5uLMHhuWNs9cYOwOgSvx8HqwrQMc77ZfIq
wB2124CsylUeXduaK3wLqVdKPKWI7CD951PXVhgDYDiIHTr0G5VQ/qRpDQnz3vFqjto6HHtfewh7
1UG5fMFs/qqQLAYsnwqyJakuqtG0xmbZ6JlWBdNYGgCOxXiJOqRWaducDtE0XNUwKNCmw9x25pO/
0+23pkRCWMAOmm7raI7mKbh2GR1acUUAb+DiyoE7oCmnZP1Gdm+u05X6tRIGIfGouQRSsm74A+Ec
DCIlnWeyryxhWsOp/gUyASgGebi3y7jIR1nrIuMFbSenh9kOwHBYfVrS+CZKL1uOi9obstGogvou
Mt4Pj9WdGZo0D1OFhGE1pEY+Tv+wGhSNGoljWj0e22gJQD5Y/atYiZYy7l0pI08EiWK7qYi6nhsA
+dPc3h2UsgnLUo1PrJXg3YNU2SNGwpo3WUrWnmr3cLojiGAMVczn/EryxKIqrCHUQgrE0U+a6V3s
xKUfaKkuYwJVPezcP3TMyOWsusoJ2nHU7ntWVBxyYow5O4Tss1ytZvtaqeqzVDZ/SHC+iWpPHQJg
mPyXotTqsIJH47mJUajUQCO7UwCE/YLh2w3MoFkiufsAoNY2Prrj1V0Wo4577LO2Z6SDP4DRvrGD
jR1haJwxfmdOvP0VCzhkaej+dzKoEPtr6eVpBE5mgq5BJApSTT6UBWyncZ8A3NYMr3eEcTtIB9zy
S0AWVtPDP4dLaTc8eSA0uN4/yDw3Yoe7gyr1WvRw3QaeP5MvA9OL1TkR1NjmfxBLbU0ngmO5vG/r
GM++PqWKy0iNItLJUJM+n8bfK8O2Vh4sAEtFR7b1GsJ9NQEV7hE20hdMEIRwovUL5bqDbA2L4zyF
5Q9PNvQqbvrP5CJ9/xROI1LSXWg8uBZtsnpCEu5AY6jKzS3rLdKHAsCwNhqkrS/OcqHjmqedVh5r
T576GFo4iktLI72nWRsBUmWmbKuAXHipLSpaPsTa9BF/huWu0qnJBB3LxP/A7+PSiBQGzQfSML/g
06Y5Z/nFJBpMW9Q6fX0QWPbkXCnO6aK3AUxXuG/nt8y2GIM2jD1QuaY8LfTfjBvaYVMEZak/BVZc
Yn0CaaUu42g7HD6JPrd1ZumE8vuqEuMmKIMZntL1u72/rnyb5QF72oA9JW15xTtEUCpdgxiXL0Ky
gkBDyOQ8NUfSFgO2EHT3LLWnHov7BPkybzOIMihUf5nvIyOY1mFgrMlkguwYFdqLtF5AWiwMZfjd
E7Aw3cnGhZ1smRWI8NOojYmxWsVpNy73ZQy+WMYJmTNix+joLmWgZARTLHQzzh6rnCrYz6rdSwie
U+GL1bwQhmNkSH11MuBHBkNTok4QncqWrUzr6ibN8pvxPmapENffQcPowkTEkYVXJ0wxjeiof/8+
p1K0lV1siUUZEyJHgL+PxJ9fe4k3xqbaLhpGT2ec6vfD2Gx0NOEZIsFgaAjlp7IR66vL1/cmFgWu
U/Btpet7ecyttW93xtMs9JysE2S98jRKtP5BYn5g5iyIdvaVqkDXEciN42H6kW8xs4s/sf6Sc3VL
j5hJxeeFi6JtMpT4lXDpd01tfPaBCmCNkr4LkayDze/OeSSo5SADY3ZPf9/A2wYpkXEZeTYrC8zA
i7U5wMI14jC9aTQrikrDhEL0R3EdPjg1tbiauuMrRH+xic1aEEfLXEKyl7BZsVk6OzGSDbWxJP9m
5e00GvDMAZdJ3bzjttJp/109KWZYDBe59twg1Y/lFoarmt2raEAFKiEPTg1ibFN1HwgDU8dwpp6C
oCTQ5cGrEjKkFpO+bEGJ8Y6lkofMd3S7PR9NUaGalJqY5H8FW1RtSOb56pfnywMU0/qrXdDzOT5G
s2kqMTqu8z4VB+K2tpsrasr1CdgIpRp+XTYH+pwZvhG3D6Lfb/1GIcymWuxxi37S4zxDjmX7QXgl
6E+xZan2nk5ABtj5OOYaTxasyZiRoCCrqcqEHoHICE3RSDUz6gl0Z7QfShnESfVoZeDRojuMWPjx
VxUe87GiFh8r5y5UnTbmfWmoutchgGxN04evH+7gJyCiMcTd3J8l17fFqFj4tarH1AU5jZHCIwKF
XjoCQ7XO10S6PkD/6sIyyMx0Le8zdsOz9foRnJGE4avGxRnJ/YSbygeDKlH0ibftSKWkiJtUOYEc
+Tzv2klGQ7rI5SYH0Ep9S06BRr9pO83FUb/rpOWMMqNXgdG6e+PvAJNrPwLdJEvpHp+PtTO0D+WB
WwVtKiFU0fD8t4QecW8ZV7BSnu/WmWEcr0hFJrJtW8vnx2cFYKyrhzjZaWYY/hLJS0IkOdgOxnbM
5VdeIT8p6d78EZftsG/7RryJ9WEZJAW3887XyxxijToYd1yt6v+VqvIX4QLRV7Y6qRlKu3ZCEGMw
Nqh9/vLQftJmcIDVztmer2RvID+CRh5VJmXiqKNpb5KAmIJuInWDBeJ4wIlypihoLsKnXkzxkbwS
iJ3e0YzQai0xYSFJEPpPFUbuprm27l/YhwbuI60DaFzpUxMwcIKfkYnyvT+AFjhbCFqBUf15T44m
DsGQri8PgRl6sv95F88YDTUEIyVgZ63jBK2IsuHpeyQH63xPdTw/duF5tdd/QHCRCVkjWBR1L+In
MyxB4yaOPoiO5mt/ucYEjCItcsol9W4g7gqyV4UoodmK8uVC4sxG+KA/yTfGerucZ9LCGxCtS69j
FX0gVElwgAZhr8VgfYvUW8Y49F4/oQq6Zdvdlft6Io5/YLgYpF7DNKnGahJkFN5F/qqS8Ln9TVCl
qT0NeA0wJ0zdVvYDfzx3R5egYFXQo+Q38xfEDt7Yp1CBdzVXCKnO/ACkLVP5ran5PO+w7gTY1a/b
Gtlk5GwppcmVHYf4FuozJ62zfgL3RW/KcB4h+XUdrGBsBBU/HjQaeSJMabItuLlBiHS80SVOILcT
0nl2aSUggEzIqqnpjMtNSPXktLuecXA8ni8wY91LpdUxfz7ikJevxJ96dI+wZ7vJtuOTHeN9WJtM
teP9ix1whuya6PpguIL8O9kAmdZSNT8GkBe/FSUk4zs4aDTNlHViexSSEBmGedDf8JojkMcYianr
t5pJm574boMXTLE1gDDRIX16XoLcTnoT1wVUHdtGAiAl8+f4LXleGG8tWCmiXjlmWzqDzjmVKQE+
DPTcaOXiyNgt6XtMM5xFx94oPvtDXlNUjuGwoKobHnroXxrMRDSfJG8zX64EYgAwJhBNm11ILdFg
qJZlvASwcdCHyHw0ZhoWBLmOQYZ6sEKiT/LGbemwPH90wLsPTpcnLSX31eG8S+sZTNGFqSxMqVTi
v8PF/UlU9Kgy1mRkV9mW/q7tllP2PxOBtCl5InrhxGf1GLwJlCBqKZfDi3x44RF7bC1x1O6nM2iw
bcK723AQtMdEJ1pUPnf6pHIzR9r78bchMtwmcyvobkfny9tkorrYWPQno0a4itUqmGsQFw/1j0jR
3pRwNx2BZNn2nEzV6WvyN2g94dWM6fODTGHEkGsVIGe6qs/fvZ5BYZ03ow8e+CeO8vI3qgoU4D28
fxAbQyJX3g3DWVzjjBn7z4MRcYy5rf8fS0f7Tcgl7rnYUEHtx74UgTPKLeHlrvk4YtURncCpzYSP
QIgFi74rspEKKLEP0mhvM46bq/VCMcVqJ+YYh5h9oFxq1BtdistdpX7kgtMSDoXbAei2CggxNYIa
jMxZESauAWAaJFHEHdjHu4JQA9CxmG4ll42myUZlpHTbYQUqFIOAH8SJI6aAHmbAPlC79zATej5s
Yw4ATV68Db/TJ/iR3C4o+A+3LjglobPgUGEIcgHD5Qm/CXH08k8YiLfOC2sii7eHNSn3PrIAnbNE
5H3skXHwIXk6+ia/egnNTFQ7Zsewd8d1VNB5co5EdZEoP/uRe6a3exUk63trLVjzws9eewTj740M
e2LLQ3lvfOtgxRDJpbp2jAkROFsQ52Ua6oJlh0hSB03A9zEj5lGREjmF4ubSWEyf4SpIi5+FdDWa
hBujFXoYyHJyX1N6MeHknGY1HzuWjlp3CAPKUXOCMorDPL2nlZk5Aj7v1r0EKBhyVQFu0c1BL6N+
mHq3OV4TUr+UZ3WA1LPUBqzohiUHxSMVaFTX+nWh6dUpmFhzr7/ejWgTH7fmt0l+ceM3/dix+Xab
vclP2FKCLGtVLiKi+gAJZVvkndRBJn1YIFddMChPxFhTEQHU6tV9quiX466Kji4zFgArLV0I3+Gh
dsCJ2XpeYrlPJPmsYW1mN4JEFuKhzffYtMe1itddN/xAwFADkG3Uu6tQxaO1/x9dYeiJ3DjUigiB
Xtqtv8xIWNxLO9fwixuWWXDtfXy+WOwxGURiGX9gfQV67ovpLPo4Ot8rark1R0rUOoOmmjyV2LWo
4rp852DB8lqZAyIXb7YxXkcfcgLiKLquOW3UIHDHHfDffeDS/MWOMBSI1UbnbGs9pw1THGyVzinE
ERZTBw0empkEtPnqJgvK4eLyqZmap4CmS/qggkox2jducCnZC7WOuMWtMj+FduSypZxtqcUmwfUp
if+JY+bsZNZNW4YlhUEdcSYd8sbvYqOV65c3dz6/my44L73csI38073P7QO4JQIjkpxnyljbo6pF
MoXJL6TVLeyPHSyu8GxdpvGF5le51rEsMHrjKj6WMzATXNkxvhDhG629V6wbINOSlitAkAnzFP9E
szZ9ZpP0kINzGjGWEnm4RK6E04A/RTkqBIpU03WF08XHQ9Rn323ZLFFaiOr4QKXTFWB76KzaP5h1
+JYlauT/4Me/oUoevLGVOJcCO/QZzp4Mj41h1Mx7ZgNuDTc9BwtKASDLQmd1g4O9QJpXg1Ek1Ntc
dhjC/wUJI5M03NHjwe4rCA0Vgn/z6REmEyqMruZSAgFwxPXrHA82PQSv20f9I1NSHIFcyuycj/Jl
UMeIKe1OWBPr694mnNFFtQjCs0T+/JT6puDIAh1/jd9j5VuSkotiS8xApI/QwleXHBTMiLZt9gTs
w6MzaU4QGVTk+aM/VKGRRK+NVSogELgQk4IBv6wPzFo5v6cHT8IbaMzF9ikmKIe6HybxhmRnq21V
wskLfIGlqPs68J6NhZ6+VSa4/qmndQ2Yy1GIu1PPcAAR7PYPl9YCIvW9YsWiUlbLlTdqb0tXAIEV
5WpOjE5jM1092MpEFSCS8mHWL42dOHtPVzXaTqz06EVimmI4lD/q+Bb7RRYElAW7WUZ/wThMc9n+
XzMgofhSHP2dRdgHvfZLnIrIkdRfujZC13a0u2LFluf8M8yj6iE8+bggpHm3jq5/wzAd19/FuAam
40ABISOa3iH+mQ9JruRF0bI3vtC/UxitA3cL8tr+CGChFY8ONpKIyFwfq10tPHS1BhwcgiZqo6Lz
cgkNcqh9to/QhacUEslnplIdAx54z8fH5GDhXTqV6X9673i25MM2EniClTljTlUUfiZG48leJdtc
SkJi8+INrlcth37l54vVAUBFBdSfFXlvWsuzYJsZDEBCPzTDa/IEG2B8yYJEOBUjaE2JfBEP5BRZ
Vy9IFMwnQ/mtlmMOUB33gbHqJ5P7EXnER4+eiiXlSj2ZgvxkIKgouqTjFop4z2CxpfhvvoW7o5YV
M2ix4/v1muhjQXx8D08/W/EzmvdIxRqdV03s4a0qv5EgaI8NUcU9NuE4fPaoNGeuoTHgPQf+yd3e
JzLTEgDR6bkJ3M/ga2TdEV2JFuCaTZx4B00HBzvqZQcnWpqhTciILfzKBN29/+EDPoClQV/XCwmD
PjCOPFLt5OT6Qn5+Uzs+7dSJhQEYpWrg6Gj1spS3ghxobVCh+pT9mSlKP5qI6/7g19XueSZA1pui
b4XUBJvdGd1klnKdmZIYD+Puut6ClBa2o3/Z3HDdXl7vDsJuHUIUw8/OwgIjORi+q/Edzn5ZLBiF
AM9bvF+zaTMdnf8mxlDwlR8AAH/CDycBdNuSgY4/K5fbzeht0sTZmRQsuByoBmznz9MpAlZ70/sN
ILPuWOAVMweKEeZPathNtnV4DiXVF60A6OJZYZ6BEemKOmtLuKaiCFImoMMVo2FYpED71KDq1ZaX
wX1U/Esc7f9RIXcyYGpEp4C6mzyIya8e73IhJ09G6LfSIl5rqbPNbWCH7n8KeaYLUhEAXxX7jopz
QMiSS3YBUtJdjuXcnBI5DCNn8KACpIkGc27ltTjXolEutHMr4z71JYRBAZn/bEgTRe7P1qR70PrW
lKROhQm34rEbV6HozmnkYC8skfv7iHBODbpnf4bUpK1jjg/bPw5iqMaH4S5FqvRqLQ8zbqdWxREw
AohB63gueR+E0XYOvtrmgSP54wiIzJoDJFLmqdeUk0bYq/LPJ3Adt7xymrmHNDF7eTJJlL7puotU
dsETvfVITSaXCb3ovZlxmPrMKZQ3EoWilgz3YIF/YHZgMaeoHv9+6epI9+9wISpmJhlbMI14Pa1G
GxfpbWMD8w9TcoMz1cVpYcA9ldNRz3Fw6xzceUm3RtqJiOH3zOhh+cQsu+fynqdzDwPo93JE4l1v
f/GbKNaY3EfsD66rEnz3rDupEGay1dbxwAy82PVyuwxeY4YA+KkpNNGf2R+o/bxVyStHDKHzB78t
2Rzzu9Eqaavhh+53k4OgALfokRYLqKy+xILoYwHgGSxAY2pmiIsRER6XsHtqrSMUh0UwCTRU38xo
brWzsXZ3BKdDeay3pQoH5+0UKuNuzBgDgUQ7pX8BGzzRqPpP/nNYN7CKi7xArInVdmg6B+7C+AQ4
CtTpuPO2c5IHU3TMGW05yfdXp9PTdjqF4cN3G38rfY5vuQ+ErnGFkokzCbalZGAYcf5dJkAhVB7N
Vst41SZcl4650ew9lg6uo9YiTKeu5aSnaqQ5+fn1OM+BVYiB8Gd0KyVc7dfo1wYbU1w27LsywIpM
3GYg12id8jV5XzxB+uIs4qCzTbZ4NWZCl4w8TjKslmUbtsM0Lf/aA0sy6hw0jxlzNhn7BT5Ss419
6OFlNuL18Vx+eotn5IHzfcsCpgghAgzG8uZHXEEbKJFSELO5+hjLRvY2CEP0aZnx/HzmxUSWtLGD
STaImcUMAKRPoEglSZ+7hjzlsdBZQT0/giFarHUaiUfRwiP3xRSIGOmc60B03ACqZp9Nw59CnG48
FO4EigRbiVPWtyaq1/6vNqmuZCZ92kONOd+72yUFYVvH/JaDBluvbprlPhpX/Xid5CCtaKcUwEyR
NkQyKNJ6AiPemKhJE36UXKB8ewTvCKvYrpoj302YchPUXur1F3zPbLNTQcBXHsyH/kO+W418j+Vh
egFOciE5soeX4+qhjOxUCJGZQ1dMrQ3OTO/XGY7Y3wJi+EiTVUOj4KKnVq5IvMLQORh/MwWP/Sma
J5FS0UpDu34DXzjvvwiq7DVISSiNpX98c7iNMtnrpFHWOw67CuqMDKFfqvx8fanR6V0kENL5v8h5
QPja98aN+zEHlK5awA3PUzAxeXEjuTarEiwp0RHhpayceeAbAmFEPhUDb3pnJzz97lxh+wBdVdtb
mGItmxLAO1q8l43ZbUAR4DSfx5RBX+kOiku5GZeyJx2Qfb5KghlHJUyvmvn+eyeMBNMtbqtDBChN
Hgq6uwh4hGCvApHpClR9qZhpExa3knvL1si6JCcL59cN9M2iJYsqi1e1icoqM9bcHNY9jCr10MCE
5G2+u5Rn2wbXdHmgpNNkEUc4qDjUQ4h7eQ4iE9ArhIKWcN8jwJEu2KzivvyQfl2fwVHLqTEd5YB4
QSNH0KmAUdOY3GmDoyuxEDDYpdiQuTjxXsZRjQRBhh9c/9VIKDRLBac2Y7SyMLMneEIbbI278EYH
ufiI/FYQVVdnmxrN1TMeReNO033HT/gdeUeKoX719kVIBcVC/HbzMtInDkXg2GESIDHmigshCnHH
U/Wz+Ot+TithuT8oJ+XdjcrLesHjy4FAWoC5aiIM++0aP5Bs9/d811XkQQG7waGtzvbOal8IqNNF
f8g+isG35YVcOqw+c6cCWEJWXmDITFgU8X+WzCba+06cqnPQ59L4+eapXYOsvwPtMWdPVspYs4Wh
3ehvSgohZRlZ5HwR/ZtLT7nM94hI0z7cSfXH5SnZiUb6C15pHfAB97BMpGI2CS9n/dFdblbyo6ls
AF+RjRP6pOE/z6G1Fth5TYzblU4kJXNbI7QuW657cr704fz8bJzwz1lNsEi7m5uv1FyBJLkypB+r
73yGt4taIAYlZDtkV0ej1SY3sI7d3Ft3lyX+sm63ph8WT5ZMg/ee/IXltYXY+uTf7d3YAyGrZcgi
Q3o0F3a+S6cCibduBRKoPSqw0Jiiw+sUOnbsDYaEEV+YEkJIovMBfVdQ7SRfkqVCU+wqHel04zpx
E+Sv2h5pgUrMgEmjAllus1TijuS+3Yir1GFzV3kkXLTOc9CUHxFi2yK7V2df8EpFIrGbDNjnS66f
C6pJsD1B3LBAt0czP1DuebqibE9CZgboCp8oidtW4lEdiJEQdR2a8nqY0HpkDBxol8NKGxfq+ZB3
NFdxkjfUPnL9LQuHIq+osqZ6WT9CKp1mgKH7XFWo/bI3XPxjXJqudoJHiXkMZxTrLZVc7x2f82fq
OLvsQjTBVfV5h0skxDBIYd6Klo+rZHDyMG0PEdBBBPUXdipnjtPURdYEWydM2Xsg+tkwU3iwWGus
FPDzq/MM7npneCREruFS5iFqxF+L5A8jNCNQOUM0TnMr+IuHA7HNYTTGlRdvZOgGE/d6E4qMljBh
TcRgbQ4mtz2M+BszP2mvZPQHsgmWwvnbnHOXdmSijXceQOzGtiU5UFpwKMOXoLuRa+lAJAFOf5JI
Z796iIZSLwZuTDBitIAeWmhg1w9Ef9PsUoBKNv2nV1xEIm8Tque3JztcRWaAh2be0ZV4ZtwXP5AI
EGkmLrpRunKUrfM+UcEebeL2nErgzCuPbf6TF/R1vM8jii//EW2P664PG7h9B/Ukipod7fVTD5bq
eKDor8jhdG4aM+h59/HWmZ6V81Z64zTeQoOz3j1XhT57ERZEdsFDALHS3S+hnw4qCbQHNZsIb/9g
uDVwBo5z1QbLP6vrxpw7GbK2CsHmE5QW8tu3QoiiWMka021+VEu9IM/0EilnEUOY1DfriZUCWMDi
i7SKfe8Mm4MB4XS8r37ts2YxdIkC+gmXHbguAshMe9hfI9jEXqkrJFWiBuwXOAVe4sSHMJTBtlbf
XK9QnQymTGCmtBM5HzlWCQ9HbgooNTGuujbUlTq+JGL/xp4MiILXypHShFxhOMRPjPNWqNLdhkMZ
3aYP82toDS37b9l1Nbl4Sp5fnSwcSclUGSyIbuF/pGeWGa/KSyUbyJT3kcCmA5jCmgcz/p7t5vE7
WnyB3BxE33W8HX/GetsFzcF1Ug54IwNvQHXuqiP1z/fbs1NRiyU+Hb4mDq3ldXzovILjZHklDevq
scS0YZ+7RsJjmnOxI0ycFiU1KQI5tozSfy+pLg7KeLl5FYZpj0DDAeO7xPFZPgTzWTGN7ot8Orqr
kja4KYNnSiRCNoUsX8X/dzH/dGTIRVliS+wCdiGVke/GtX1ov2zC5UVnXg126L9XkaEAyCb72Yq+
Sz/XWnbkNlBXg4x7xmo8yEzeCzG5nwfEdpwRpTcz2yzmTP8nkMiIZoxp1k6FMq2GD20dnl8ZTxJ7
hnw2/C1VA7W6kwhmPw7RkNWxKPOd5t5emrpAgdCzrUM/0DSbnViCsChrwzmfgvEhqyNDmBUW5Fv7
moFbYrQp5HABmKxNpOThGEpYa/rAUouFPngYlw89hlbE2MTu3XpQDBfMd3aFDWZCtukNO9m155aE
VYNyo3koGWvw+nzNZh3tpG5EfGv9CF5Aa/Pm3yQDzHU9ob7uGnf3tvTntoeKrj2uFpu4jEoat79F
1d1PQy6TvhoKtLtbexhTkAG1BGlawKXLhZW8i6X2vBQy8OHxHcXmW22Djum1/Ns/cKyV3fdI5SMu
rw4Axoeosdk7fY9p4cFskEyHDDZi2iyDpSw4Pd1aZqcWjDgE3HIf+4fKDN/coDUBzsFZU5bXx5g8
uUuU5FllvghhMdPahmbQ2aLlfiOwwrJUnnlRrzxMeywzoG8jK/FK2zK53UcqSrVgNPT4zS0uPNO5
PQzci6H9hc4TPlLNiXJXiZIXxaVUWGmYFLwiwfnOoky5TaspM4qNBwDQH9eF91lkkfidccZh6wKY
89FZhe0XOVMU5buOw3NfNFcOag4KmlVWlClAsU/wCbBASeed6ZaxmiJUEMr/qLN8LSKLULJo47XE
6n7T+d7ilQuI2jVoGPKvdSQb/hqlX8l6FjvtZyG1909XICDTmcyItmWk8jpk5hJSzKDzFX/JG4pW
LIj3cZLphJx5ICulmxc4ooyq8xJDy7LxrOG0Jr227+ukgV+VByG9aRz0qXtTwlFI9YtVBYRIYgAB
33shisA3SchLz3laKv862J6Jaf628uhZagXVozNg81GJ+5vnCOfBrI9JIajwB4fe/zeq2v1axF2J
WPchvLiSbiR9LFrx9OXrUZ1KvRSW7qd5NFmGgEZ1rWcVcRYF7g0TqtLzdoxSkmsTjLpw5zu8b5XB
EJLwJ8tcKumSM1OBuMpzirAAOIHHmyB00n6Gv29tzV7xL2fU1tkRkuu/ixxfqtInFKU/bTxuuA+2
WLZcvOOZKicGWaZvBSvCW0QYbkFQ/JJfYK0PX+YGbs41fpO9IZH43caAm6J4n9j6kfuxDB84nHcV
09KqtzLAVJOtisXI0biiReInxjxuTLA+hedhTJGqQtxVtoCCpWTtgGx/2rdr9nKo16+lFRvplDIA
/oieJkipHtPIkZlLki6lL3fG2CxV8wir6XW608v+qe0KalBRSscz/Tv0OUR+nPf4dfKEUNK07Z4i
SWg4a4iLXh90XbRhcA4YJT7gVgmsR8pLjFd97bIAuOXzcCiAu/u1Fq8hHLB5Abta9xPArzqZ3lrV
870WhXAk5tgNZ76W0QfcGeLhMXbMpjN3GnDnx8Z7J9kK1TWhhGQetC69eo2KyKZ4hzprCa+QM3fr
2PWnFiFtOsjWUO3HPOUUueG6vm0dVo2hwsgrj0C08QIC5cvTyDngQZQwKrDp05nO1gBxPfQYXZPe
0AkO881xtJaePvEpnZwO+etH67o63EdhpLwW0sEcRYNwDQfKuRkX7HK2arYTT/SjlL7NENtOI4yZ
AtGN0rxumFHcXCYcmsKPD0wsOGquQkRYpUGCbJfrCu5ELFVcWjXPSm4z+hdCk3NvBmZHxuPGb3Xm
R3SSBYWNRVx0kH9HPQkUwal8iVZ+NugvZfqgb+SsDpcOa4AdAVM3TzEebSY5+rUtW+l5Rd5wFALG
PqxXhbQOynZMnp/W/kdH8ohvQoJ2MJBiuICnPrWvIWwLE33F2Us1WfM/nE5zU8qo0YVNMXjTnTBO
qGcjIo2Iy/khW5Z3psfU1NReuDN8W+ie2pi95rjOxSuqrv+URinfzPL494rUGcWf6tZ+Hbh9WxAX
8ulEcqmmEaDEsOiuUIe4zSFeqcbDO+jhpAppDV8fCBRLeeGga4BJ/QJ7DSSVZO7k7iXixOzkVofP
RIC9wjzjbE4jwMQ3REbDRu2NES5t7qpqysrsRkBmSzs5+IObFUEonob43beJ6sxfaOeLS0M3KUJO
XW2i1gycmaREtxQOlPXBvSt2R6I9qOP7K8YJFtDx2OhJMnjSjAFR90sGnYKcE8jEanf9EzzCgF3x
WARRvkSaZ8KPrnNBni8VnGWm8C0eltvHDahYHiSnt6pCNAZUflvFqgeit86/miMCakZFPfl7IjEd
sC4Zbuz5buB9GmchqGsxfSmrkkl4lKSyeclWFZUAPgnIa1NF+57s9JPzoxnj0FyqoNVzch6desHD
ztyVvne/zbafwdQw49sCH6Xrsh2bhHf5gJxems+51xxG2zm2tNC2A/FcrKYI8uzsok1Za1P+c99X
FXYQXXXO/2cK0Kg5HSS4NbAJ/1mn856BMJMcWHy7AkdHpTQt3RWrIsezVA4EVdL5XReIpnhV6mUy
4iW2ceBV4xntzB3+VhDKqi0FzQh3JAc8RtWfFV9L5kP+9rnpzSZ169sbjF5U0+mC94nax/RrI86y
JvoYi9b7pArE2A+H9brue+G6tlhephAUZLZdnyf0Zk9WFMfABMBkVcIEG+mR95EpzvI5S4M285GZ
YuDPRSi0i1e66cclPTQs4Ck5ZJjQ4EKhXdCb7dzNyZOl4WTD6qqj7dXZa89xwRbeHwBUkGuDWHDf
BYsJldP8OJhM0rfbZY7YbcENaE+XFrsK7GF2lA2xvLeCcIqASJ0CDV5UhYcvqpuU4XSxJZGgKJ5U
KIgA4z+yf/dvM4PtvWC1KGK2QvCpqLwQXnrdEtm0Gc3Clha+Xc/Bm4dk6buFyQOCOr4vktVKnseX
sRcnHWWxhyeJaGbJ2dPsmhwPegNFWdkuFBYtxmcqOsPPAHe43gCa06oPmxHIdCJaK+ORQ/FY9/gz
6SJZP66DXrirwrWXcXdlXgmYCMs8pq9CTD1eE7D7HueFVJ3pUqhRAbXaa+v0VAhfunCkaQixy/u4
SsZTNSrVRl3w7GmbwA/TKevXgfn5AbpINwzqZL0kAUBUm9b/v59Lr3Srr/BIWsSjW0jLJauScFJ+
M9tCrRPCqnBstSmesZxr4E9NzhlBUNMDlR99k5sLNGcXrwnDqZsSU6CVBzNwMJldFupbo7FKkN3r
fNaEfAe79ifoyNuH56gVRQIdjfsMpANTNCE0SAAiJUzQf71jSl2IGg+9Gr7bamoCHNXSdK1a5X/T
pFR4nvTJ7ruStBZcFIqfTks7+wAunw6y2kXcwMQchTBSEJCtjzLerr/7aiBEe0/2U918oAFhdT2b
g487k3VSKDDTJYxYMvR/gHIoTsADtkJORHj+mkMe11DTy95H0K95cKy51e01JDhs2dGaTPwLqidZ
r4Ff+c0zvKLM3yimBfHIXsf5AXlZsGxFR+2lsJrabLWHFqQ49Bpv+Dpns1CwXfXi5IAkxX+iiGs4
ZuyY8oO0hF2hiySdOelgdo/4v6QTDaR7NeGvY1/VN3Rqa5J/tqEBO5JiKJ0Qbt0wTmcSj3iBTMUy
lv7N2YHsYy5P/l0yKw3cQFChQbARl39DnXFuvfr2HrW2AF+ZCQDV7817aAzERBjX0aWJwqp/MuhL
toGx7x2mOoCEaY1oeja4A8j8CHDFdnn4sjermE+CcDmV5Tsx1xsPlKbEut9GkOUJgCsDpnuSuzX+
xoT2tiiQ+8SldPauolp2Ivbopxa3y9KbatwT5VVJeRZBbJpjrOCslLz/3hygtJZ0llUS/MFzOnKD
utaYdxNlly5xFQkc2rAZk8Z/ViP7TmYvhR0ObnFVIDbDAg9fKDt9DRuY3KC5ibBnMC5l3Go7BcSz
ETTq92o1DrBCjA+I+4YQOP//n0TgZosscngJu0a3xH3Fs5qOPAdHXnJjdP7X5ToVBZXxPToPYMl2
1rCsFZba1qt918tbPjJI3WezjaJmXLHzzk8rtgRwN33DOlVgIon9pF5Lo+GXheV4C0gh+4cckRjR
STo2fn3D++CiVuC3LgZoxpeUAs1TVXwKgu5XN5szgwZuKBHvvizEpgcc6LcBlhlFiTbPe9iiCD/T
vIOv7+Hoe8b0nnSKdpSxuzH/ZAfw6FF/e8KOEemQw/LljbC/bRnV9B1rCkKkZ5uYUXZKDdmMDONP
5qkDqORINjUkH225eX5DIUsoKFJUceB0tH7Bg/OgiVJj2t4zagY5sDIu7lfpBrs2estkDE1IBhFw
hftJ1FeMoRm5kcLKptnVzrH6uffZhuDrdfRiEQOVusOcq5cYfb4s5cekljHFwIAqvJM1p1dG1U9l
rB+DJBNEl4dP47Z6CJPS9K3Ga0XIaeXMX2KLnR9tWCyW6A2JznJzTgkb2E+FVVcfkqCr0Yq8FPpS
+A9QdEerv1lbqOU1/xpA8ew/jSdeaEy+05nM3moWjDvcLXjIL22A1J+KGILdSJwU/pq/1HoznY59
SRGZCzYkbQUAKKaLCCdAlgSrbO0aj1djym6g0rEYWD1p6YQHbn3Mb63Yq3j3LEVD1NpGMlC86Oep
9iSA4inurRQJuQDiKXIDvCI+M6MBzlgK4WhABEo/LWXjIooiEAnuUKEv0BXb2WnLAAUKaTD40xqJ
cfdQKSLYrq1fXalspR2/r9siVQe3Avh6vELpywxsl75XYTZp+mroka8VcJw3iFbONsN+rKPV8pE1
juOvuoV64cF0ccOIXYm3G+H8695K6p8TbCZkJqP35aqYe1ddiC5KjLO+iYDzA/i0tOMU4WEDYbv6
/J9zvRMkCjIE5ualODN7fZpglJNafoNwSlMVSm4KdAbnbkyCSFJ8TMZaN7UGvn10ZzroUkxTfQE7
Rywr29lAky+dQYXC3jBSZL2qcVnOEPnKwyuqDWUsFBMbPNUUjWVyCBrKokOTrP7Qb9hst/hqQaYm
AtuvTDo5O2Fgd4bI7xyUgsMn2Ab7ZeXbFIM05R/pD2a+q+AY+7qU12m2qO3UoeSZ47h1+a5U++o9
BEIclU2Y57RqOHv2xD+KmQlc31P9Ori42lV0AwL9tkI93VQ/Q21boNSKvb6oOwgAk6xctTZN9Caf
nhKu/IM1pSZr1FeOMRz0PAsTWtJeOYyUrJtE8Nc9rHHgt4/m7BbimErdAjFQDEiT1dQNV5xutbNx
wuDhCbxsl+RMmnqXpFA3sg5pq90o7SDr3YMPIxXnrRaKrn8z8oXFHNQBg3CoVlOogDZoC+bULuoE
9VgYVXIfWEgMRADmm0+GbIXBaWgQInCQUfIcd0bt52UDSA0u43wFhHmz5hJugOb34DxNc54DJ4qJ
afssNSTyy8MOSCTmGZ/k84odJTck5uYkd1EqcMPxxKH/XdLG19M82I3VlJQ1RpuwgwSU67R0zQsD
FDnwPzHBpi71J6TGQ7mr3tWDlQMTcYwu5IrSlaGUwI3QPj2Epd05UgxFTHX0gVcCcrEET0k1ESrH
+YpvTwzzbAl7GKpHHbX/2KZQdFVQC+XbJSRtjj/DjIDaeYxMOuJ8dtrJEQ4PsXsRsl+6Ygc3G9iS
WKD+HHFytKEFFn7XiQGTpIKFJzj4LIZaphm81LBTlsuCBEJpuzb4baxwLrPsZ2ORTlQ6XxMzij1z
+CO+w+P8jZaGyysTrD6y3ePk7QO8u3x4NkqFsRWAcdyjCYhTzPVQ3pTapfMOxyGtmdqryfyesWGw
fnYy4TqDGmdOF5s8aYW6Wt271U4Ah8EcN5veiEt689Tennnr+9ve2xSBdRWL1b59D/b6OFExj38u
SJHGUH8vSNYRlWn37ZlqpaIeLo1xjKAQhstK3IaYM2mBXQsqbXOmhJPNUFHkhyJ/QQ3Kk35Qvwtf
2DChvAnyZDQ/JU86A+vxuqcFVmCj9gGG1F8+zyW/CJdsMYexV9ktZlRaUMdYQ0qSaLIdzMbhSIex
rpyP6aUXtGbVuwBrpmM6tpm0kYaApd6gTidalAWAeYyBOHOqpAbDQDOKc50HyYQnTbjLkKVxLOY3
L3RN5KxBsCFVmJpW0o7p3CmXF4RqWQoKCra316nFujmGdjP/uQCwZ29uAUJfRPr9hnsNWF9XgwQh
vvedBBFEYiVyz1PvS8RNLB/ScvieAdEF9Ue0+DjgSCQpD9kjGQlhtpjhbUufHtwC7pwDEJByEorb
PhlOpL+4Eq0UTQbHgE28pjBKQgc8zXBpNRK0jMbeRzN7mfixmZna0bjZsVs4hzJYpkD4x77hhwWJ
hO/qVeY9/kGZcerW6P9Ri8bqvQNoK+kxTlY5h1/Cf0YOu5bJO1rkwRS95lR3+iAsPnS/sYz46xn+
NSpI1xFjttjaIxDGnfLQ2qLhRh0WbP/PLG3rY0MvqjrNTpjU5nyagV8aHzvsedrdJ1ue68B5w8Ts
asUc0d6QV8/f4/UMgPuvJMVqlou2QzxZdhyxtUbiExaggVQJ0Iug0cTSfST9g3kZ6smArYmpI571
s/Hm8Vxm3sprkV1QN3ICCMUDTQhNR7JCCd6+gQwHBTKCUc+VAm/s7fRgI8wFK2G6Kr/Wpih41sSS
zsIHoQQjI2kVXm6Dy4/THuVjbH2U+YwyPgZ0e3M1lQ5ZGeP4hiS5JrDpNIa5PknipumxTmNiMKMG
UhjrfbBCUFiscwcjkLrmZtXXsUSq7yovrXBgSHmp1/24SfLZpwzotw35crQ7gqRnBIxVDSUda8cS
gqf5CaUHYp3p9eS1B70SLuR+bWinTwGbu01Wa850hl2G8MmkvDpdr6YCF1k6cnini9nX/JtWGBtl
kshqRrsTI3seAeLkP5ecP45UKKJdLC21gMo12bzsB4OmU7OgZ1yynYU8gMt0Zxw/K7eTNugVFOGV
wTYe0nHVviroxezA5HjXDwC1sln6m01RtEVWEmBJq84H70rAKXKnCWXvId874bxw4NEtFlG0UgfP
EKOUsrixJI/AVcbnUVluLG3cJk+7YlZ0xmUxShUUprchDmmdxdjd53m1VJFxKn0uXdWehglsJzoy
HMM+GYBGbu/Hrl+yfUP69hlwpZsCGjt8Nwq3DoUVn8i/TyNFQpvwP3MVAj6GCLR98GMW+QMrCAOQ
9g3AYfk/TUtyVAjgGlJDHQkTMrC1hGNbCPh3g/M0KVlLiv4yIejvpMcVi58EadgrU7LnSt6SkXhN
d295OuUdRyXIXh6oWr+8psk1d2o9cA3zGyFKcKJGaBDpmZAU7pKaW7M+L2xFT1VAcjWGk0cJLWQW
52Bp9lF/f9QSxesQDonf2ZQlak6Y4Cp50rNYauuVDzb3947PjPycLByzP3RrTH+iCodvPrdQlYKA
3IBHrlEooFHTZd7fSHUPGHexcCYxmr/nOXGAHOKDu4XXRxBg1NDnubK8G9XUSEgAxL1YNFSTixms
8uJkLk6K3Qy7dbHaqeIGiplWA5/uJTyzaqRMSR0UZlDTHCr9lV3gYsj5W6C7su/rIb665zQvZOEb
MR9M8hoVvpMHkBWJfpWzWmfgTGumJ6Ji/kCfKylGGLGxQY82jtvEjGNi+qaplsxXOsacHi/zoLcI
flGGTVr1cdfGEMFi+bc/rjrQuJEdBU+nm964XkERPv+J9/w22hki/ddFVzxz344vEdkSfBfxepqf
bKW8ri2bO1d6ffTwxONqKYjmzUDhHKF7wOZ2j3QTRheKb3uFU/f98jSjaqqUXWumMEjqGjFdWWGH
NYGfDGBMT1ZGV+HzcAUh1m0ENK1qhJzuxHK1ov6UwWINEZAosf9En8UM2CzT8lI5+1702hL67ubY
K14AAP5hRLgOZPDbFEd8QG6lnN8Oagc21sOv1YimWuPdiUw8Z83zFBw4MiywLwUbECI3fkk2T5oS
upaTVOR6+14RqjBv2KwXKlxlvep1UIOPKAA7DR5qxraKn623a3L3OODKpAHq3HAF963XGlQAbO6t
VRNzm3UWvkhS2BTLSjjXw0wuoogIpJ8//4O117fCrb/Ms3LfXaPkzekd9nUMKoBcbDmRtK6kz3os
kTqMtSKwIbyvCsbrOZ+ThxaJasU28VOABXUGcw+CLm463ywYo1QGgcGxPr54immqaHo/SQUtEMN6
lpqkwP6BHCxErlA5vUjgSzW2Vvnpel2z5Kk/tAkpkJOutG3wwtHQ1LLZaS+/o6J/CBrbRQNWM+B2
sYGDQPcsvxkSYlL2pd3ixH/pPYXVcyaFaT9bVT/Y1fVkjZ2DHRmusT9bZo+s9J2z2T3ch5+hJFwP
G3HvrqfecZjAVyZNE+thIf5rrb6mpJ97a0qbs2CPnM0WFEEQ9dzFDB8tpCUwjVEwvkJ15F6f3kvE
7c+0uDdOBwbsyksFgHR1lNRk9Rsq7bQomtrclWvulih50GIN7jgx19gJCnh6VVMkERV9YFWeGP5h
uNmDpd+ww5KcdWEAt8tF7O6JKUJt/vAyLGrZRQ6n8+b4XAXJ+50rQq3eWUEuEpxOFTpccfYPfCuy
fPKjBU/DUqbVsmTr40geIp1+jBqP4PJar0LyRZ0mQ0E2M06hpuV7clSidmbbFDtQWNH19HHf/Irz
l+G3rpO66f4lzi/3iMYXSiEYimwFSomQwwZzws0qPSH6oUsiok2MnunL0yW8MaX3S0RA2/BV09S5
mJGdPoJHKKES6OPEnMfztlG1VfVxjkg+lGVimNEV4KtTF3dIVEmx+M3q6GCOXY1LeOYtmAiDzdTc
Cfj5H0M17Hr3xyJ3B8oS6kRo/nciL+w0Re7r+bXT08RE5HBIjPhcO0c1FcIHgvJQtHgRFGrC+bJ5
P2gGUkMQyqCJcKiQ8x31I2vg+pt21GO1V+le2Iptg6D9iBdArCqNoo7OircsMlCv9UpBh/W86FFA
JCTV6I4vbwSRAlFumt/NlrS4gz+du/MX+gGBhNBbbsJxkiAqphyT8s0zjrvB8OUHGMFwBuAK01Hd
BTJnE3LXFFNxo75hxqQLEd9bKZla0JqxFW1aCxdXGzMkpjTfhGiZJrl3e5AKcRCncgQufX+mhx44
GXFukKT2p/b1Cgo5upVeiOGCMDFrRhDETYIyHmeDqt5V3EKG2qziAZ05mRBEERpJwTWxwUJik8pQ
lSh2zM4O09qVdT0KdH6JPIrxbg2ZxdWVcixZEiHgkHdUXrGkVDXSHWqYGjW5WwSx53ubPefqk3gS
NpOsoICfUj2/+4GjG0UKxuJstBmzIJygr7jyzg+fO/SnpcW2IJw1gH3egps/bPI16KVXBczdNEtl
Pb9+DO6gBxj3t7ueDZ44q+denXZxcC6sUjhTuYYNZrCWuEjF50GW+x01EF0bFndj64pRjpR6Goi4
9rkiMbRBed+aB+gE1k50s/cTXIbSThqyOSG9oa1uWB6shxh/eR/bfQcIk1Y/+RLB76oAU4I0sMEt
h5OnfD+wbwFiMcPa+9eM008FgnvYVS+g1+ujHAGj1a+i36dpynnixvp2djoPqW7aYBzkbYYpBSHP
kyWWSawaNcxKRzhZfKXKekQhXX/8p/XB/6aapB8gljoMGwIbHpUCI3+Od99uXq5IWI+eKw1eyNMc
NAdfNLvGN+wX2AR9iKY18OSO4mxWcIID4HW6TsbvJWH7qA/UobPItRYofYO8C2iFdooCeRk6SKPA
ieK9+AK2w/o4EjHGcbRffWlmAKJy9iAoX+cr6nYH2mhHJIHemKzQyplabatmvSP2kMwjMlDQrpFn
HZEJcn6VZsNrEbJoNumDsTxMvhCyx/43cGCwpCFoeNxKsde2zoMw1KRLuJFBmRo4OfrSeVuB8lxj
UMzCRUiBek1mqGV67K1vnADMUqyDBjJbnOJjdzleI3HvD6PRpaRZL2pSeUIbdTirxKXxbFkAQCuf
4wfHNXRaBl/YZIQ0CMxA/PQgezzitibUNIyAgwc1Y5t40vlhB0SgXpi2cm0DqJZVj4p/UhNd3UkY
AZ9LrI4SCHEiEvwEGvTOgCADWd00Two1WqSfS+2tqmaqRzBIIGUvmZjbCSKiRvkahRz/XRZH5kE7
FCVs1VMF7PjEEKmVCvjx3L7ULzd0UGESbRRpZObOinfDb0aWNwmjZ9WFyOwWNGA4oEPHYdxJ8ahO
thmxNcwETH2wZ+trUs8+2QlocQvbDZKBS1LFM5x1hcWdvE79BVFIN236G92jOuuKUjdpnJr/qLV0
zhw4IQyuexhTIRyCwiefxzs/dg41jtgg9F9Z19Ud87ABmZpePUrBHZQTK50qkABNPrwARX27lzJY
7PxzTPP0EcX0dnMTTSREMsJsM6qIFWWdt6kfYE/lkNlAy7Ho+oF7pdpJy8XnhfM2tI6oSHc6Ejx3
zX7bq57QRuWdw1/8Onf7nNKkYnQbnkUiIaobUjb5yLyna4saRzeXHSvBT0MObUBkOIrZU20q8mDG
Nh6huLCskm9ekbCy0z5edAbC0M63amhmJlKsQ/Ht8PXser8fCrmVgLUWzINgJJvyVlsYNgspBw3z
CRajJ+s0iLmY8WW5CtQMgzTKyOLqyvZUP3oJBbik3s6gIXV+fqnlog4DLtWQ2ZNrptSRLABylKkC
M0lUkFlAL3kNzSwe8TymrrQqd8gv6eYa+TQqKNgjaowTPLRIfyiSdJQitkFyzRMFg81ZjYDIqp5Q
BmY+b6QepVRirvERJIs3LseLYli5iFQsvvHX+YUSVSG0XnFlmcbwaY12S4PnfhZi9HjYE8d7QDje
dwp5SYA+t+ltb3LO6spZtqtdNjMTCTDDKsUlYdxjrc0FHOT5BEecqLh9N27umBTlxCUZHI+8Kwf2
HKWWh/QRWCussflblLkdQBSxCU89FcK+H0MqPYvXYvu1+dvJrsRPaEvjZBgKHnurk5SoC+xEmg0b
XXpvYFtwnBJ6b7ulwdyW8zLrtTylXKVmvVDCIlNGVpZv694Nm4aEOiJOuoAwLtQ5n7n4CQp8CuXH
imi1NoivWHLb8be8AlpcKD+2WrdJvOj2Oybx0QB5rr1JNHbxT5TA2sXeov/vLPVSypBwejYx4/cA
kSZj3+xvt/2z685s0/MFJ0ypc0PSX/78Ns6LTtTZIVqKqMDG6ZKB0DhJSLmcyvLWtY5WnU4IQZZD
KW8uv7aH18fqcn3YYVHYkwRUG9V+Eir+40KVWpMWVSKlZ0iLbXDpWOmmoBjXLW6LM9uPkPj7tSzJ
ADRY/PZV2w19EWsZsN9db4hkSf1cD9gDIWLEY75qkIc9wzse1HUMUjWi7/z1fvYo/7wpJfVELnuh
ykymqvRAroCabM3Du5eGsRUTUVE3JwZ1Q7ciJbVTD/sPihFL9U6xVOp+U+WL4Alml0sjQlUwNiFt
ntdytkA4tKtYNfMndBE2s8wpSbhL83sLC8jFPtzc766JMkUG7HJ+6i/HUGcFj8wrysrgJidDnA03
63HeViQ0bKgHAbWFnz1bQU0gryDzC9Yjv6Nv3Zfb1GdJ8F3k/6fb7OLiIeM7MqMwvpDPAW2vmE6O
QbWSLde1b10d8bkFIMNXvsw8vNOu01z6IZIIXDnWRLN05//b+fi5Xbo9F87JHOo63t2uaMQhnkGM
GQ8M7APwSjKDE4IWwwqvvZe8ZbQUYrlYS92S59AwZM0nfSLoMIHY0Tvx+1QrGjy1UAbNdA+lLaiu
9sIkuOefY9aZfYxzhBgW8e1mrQvz4Viot3IgEbDWDH+5MR8Cw41afGOscZCmxqipSF417ytD8ikF
nLf5FOYhhwWqICN5D4ZTeey92nbGvKQ1tABSBxE11Y728bXIPGzXGnFjdZTGp6D1pibB0SeFLhxB
AVK22hvCJZgPfPdNL/vrc6IGXL6ZJ0CplCAw+7YytznAT2mgLYZ+PkiLUDRD14+tGxRvNQ07AsxN
+yCv3vU8WKeasPwQo2It3d86yxkf/yV33ceRLmb8wniz4/V/nwc7z0RzT8m9dDKJ8PVDqjt5V99n
oGa3D3tcrFentVqTNfkR5Euq2vEV613Yi3bU4rwW4ok5tpXLBudSk12/PYLy1v+ZdC8ojWEUzHOH
sfhXVr2dk2zqR+bWeuQOE4Iun3ONM0GSfsCwVcNHP7lb/AOzsUdZXa2oPBwACU5KXYQcBCIakECd
iwlymwv8qsW+5NxXDWKWzkEJt2LFxk4QMKcFMncWtYA3VQegFGSS4mkZkmjqly926GVg3fBsqdfQ
haebf+Gb6OubrwXWb2iDgT3yKrqiWStQA3OoufEOEiMeFDQZ4rAbcP9ugx+8ESmft8U8icXthm51
8Qc7tiTKqlrTt4LC/nRl1gfULiOq2H7kSi4uRw4jcGpl1Bt0KV3ayp47VWAn7K3XQebg5d2c0gW0
2J/32jWNcyG8lvgVMz8N36dGIc7RbTk3zg0eFwWYbPtzkPbMxhv6SQjW8rkL0BWF5EF56AaGvgtP
rr5ZUdBd44ADDg1qdCXYEEUzcvDF7iHJCfJ6nXrXBKzqoS6XhkN3uEjAlnTd2M/y01Lb60qodN8Z
uKxRZdD5oCOJ4cYbwPwP5VfC0yRFlH419bxzfV3AiHACk/Jc8jHHxNjIz7mvsh53G1eF8FRgm1ui
+OuJEmzf4/BwLqyZyA/ixMl84hf/geqb8cHP2Hrr/gAAmxYmWaNMIC2w9Bo09EDDXWQdz3YGeFGw
zWi+MMK6xaERM1K1zbdkzlde3RrSQ1TcQuCshGljX4SN0vQUnw7kL07/Kwc2hyrfj5rhrE2MWHBE
kgeNT9Zmd2PiDwCipxXsi3ilKFccWORrixDhWXUHS+vsuippxCcvY9rTov9gllqXNFZXTjTGyuCu
EFz7g8rZsN/5q0qyAH5pVjWm/UTTDJ9FabVvxoezQfNa8Hl5d+ATJ50ZOacFK4hjTmIRUyhv1bAr
4Hpcw6qJdOHQPjaflIXwDYlJfJz1663JXDU1+NSCNRGd3KYD+rtlZt1da7wsRlZuFbjAuKIr/jnB
Bn1a3UQayojFD77TIdthT95GUP4Hy8os3dmNDxUBgZtZ7rfsoq4msaXrlGcXafC0kmpZiL7Ftcrw
/NZ1hXycbC7BqEYODHSNFJw9TL0ySmRqLiIX+ztelmwMLDESZLTGhkyNX/2Sfk2N4yrH5h14h3PM
aEgOdFgdNSldPjacn+aDw9KJDkH5uehwWrmIJCMUIR8ZzRk3kTEt8djJsFMjqeOP1Am7/bXKqim6
XvgGI186VGP3lBAbx5LGdP+mnLnWI8Vl+kL8ACmOXbTFORs0j7a+HqVdfu6Kk3E3lXTtIGQOKB2E
t5hrLnV6K+9PvgkEijDyFJC7WCwm8Ppatxtme8AHnEDX6nbydVrir+Agsw3zv3qWbiBK8pRyHZYv
tmjQqX9gSZvyr5Ure/G82qbd4r+yM8U7YB6m6s1i5uP11YIXXWy+v0a8p5OJrv0K2NMPtyqFYxn/
+hrmK6hMMXifyjfsI2ezyqCYnACKODhtlwnW28WlrfNZ5G3VwDD855fSuIwY8VLBIDeZYsn6hPJp
d/oJsFfTbpkm0VdV1EwH+CjX1o0hFGVIWn0SuNpU2q2sUhiGI1njOfCEm83j2Fh9Dl7YETjY2GKO
i6a0I5FHLedjlgqUT4VdPqX+rvtvXHypIxzS5LLsRc6SMWYCxoRl7eV3BsthH/4kbf6Sw5d57nVs
v2gnOq/hEST/GWFdlqnLOamNlt2bkJCLJ2DPnbPAei850TDNzsQvr4JqjHOMuom8MHFyw8Iz4Luf
5UUlmkUYN8rSWr46yAARsau/KBruR3YDTZq1zurpmWmjkSd4nxoSxro1dy9gZAVuRbvQKzldpH13
s3iFL8BiZRbZaXrt5J/C2eQJGwpogMX2JFTZnMaLYg8guXZcmDD+OZUvJcz4F5W61kvoJJhPU2em
jPhxIYsylMcu+BNw3XnC2H9pseSXsyy9B6JVi+hGcRqETSj2YVJBfcTIREMdKxssZLRC8WJIhAp3
G1qFpMP6zpM9y/yT5LKKHi4wsJsmCsLRkQqLiigxWb9Ft7cGONr0BfD1ZlDEvizBpGyUWQKlhI5O
CdVvy5n+Pob52KI9vfnKCahg0L11H9VhiNh0+1fQbjdgr5aH7BAzrI3s8q+ATUjln7h5D8mdyJHk
AzD+pMiAzDjJ/PnHOuMEWEnmDxlbN9MMcVmTqAPV8jYWV/BfH6ddWhQHNcXLojPIcn86KThxNQks
FWWclvUPrHDM/5/HoVV776Iew/y8jIS3t3boGRyeUgcDEpjyjBsLH0GuByv0qJlslkWC7443xWhy
mlXM5T0KWd5Eer75NpLdKCjYxv8Nt2aVS1D9xaZFOdoEHO1y0Nwpva4kXdZqHTU1k9FdrXjYPjq/
NBNLRQyhp5rP62t56cYevp9EhGbN4ENvwoJbO4jR32VyVefjwysbo/LCoIRmP+ReZESn1CC55A6H
/K1kfk6YY5BhCdOw259AhWXmbD2a/J1Ws4wjYz+APXfMguQ8z6r7QlmYOIVKbHUgFBAeTpZrb7Ir
ZWYDxrCJAC5rD0iN5VEaZxblAbg+juHbq8RRIkWVF7RjVrluO5SNUWR6nskyRrck5B3a5SOdKL7l
1F7qObQ2+WC6DCweZBFVTGzBbLrQY6IUgAT8K6FlteH8js9od6qSNmeFt95Pda3rvakX7uJTJyqd
A/3WQgjHr5BdjNJX/PuG1OoFx/FerFyIcaKsO2GwaRviDh/Acd9y3TBMcxhSkjvaXbbG1MJODioN
0XaDeJMQJMaNKvPFjZJkybJIZluFSbyzxIIrJ/wmt/y64SJPVo9xj3VEoQaV3YZYniS/BEhGQyIx
DlgZEUUnkTTyltNq+AcMkfLPZx0we4bIkxlppRyUzf4t5RDRdKNe0/hL7PDVvZaQOoLNkXL4AUEi
zPn8N9EnJwlSn5FTaotaeiMmz+W15ak+5C2nUCEeikleIpfmuoYNhTIeJONT805wzf6kKkP3K5Ax
IMazgXN4aOcWPcT0OdUSnJa4XebE/kl3PEAXYQdkmkFU1hkEGkq4S70DlGfi37viZywKKF5Pz1j/
Q9OBqZvlDh4sNuaDFRynJAXXCmutI/PKdWJFHvErXlsH3r/OJJfG+Vj0QF1Z7YlPeBHk8CDFSwfH
s5uFiVSdw5/Y1o6x6xcw5H12vlY8M0rMTe5nh7vBunsqUAVlZcwseYcZiHZ/83UdviAmLjFVUPpY
0qgLwB1xFKt5Vz2Lr3iayZltUFbt/5Ppo3aa6nrMjGjY2dE0nHhV+T4xf3a17TOPQ8gI/Oh740EJ
jfm6y7ZV47APgXNqKkF3vQviU3cOBYmQ5vBqZNWt/cmLnE2PpIIDn4clVxflCEWXul+w/D/n+CPD
aMtgZzIy1LDKNCWjGz28uuYV2+Q/cVaykgVA3wAgtHmlxCsxa/HjL7IeROXeQkxzSMzQ1cjI6lbO
W/4MEsRqHYKuir8SYv+8RUhZB7B+9Fr8UsfbAbfX2+tcydSBn8cir2X7kKXjcQetUavkhVomHjH2
jzecdclggmOUz8Da4dAP0gbUdhQnf2ZedLt6HkyaTjK8SPZJolir5efxFHkqrJBE7ixm3eer5X8I
quBBBn+lmj+bhw8A3wgcdg1RsSlKWj85qDjZovJ8K339Wi1lrzXq/WSLpcd/EfbgICuHHyBfehOQ
mnlDNNi5EOzphNKVkJ5WUTPYUktbWgEqqVO5c1+hkShuA1XwizYw+yhVfSkCZFy911Y+4YimxeAH
S3wigU5tFfVFqsN76Us6yuDx5mV7zR5DjwPN7aanA3I5mfqdrG9Em6XG4Hw7MDFLBP9GQAZdSdGE
aLqlvf6bPr/ysvVWcmvClU1YPDmvYYls/ihutciVY8v2yh4vbmuDEAyA3IZu1iBFE/Jk+XJHoHx6
3VijREIn7lJlkfz6oxtSP8p04pBzrEJGIUFtY6ZW1eckL+PehbNMHZiWUl7uUhFM64193jFb6qLy
wwUcDYXV7ePc7JkD1DFR6HHJXuctnWa2JvFGy5g+f6rIZELoyC7qPOwYubmj40adpfupv1Glcxr3
LRWd+r/qlLlTSCo1S0qGgNGU9RxEEfc1RMjXKqrteDMavLHlXvDW2zrhgs5Lsj5U/cvzsZm/HEPw
W2DbYgNwhcZvIsYhoXb/tWy5JJ3U4CMxnve6ZwaXgGmL+8LAXLA7hTY7NdWRxVkWUqqBD9s1d11x
hA+DIi1b0f0vAHalAlCI57Tx6xcnonU0/Uisk2f0VqDU2AkXNIvglTxma7UepeQtRObJH/6UkcxF
Xrldcdzhfa6P82uAdHqHA8rO9WQqGbY284EFGEeJ8VKrEDdDn1pl3UL9HyBfQHeJVIpw4HrwE0ux
ULH4N5KyO3OmZT7Cb1/MmWukZsECwdq9tIIo1t5gBRsBFzopYMhNoPfpGsEw8LIEmWsJYVpxZ13r
OUqUu2SBfx4eKu+i65CZDdaf2KNZO/hnoaQecR8gD++GEGU74+t8rUWd7zYyqYQSdrmROspSluQ7
wsB3T48/GTE6X8qLJLraz5gRSSbgh63k6GM/ma+utLOsPtow+mNw0E8nWlYIrH4NSPAuj7NHbt2A
fylvArug6rSlsrJjeq4IP9F7s0JODiBHtNET9iLC1sTTx91Ya5tiyInYoRnsU0mK3ZmWMDLOQ6RC
P0M/qbvgsbcOEE6PnsnSBlM2PM9W+Dt65G6Tyek+gaER5WNkYXcwY7rPBO2iGotANjHA6Cy4/vXN
WsfKTxs8E3zS6ABy4P55+BtC383vTRDGJFmWP7scFQvOMSyIfyhKZneW7ZqfGSgnYM76I9os4EGp
OSafpTuvB9eY/h+BL43irkRJuWSUeGW3CiiT12ZAWFCX3ET9gkkYWi9zy65Afj7MB6Xt+5FH/H1S
xgdYTVY40Jpv1FXnr6LKgKK2hCiMZaWgbmHrqaGmhGx5xo51lRHBG/QyrjWA4tMK9DvrY4gOMvf3
uQ9ieNZrxKRUNZDnskVgybZ0oebRaLWuDz/x/tis+XiqhhW6lNqxzsfeubUoEBR5SZoIDPbzRR0i
Txu5ODmMhUZI/vhxdoRLYlUa31U59dlRJFF2bX+CNe0uqJ7Kktuvf6JLjaYoQAqjucg2j6Q9Ar+W
824vfJCbUi4q79cDiVCnVuS1CbEhmI8eozBK70uc2N5W5LyLBU1aU3G+SVbD4jQ8+IQ7vYpLOEY4
3D02oGmV9UGVBmSUzY2sV8/uuIelNUYeRaXoXg3f71x9bn0q0/XV4QsL0gW0btUcV/rNl5JSF0hH
YAQqqeozmB8RcrxK4BQdROBRxsn6AZBMBqcFdeHgM0o1Zh7NjyGQSSWjYvTasOzjVs0qSsjSGZHg
yEMTyLhXA1ATe8dP/14TK60dgqQzI/sD3D6ea0LRJMfdEUHCqShRHN9l6KL8HC2MSvFGOqFYwPOQ
q9xVydfTrKCCSRcg5YJrNter2hQbUCZqfnXRHNMADFM6bwIDGh4SVT3J1D7Qez5eepznqAIiXxrU
qV4uAfuxa5RU36fmJ57rfc4GNyx48OASz+qSoKgpXVAyjnp4VM6/ljNqFnGU33sex6GHFjj6L0da
PKZVqWY5/b/v+uzFniIL4XffFzzk+xuGcCSuYOmpZtmmdwVVLCEjgMnxXc3S+TiOGd+nE/ewMGG0
cvMxcMpXTNxGL7YJREXerhSV6WQDe2q40EbOExfHRbYhvuICw8dUsxN+cek9/ZvC2KOi1MhsyIj5
DJMsIZYmxlgxIMy2w8G2rdNV3oHeB8Y9rkZ3316prG57Wk1YYi9NkmOd1FymQ5xTflh+Qvx9F2tm
684JXaalHDXbpAX4Bu5FdFTfw0VTPTh5URyUsPdIratPHTQcG8YPmKwinB1pD/FoTIeM3ZMn1Tsp
9sCdZDT3QbaBM0BUxi2ebhVJSFuHe9rLYRQR7KE3jrwp5h3ExJpAd27q3J1qPqZpjSoQCh9cS7KT
BOP+pJNPQqqnQx1fwrnSKp1trBNb6g/vmYzjyuTTTMukQjBwypxR6k4MhGb7UmMxOdVX1eJSmXcZ
xrq9Mb5dnQmTpFQnqnw2qZrIePCho5A7ILfHUO5As6SJxfIIiMjrG/tIadhg0pIv+dKsS4HPv7V6
9pZII8JzVoQiSdEw4Cnaz8sPgOkHnJkUiPRHm299l8tVZynk6kzBP0An4zlUPzzyBMxMj1Ry5zia
c5Aa1vPzIS0pfYVCo9mL2R/SJpIKmJwWPPWs73E+BIrg1e0H4+RJrvybd0nxs8jR0geiu3Hf/9ud
lWLKKA6/qzPxOXyM7S4U1EznlbcQmPFv1lBckoga9tf8c1PAUQFUx1tUmOmJVlGDrUYXavzcSBDJ
h0OMD3JITV3Kd0/cP9NMNiml8WCnZnUmfFzTta030edboi/gshbilYhEw6RIZwN8Y4k95aKLCVIv
4h9F2hUN8qyRAtA3NVp0b6lTD6LGUBHrYWkBDVyu709+us/gPOBPYwhIJsJ+EoKQw/zAj9HwRi+n
USo0Z1Poi5AFQixdqhn6qYy+ukdYj8r8FbOU/Q1YO/vh3YwQ1PT8aKCK0g6YsBE0t7GiFYr/Vsh3
TiXSqwI4a+FmC6MGJNm4MQZDiRXoB2moSGYxgex586ASPDJK3PLgrEigCZ+Kbb5dFYCdMPIerXJ0
y95vvwVCN+EZtM+U3qr1tTr8kBKMc3n2wYnnQvkRKLxTI8MEKvcZNp7Du3cKpprZMrcH5ip7bW6D
TwITQQBTZUvu+a3UN6wlBIVciLJHiHuyOyMkBbTml6nmH0Z9wGys9EFyufDlisKoUk+YF98QUAQK
QBIGLSRB+LTiSfmgLt12Ornto4gRzXIO8AT6S8joLEZ2kUAjGRbPMRCnMu0TCxIZrjdlbL5ipNmy
j0nNK+7ZcD0Ve4R2F3pSas3pBThDgPoUD+5Jn9AQGudOIzOYButhPWX4PwKI3CcFQYsoAa6bbEKp
knDkCqvpDWNRLWqUxPqghVt9D16Ms6/vARDKsRF++eBloA9l+b6eRHW0OzKuv8j8t8WkZlmgfVy7
t7423qqPXl7Jb2E/a2ZeMWNCOvEG2XeeI3au9nyNnLiYbs8XyoQ54qXBF6EBWhTVRyFgVa6j636U
3lyoU6k5pEmZdgHQbdESWvlEWLUH/RKmlFcRUNbAnVyjeI0VXdcgxx+aPxzhaiJajFcjnZ1i/wC9
7HQAVEe49X9IOGXanegbrhl/cr5ZA8Zd3fGJMsClHJgk5UWQGeP0b2KiboXN7tP/NanQTA1Z7Qna
vXkUH8tiWy4kJfCgMipJIMT7V5FcopYwQEBgD7rmH53zsho1ImCg5CqrP1aLN6cn8ULwU2bcUW8E
bbjCqcT1V6zoGExPzc2y7FUUZQI5+JXleQ1UdiSD8UdLYR2R8Lj1HQmXx24UxDfXV/FrEJcWZPYk
XMEqZWEL2g7ymAnDCEfI4uyoNyOEci9ZhadXa7E0lVbgESams52gtt4tlHl6U2tetI7kM+8KGXnv
DKHq8n4T4iUwcJUmOIR7hI14j4niVFK/O0HC6cV1To/vsY4bONokhX2Z+8zqqJ3dHJnhPdANdkD/
lCNM3Dgpdip4ths31GQBiUSt6n8DyHkC5zOEcUcLTLPKLibICr8EJ1FptXitJn4O4wt6vg7ZjqmN
ukAsjyTPWF8j1Wu/694YbsDPJve33INOIkdo9KzQEtzyH6fihhwbTc8BZ8095QfKAz5cNkQbPK2f
C7Gbb+Pwyq5gX/a7ejXeygIktpGcFfUcZmzOLlCO6T2U9TGSJfibp7ZTlBECutEQTQthJL7bnoyh
tSE3RA1Y+fWvKKmEnr+EZz0GXFk0zQqxFJrzJsLqv+urlYT6zZ6Y0GvROlcweIy8JK74wsY1R1pl
Pd4VF5Qv2CBz3LLEwMihINlH1828/BxUE8ZSn/XVXwOnE8E4cBL0vXZPZF9Y43fXZAOvj37E/OSG
CHD/Qe668lAgEHkdkwDZbb2qGzkI7a/yjEU3/IH6Dj7ucOFizCxfgTC78Ai50qBJAY1VXw8LuQN2
PV6yqdOZ3FtHFkchhK5ZnfJhsiCL2aCH/FYhdxL4RKTfUh5QjxjfQv1f41IL6L6P5G0yGgc0SCva
jAOsz2ObQApDSiy36VCRV441zLEbmycbTU/d2Eh4GLBOB5pJu08whe6PNIxPocdyZOlAFQfKQmsj
nPFg7XZxJXb7Nv1qjMMcsmcdSWV3Vn7mBPU6QiXzjy+Q+NmHuYDY78/8rTm6wURbiu5VVWXZwHtM
S0ocm6ZVhZkePfMr1ZYqJ/RFMkU6DsErrUzI0JnaRID3gz5spoqeV9EFxJUihed5wkcLUnqprvmM
maelAY2FLrP4+qndlYT1VW2/auzqSFX1m1pTTGsultyd0RCBHdeVVSzh5xWAPqjO5gSOkAxlSb6h
p2McGDbffHtNsvxy1lQM5LzLfYPIQ7PXu3B93betwHH2T+RYuM5B8nzwZoufR0D8r3kp3Jzs+PTx
QFHzKHrSl9NqwQryOF4MiZ9iO4PZUq7krQeinouarSjVlaGv0giAMPqXD5/AFSP8D3qbQiWQPoUU
S7OQSJPOxobutozoHdxFRF7IEbvNUQ1MTI3pc5wUA8KBOZiAZqsNWBRJpdbu0f2J2PIFQ78GaY0+
GQBG4EFHuPw6V37AfU/T3KShA+gqcesDsF2ofnfSYnGd8feKYxwQtmpH93ia6eWJxD9pFytTctLX
dZG9gXSFVlnPA+xjwqZKigh3E0A9HYTH5BGgwPDm00pG8wmbeuk+Pc+CDI32Ph6ByPLChT+xEiym
ilbsgcq7Lm7Pw5ugeC11hyy0XZgveM/wTMFMCA5PQW7Y3/JegRy2P43mwwsmU6nQnom0996zwapo
Q01VxpN0fmgZAwHBIVEdWzu5gA6IzwW3RcPPqb1b6XOSTjJWVv5Jx9c6eK2DmCJUsPGimDNN5AU+
3ojz0XhCxoOxpKujQdYelM35L96RRegVhUx7UU0WB1wkMyWjyfn+l/TmMVXgEIy5a3RKBKfuaSqa
6j/+w6ab7BMgRizgoOG2CHMNhYDUqfjb5YcrEzqiG2Ux8hjSoeRS3yfA/HlTZtB8B1O2KcD8GwdV
q4/XZrsnGsvBYgmKKgNB7/XX9hKu6/BCz8KMdH7YitqGqEsUZIaM3HX3MXbhxFa09XUBhlWQJIbx
Z7vmqRBFHO8nPQ1397AcbBeQ46y6KpXpYLFmiHu2tGQgFYt43O1GPv7R8Dm0PTGIx3nISaf2YIw3
r87C5ok0N5/9rjDYBZ66mZfDx/tdjAhKDYXVn+4y8TI+fENHTY9HszOXj1m3GQDbN7xAsxcQgG4P
IojHUMSJg4JHizmygeMXtPRauMINkI8Ub2Zr+2a8+6ExeDdEcx1/l8JkNOnRYx8YjZ9+sERsA41A
gO+EvONSip2LaIEr7LWBzPiD279HC2hYA1BibfwZq+BAxzo/cA1jH0wottsgp+hA8/pmvqs3EJSV
q+KNZt3bpfrY/o56Or2bR7uyxGwvwW9OGyMyK+xTZp9es3tUjNFm6R5mCGXMnrASo//Pyqgjw9zu
WuBxQFcnOUJ2W4Q/jr9ahEt7rPCV1kb9HBuuATVjmhWPHS6sFQyn6DhdWjsgrQ1Jzebtf1tzaABL
uQRrPKCxxRIfzbMXGxyXiUR3HHIgMl24GSwqwUnt4G+3CiJkfNCKVyhMe9gvftlloYTWSRMcPgW4
CYAM0umV5G7pynFYdzfUPc4tMjCnd9PEbqW0shyFRXDqYKAnX8eahh+ZUCpPlC5AOWmQIOcjIDQ0
wuvzxyCRr6x+izamD5fIQbtU991USCbmNpw8UgjUbmmmQ3rY3/U3N1cre+qg6Q9uKDYqNk+L31Tb
95XLBs82XPnYmljGcwcdmhP+Z0+ITy6djD7ke2J5TJ4/vjzdvqiVzCDckj/ESGmbht2UrRdNuh4O
QmAliQ2sy8GPgztrfkRwo2NdLMdUFUkUqN4o3pzYVcx9AKZ1tmgdVAzAM3vKyU5C4Hld4sR//oWk
WIOuxpOT0rjP7/t7BaPF+7skQMSxJn8uy2Xg8vVxMMRg4ZBu6gewruaXwNJZUwfmGwJBS7qHpEC3
pN71/EinD41MyL0FTm6J67fCDL4GG+uqfuC6CXmKD7THVi0xY25A9wnmHdgxfPJf2LzNFLosX4kw
FuZX18H2OUSDIfd8XkxpofdEL3cd39/uIQa/SfPIYS8x89Q/qte0/HfU0M4tfsBkad3OV7ancNB1
ITOvxWTzfE9/kWjepnvLFDU+Rdgqy3JkKnmSiFswoHQaaBfyEOSpMYlMlyh3LVVxcjKH63A9hUrC
65nJgHLJIz9YxhkrGvBzIPD4ClOLkgBBpihm4P/1K3EHvwIGK1Yh/ldZEyEb2oUA91kCit5Gbpnn
3TmOESUW9mTpY8lY9HfQYoZkdoW0vbQbbY8ocrYe1B+r6oX8xE7RURh2AxEuo1ZU3sICb1lRHSpJ
uCi+uI6uWvb2q7c2grTXDHyea+focmK5JLHJZi8vHlQnhbCCcplY+gRfysXomWB7pBq2MLwxUPhs
BsQ4eIfxUP4ISaDLhdu1vKtzL2mjt7I0xGptzsb1Odp3XHqjEreGEfsr3yxYUsGfO23XykFEkxjl
35XROt8ZAXFPQ1fM+Lvof+ev7s7v5hAJUYiNVxX6xPZrnW1ejbM2XIkxkkoE+xoxfqNWqSUox97X
SjhoMYto0UX1C+BOlWE8b6p8cE4zaFRh5UsHPPXvmYkJW3WU8d44lVY7/imj5YIhD6T9n+z0A9Z6
vP2PzS4ClpjxNLHSAt3hFYBqBNh2P4mi8uNAysitPzjohgjj8eFwK6f++2HziK86cHKR6MaKVJdr
49SOs035VYJSAKjec8RPDtyv7sCDTJVV5JhF68Ry/AsaCY3j76oZACY/WTZBZfNIaHuNg5u6E3/E
ceqZAJTs7B9+gU0ZJVM/e+mSBJFdzW7QfkqpoWx691OJBN3QYSyI9O+B9y54ww1uVXWA2gMuPJEJ
s5Z/Ar4iUuphfqskfH67nRijCbM1jJ17KIrmifZSr+pGgTDh2/bhDVXVJCIDPGI5dl7FogIU5LBH
ltGnkkPQKpwlOS4uMtElCZWXcf8jYYFNtyZjj3v6UF/Fn/gfpGjM/nTq00UJ9d/JzaugpX92FAwg
Wz0uceE3DRsB9P+A/5dWqBrEGZYr/pjVbGhtv165pTRLnVcnDMYXRiV/mF/KsjhJwUfgvjxAFZw0
Rq0Do4Re+SRKx4j5N+nYSwURkwdP9IfZ1YvL2lrzuTMdkn5LL78fa71GyIgkCStONBKQyiwNAVMD
xEhHSp7g9fqqAcWrzW4hkgL+7Is4gq4QaCM9veAjUzdgc5lAh9YILzcIuioe1AOf975/EoZ1SYuB
peiflGZeO0UGBYkwC6DaHy0bav3JGt0I0PoJmE1hJ0nRJysTQuEqc4Qaq/VsA81lPWa5CIOUyDCV
T4jhhb99fAr8RgZTz00IAUcPcQT7EelKoiPHfoDIg4OE3LHFgBO0i5jhC5Sum2C3MDEXxckNoTTc
nNwZwsaXHkLHTfbPismVr+OkrzOV2DSBnKMFy4x2AkBBHQrCgBrc+NZ6dO9rg/eBGamYSv6gJ+fq
eo+hrih3Hr/qIh+PN6MeZyc9eYXyfRh9GUcd5k8w32chMWStb5mFJFp+vczQysT32dyiShi19q9l
J+YRT8swKZLc/DzsYMCtMNlxIDjge/29PMQaW2x6Rn5DvN4FQh8yKunOxndSOTpnyLZmG4OeiMiJ
mzbfy4vSuoSumahnc2uzJQnJsPZzfI4TkdOCVdE7AvNV0+U1yAHloxbg0AH9AHJMtuVAzP98t9SG
XxZqdqVTptj4g5N1PLaSyQkFyK3CaTaeDpZS0llbmf1dbjDQ8460bFnfcT2FNEdnPdolFmTj3w3v
BYfD7U0vSXCpsQJiMK+V6Rf23wuLOGhyjoiDhlet/D7ok2oHJn0RGCWhCSBuUAnxNotgAJE4b1xk
sJ7ty00jsbllXMiagpa3UhAZUSeDiMBg59qe1rF6SehNVQYJnvnjfmt2wOMKzoSaeZfBhV2jLG0W
RrpELWTLZMDR0cNcQHKE+c1Nk2JK2NpNsKLwDj8SgmCKpy/q7QW0fcve5RE1/uY0vK5AWZC1qEwK
r7KyZmewRET3y8f/tLG/DMx6o5OT4vFWIXZ82x1/w4/oUSeVComSByWmCSMNnGwi2cyR6KGFuHtb
xx/6gK9RVUV43lEGiijc7wAggI+Lw8le4vJM/adzqAZFIHPyqSJci6EgAiw0m3Ui2jwKKGOYw5wg
OenPTsBKBtMioaO1TIZqsMkO3m6EAvS1UPFwutwbnlJe6169ndFSJstcDUvden6tQzMedRrpM+JL
gjcC5d8zdARvQOKL31yb6F2/tXotPtzauB0cKA3ZVIlHj4fgY74gVLOv+kYPT6xH2g0Nvy/OM/5b
ZRmUmqT9Z3vhM275XZgM65XjZwLTleZoEwVpqZViGh7q8o9fPnfDlZKALTSGF+EjFOGejFB73Lna
U5pj0VOLy0VUvc2en08rz7ZNWwd3M/ykqzKeV/7tdFAoy4pJqW5lwIJtGId2ucDXuRs35BuvvD4l
NQjHErETD7RjeEG5rjfITJUwH7MWxQDSJJUuJLWVx8kvp6eYPZdkD60mNYg9bcEjNail1mfPRhL1
fD/Rnyi35pVl3jmb8x6FCXKWIVWzp0au0TQ6APdHrSqrdeD3Ue0p2Rug8rC/Ch9cxptxVRIsjAsz
UQrRY4HMdw6t2kT9yoKPtIHhtMozoTfwss6Xr0CDGS8yX9CZGfcMnWKb4SoyVQIhmQdvx0t3xOOQ
T7ZtZq7V6bB2hYm3Y4FPw6cyCOpiWNYKMIsZnF/mJ+46wOggu4LVhEQzxDYj/hZdtkcNYWrqLN0U
2YoEsScxGdEsFOqMhcihyUNz3XkamTGNB5nhj9QYtfXI2ggcfRz++dLZhkcqL/CM7XzcjwFBnvVs
WnITGWz4iuiqtxBvC0qNQiT0PLSCa4tXE7ZmLOtPGtEzevny0WsB4q1Bl/fglcR6EIt9XaRr2GEC
VKqxkZVszSxMaJAQ14xNcbXnndzh4nbWJbLx1WEhuhjyH6f4ZYqm69/XqvJM5ixlXCXqFap+hUsC
JDDmZ9f/LyWQe+GNgOIl9rPyouRXTn/yauz65ExiJAbiswD8tzurhDQAmB/RpWVKKb1zJ8JUYLe0
gyT0pi/xFybZcMzf3NRMpU8ebyNswxj26xCjvbd1Gfv3oiGr2CmOBsjR9+wE61eZlLi6YeOQVjz5
Wo/O2mQtzf6/fJRoK1B81q340dpMsWOCYLasvKDwXrqkXkK+wnUGZpBbu2oaL4SSBlwH409T/5QP
8IWkUR+A2WVuDjdw4Fkovb+cO6/7G0njwv7Fm3yZxSMQ+zvwkYIB/7OorPb5aCpSTjYqfM5zbmWw
IW8x8mh6PUQOjVsh/+5JjJgcuvWBajfCM8RTzhogwzpDqtUPFZvRdZLnDFnWYFT0eYmqh9yri9cN
daca5hqxVEEtVA7fL30HHI/lx0xt4VXZhjsLDQ7RxfD1z+vxxDaEDOUh3wcDI5ci4yyFu+alN8oo
/4FSNZGTWxNWX2RzST2XdwXwmaZzsfLn/vPCH9HPTWA2R5QPiK5W1UaW6qsmaizP+itTofMtZmKV
8HKEubKWN/QKedqZmvxnghluqocyvrRR6agsXRIr1bWvgxED/H5GqlFfDgBpovKqmFf3KYGv4deR
RN2yDzrOZHv2NjhFtxyuJ1rn5u4DZ93baMmIMML127UyW+63bJYqQXUONZhZKEvISlCD/490+E9U
44ZmFSuI/6KfW5bf3Prelg8mlOLsZ0i3YI0CNIV/qi+yjolU0UfKJzYbZW3tEUDY4Yfc5fvuhuTe
vDFHnd7VgW/dJlAWJN4Czd/Wc17zVpvD7iLwtzI95l9ntNBQUlh11dd1+pHEX17U5vwpERIP9zGj
9hlNbtA8mCvNl90shEbruMm87SQfXBOiHn7zu2R8PIwQwnJGtcm7apmA2CTVX7xyKOg6ar1unQ70
gANRjOrYe8FZKKa9cFdr0IGgQAv227HpvbEXPpEsXArbdoKv58pF55KfM0XPEuLbCfFq/hqEsphO
Iwx+ja1D1CwJOo/Yst/K5ChNlWbJR3ioLl6JuduVSh9Y/ASdSyMcclNHiI9Y/H1/xflAyQ5cRR5N
jv3eUdtMyHAvAaruCeoQvpNoly29bms7jmS2DXXLMR9Se8arkJ29jUPxsGirEi32rwUksRzaIDSD
zTUlElIqCeg67tGicYsjgWy1DmJ2tKt1A/S+/SQz5gTQCELhRw8lgxszBNHYo1TwiiDqr3M000bs
aG2TAmf2iQLsnGT3iHYH9rQp2I2Xjobq2lxA7bI16PyTXxlN9ZS64cgZUudne49T6Z5haZz39sNi
ta8/8JVvd0EJ5N+17Q67oeRei2PPKs/dIBoQRXqPDaG1H9ov5WZW5n3SFKLH3LY1h6OB1Ztenxqa
kU/Bon2ZzDZRGzpKYdDwHzYpkP6o88ojD0//7z+s+lqz2u04tTdMlv+YokeNROZ2U0VyV8DAy+GA
QIeMrD62uofJyd5NJDL4EgnYPml5RFA40LQZQAnd8KxkrSUw7/8gMeEgZm406vcNUMf1gHFxrhsL
biqS31I8RzBZLvNxBHlZLRFmJHWt4WDtbCea4JwDbB5PyvrjB4Ychsz8KlP955SyqI21++ZNwTkg
PhjSYYOGDv0owZ4P1uLIX7w3GL5RSZT5xC3l0Zn+bnhdDR+MeY7grcleJQE+1JzMaRxRV84ItNKI
d2ZeEFtxd1feaU13MxNem+qZBuq0UxYHc2YxjDH1hI08gK9LaJHKqJMeYEh48RoNyBI+tnIeGfoi
IYQcYg88xEXuVLuztU7QW1XDV0XS4nG1ao/YYqplGTFOpICDlss+qitTSpANaBz10CG7EUhezyn3
WqfmACTb2ox6lBHNju31vEAHcTvKiFataQC2ayvaf7YUefLLmtApWxPmBij92llmHF1zujnzDt2j
dh1yIWSlEk6SVIvFX4mhSsAQ9yVNTxINKVEagNbY4cYhZq6yKgg4zkL+cmpfAaBUaer+NUNU1RYG
0ZVJhFE68ZDohUPmu37DLTANPOEJ/Aee9ReN6IQeldPgorcZGW423O63wuEbzhyOqG3v6wo4vt6Q
N58O2KnWAcqtVWcEIYyEa71iGPm8auEpgcVbCFzFC9CYBYVXbXtGE0j0DXrScGWaNgN2S2SDGpZ1
2DoeLBG9xAlgbAmk48u6H5TVuq+0kOaG7aTpyLO9ATX/47xKJhKMB4v+DtL+KXAB7+davDr9HIkY
K4aujbKbrz80AwdLMOWg/KDJyAcVF6VJRx9nh06J8O8x1L1uYzWf9VGZJOX5eiUbfsvj8rYM8l9c
rWaROF/ci5ewWnt9q4zBCkfdwgZhFgMii0IdOh81yv0+GMMA5ANt9KssSufwi6829bmb52sUI7lP
mYQY3WflG16FLTpryNhWQAZXGX9dE2Bv/iVTBjlFg9DSGUPUnZ9HfSn59L1DmiKXr0rsd9i2vZUi
ODY4iunJJHk72w3GFrfbVbFUzJKlwnBLJ8TOKwGYleOL2UBGzosdqtCPFuo84woVZg1zt34vbZ5Z
xce1mfl22NTHa3OHnAdMFN1hudjFCY0pncf8IwFsDddGQfYcbiOT0dRsL7HgDDQM0vSmtLv/lRO7
Os+2kFl19FNBa13IuFpwVq3xrWOBfX8b4m+Zcj9Yzfsdpx9vd7PppaIz2xuA9b4DcUlqw4DNN/K5
X9zUqxdCH+XTxYJuN2MwNASJ+h6qbiV1PgtgWai9kQvwNpipHhMmSrp/54ZLeMzsci/cjKDy7Ppf
ild3nCZmKnu0/ZzxIhB1BLAnRkhYELw+9BnC1dDSa9dKZWFP3pxktG/voJwrPQPtkTMYSsw4sTE4
82Dgx3lspltOuVPllk4qXq03VSX5VKc4/SWv0PPTQxLvgKK6ShnD874/eoJ5MNbUjJUfpF74sekH
+t1ctf0Bwv4gG8T1uBhuqgv30k6jE5+uuuC7x2kZk9j4EmG7rUnCXmWcZXI7beEqgnAFlgx8sXCG
++FNpCnKae+DVDhmNE4pvlumPvrV9ei/jAmdcwY4kFNR0jKhAXznlAwmdfqnEgrOCDPFDF7lBdcr
hUmu4l8iNjxOUTFG0aOJa6vOuuYtBBsuWvCkerHP+CvAqzbyK0b8SQ1n5EDHNC+MmpjC2oRPgO2x
RhFjq1wMl5AF9S+gyeUK9WDJREeL8tm5L8Mr4zdbYosEKY8BO6twfoFknt6PoVgbJv3nB8l13w4g
lf8zDl4/HrhvQIyzWxwoGalR2lDSHTh2khvlN47uCAkg3gcYpwBlr/LMpaEkgzDkbMA+lSwvjH+P
KIPqqG31R68ItLtyXhaSGNcFtrZYDqympWmsBslBXnjiZV9c2tSP3zWbyWYI8w0vDoD8hTu2fbTc
m+9eeN9l/lNN9r8Ezs+aNbroRgVEbnbq9kQ3p43pHuUMTuj6jW2FpVjWI9Lg9QHvcpE0x1x09pSJ
iXmtLr4PbZfVBX95EjqLyxNkWJ3/kTTIB/nLr99Xn0QlFDI2BROgdcLxhrgsTY/5iG6HRlC+uHrm
/PfhwGB4NEIgv5bYByxshf7vXUh90CEz+OUJGSJd4dowX7M+TQbgPACbqmG9jrdhXIMc1Opb3jyo
w7KU3ZQHlvWw3GlkTYmzAsJPp162ZjhMO8ewGQXjlaKd3wdi9vcLPEJmtrkyxDvF/1h6whfZxWkz
WEBOHZqDt1imJLLrY5Rukv3GU1dQl+SZQ9DBb2CWTfTJGXVwUv0tNUJLL0U9i7QFnWnB0f/8rGjW
Pg15RgXxlqxGsKuVoSZMlvkuziE0fncuIQ4Cmss3az+F2tqJajVzfgbbkbbjCaL2SdiQYacBIcr9
XkgkZBE5Xt3LcBPFu6+WLc0Reja9sXR9ViZC4VDCcJq23UYu8FhXwfOFubO3miJdmoaP9GlzQ582
3qgoAFqPcK8LMMzgtIta4KWFN02h5ZQzn0BPrQsa62RYGhP1QIBzbhQ6FV0xL4R7xgRN141XYjmJ
ORq8vlWnI15HcOgaptrnvYcu96ebzWAWCkTIduVsV+ZBnQ1pGKyD6FjHw6yzf4cLPY5j3neRliHT
R2hOzN+Zfgv0D3oENhtODOcbEt6Wr0MGyzPHCN5iFNvEJA2+t+IzTHQPu74l4dxMa2IsiGZB5dmw
kA44pAbMpUZBqlVdNjCt0zbu9+4oqbVhHLOSWgitM9oS2Ib6TjS3ohkkUqdXeChxgWocgY0mOQbE
oXON/p+B72MaoIaP2SyCq46DXh4cHe4/saPdRTDkh87DGRtR/5fe4ZJ//eg7mMi4N3HlZJUqSuqg
O5BFagyp+MyViYMQffQs9lNohY9HBLPmQR2gK6sMiIEKEP77zUTmqFBoGSogtRdLQYkpKddLgtGq
SONnaFywymEtH4247Tp8vFjkV9FtSX8yq/6SfKXgikqM3KVFaq/Y/jNwuqsOsimmDMEibOvJJuc1
InC8dP+0bJ3vCUmdHfuheXMx8pI3+2aHAjebeYWYn2lXj2sl0c27tI2RUQ2gSDKH5m/32w5Ho10e
re4A2Q/NaQjEvIJ2yulEU3G0kaCbh+vofShVsLRFSmTvVaba/0hx1q0euF1258AEyUbRJP3Y0bNb
1yl5rjsJA22CLr/FPQzRsi1C/bkFYAojd3rc7PeOWg0wvUlc7TNXQWq8zx9cIhPWPWPjM2Eg1htV
Ofqqq4bl/eqfdWhlwPgk5PDR7I32Lcmm1xfb0rLgdd4Wy9zIiePQVnUoKdfDzXVWBJCb/S4Qjk87
WngPVAawGyYX1nCKCKeTk4ZrdQuuumwLOo66JyIxUOKQOFOBW68neGfdqH7V5VvBPjB7D+AhAJmL
qXs7LIcIBDRUscU/KuGah3XaPr1lhuOiCjV2DjfgaIk9wGpYzO1X5x2Adt8ri4//tLhW1/JggnZR
siWlrVSROSv08zQXCgDSa6FSb2kHzcjG5hP2AcP/vhgcVg396fOTAAGBTYp484uBj2XQWB+y//bi
GJg6DjcVoKUMhYEgIQYj7dqsaSwu+k4Tms0rl6IeciucrMlQ9e41PuNULt92L1nwLIv+NqSyxiRI
3rGco7EM2A/2ts2h+D7TVRKgT7GN3eAYLaPg/cVsNYSU/w+ACAxBpxU4UX++GY3Wsk+qmqp/Havk
AaLs2rCeAONowB7+To/oatDr/jTo66cBowDb2xaPKjys4YvpbuvGhIrMl3uvyQ2AUOxRMoqtZ+LM
1J+R4tugkpIVsw8OWBRVcQq7wF0p4TjmmadODUIGLJ8VrRMfvSC1bGHSl7JKc/YQWFfbX4IBM4vm
g/G9HsDCd6g3ThuyqhcmvF6Dir9I0gqTO8WpCfSLwITEo8SZDmrxcZZHl3oc+FEliPMzoFA4u9/f
m5rqwC1TgsXWWHnQZJ73NzjDiB4i1EdTWrx1c3z2MDX5FI0Pd9NuKD4b4HI02LHqg78xI6kAeb1y
KSE2hTjrvaxqgF2t6iGHKeOPO/2z1tFhr+hRARXt3djqxcxKKhTMKWUssNW7sXvIkN+kYwfrhlzN
o0t4Ci9iCX37/6QGMBdKtIqDNCAYghH64sm6SzKiWFOMYpVLKCI7/aDUFC1aiuCp2d/NVOXhKy/B
kgNlQIGaO1bZN4rIgzAbMIrVBpbfRBFdzOXzkkzwsJvK5Uzwc0jC8qvVmR94EdCM+jX7e3H+kzz5
Lp9V6aM5ldRQplIhmMHXYdFcCLMW+zHwGwNFd+lqQoiklsv2ZXn5v/ECtLWxphZgMNoa4+iMs20R
iggG79+21P00AwjfNSOC/lAkLZ92I5QzU3o/1esSBj5smdqHt75dVX+PgfQCCwNQWF9o4u+922pR
RA7eI6a6XXItriUOuennSyZsDdCqn14tyC9dQOfsvzvB63Gdcq7NALc6eMUmZc9X9WkcXJMUWNLN
mGrOVtC76ysuETqBWncc1Et3VuoXH3Tl1xCeGG1AoIkhqRBzkcP4bXGrWYaBqQV7NdTPK8gVFHzy
ZKNYmaiuopcR7eM4vjj2LiKroCOWrvlCtqM1qXtS5+lsgAxwk8cc3LsWSkKLuj8QhQ0XMqGx+voP
/Tc9Kduynj1s4JcNjGArpO2c5cJiYXQoyAH9Q04UFFnmfmpjPHd6vdYRr0WBQRSoGXeLPxlodQBZ
Gc+HwpBnVfx4//MEyAG06JM+4mvzty/h8Got9Ix5TTKldh6d2XTJoiLP03zFtQ4xkDx07xrk29xd
pwFsunzqx7VWHPSD3T3AM/duQKMOC5H9BT2ShgRhnkl0BA6AOsKosKF/M0Y/ZmimNAZxWTUP6uEi
z9mSBD53TBwiZqpYvAGtHXhk8bV9XJo4EoMkht5oc7DaPhBKNKSyiBsQwJAZkqkFIhCr4aJqFxOA
XTRaoPKmOHtbAvmvAz3osr8wW+9S2KXv1VHgPXZze/BZJVmFyBmTanvi0T491q4CHl99G12Bt1O4
eskrH55ikRiLTV6BjeqMBGQhkq+LhqbHelq1HVtTB/1GdzlPqrolOtKjpQZcfT9J8GKv6HHanTDO
UdUWk6/1WeDvVdlN/2XmXZ9DvRLxGv/GGDqvfm/y6hkSO1SXP3fZMOv0iyLdQJTsyTk6d+1iLNp/
rm7DDq4g3hKbW3gt7vNEu0/Xn/GwTppdKWQEdlqhGeyt6iH5v1ueGqug2QtwgGvBfP77o8wsQ/YK
8+weNgVtxPhDMB3Fudbc94fH6DF/veZCSj+Dwd+oyPAr6pVe5y6HDW2O+zxjw24MNIxMt0E1Zny5
sPs3LpoW93GfJcmWDmm0FignKZezfDQ71gknneqsevA6W/NFBXkCizazJ+xR1/3rXLKTQzs8x/dl
bONhHXeFI8fi8+iuQ+ZFnfak56FelYIcWxvYPqNIFcqxNe64VqnJbGjHIxT5Z0SZYAnVleIAYiHz
5pb+RAzprportCeuiAN2gdu6Nj0vY7Omt58wTwi+NSWJqHf5n9Hx0owRl0JDSCOveCa21zbAvApN
sHy4GPd0XV/rSP7kCMHu3PuIRv1ccK3u6aG69z7gfLEbh34uogqpw0HGr3m2dhf35yN6KU/V2oG5
CI3iKi8AJBbK+fAt5iR/Z3jpgYdlMJ5OaNeWp7Pfgk5V7jH/PKimn+J2/dD2nADcbo8Bfce2ebP0
BUvw4tTY2iIMy2XJs4jHvmlwOMQ3V9xiRsrhASMZZCHGP1FewKisLSlfi1Dcb0iu5CRWg48aNIkP
33h2P08od1TroOxPR4b5BLPZpCVP+wLN/1D/5v55blOEoOw/eWy/MXhOHnqOAJtf5zpWDurG1EYg
0A593KhnfsitgILk5ibXk/HOfLgJ9jnXsIlFwcktRDzonn+Fq3GJX8sXdkxwVdJ6CULNIkHz7JoB
HmS3bNpmCXLEnEL6kVJeAnAXjpsUly2FPFn66KLl4PbnKRJMD1yYqwhcDmCUrE0Z660KgfrnO6xx
USxt4Lz0Na5vPYUOjrz6MBqD47dRSh0lEZbt4U/ppxVdp6SRWgTriNmavd3jwDsnHO1XVLRQc/j7
0rXq/NgYQ+gGxwG9WFibAKpZcShv1veLOhf4tm/vzKn/O4c/sTgljfdOT2Kp3Kq5Gw37ihxmjCAb
61htwLZIwNl2xcGsyss21JK5ePugXH8tS9rIS2VrvsHggqbtWKtNvHjsHzl0LaasuyhlWeT5Vzu7
Qf20PN7exAqoCCcovnA1GmhEQIEnRCnXOx+zE5LzaQHl7r6AFgnfNAEyLXbq08MIrtsrdVNVPlhd
9TdsJL/c0KzOBLFaNd+ocOBk6ZMQu1Iqbly2uDoziVZ5HHB3FnbNxeiWFj5Xmzlnx1VIy6vFyZ1x
bDNDx4q2oCBpiFUJqVr0bLF012bbB/umfjnUTyD4nF+0QCmm6zMomddFW5IpNAgEO5ygEwAkgbSm
yIkFti/QVXHSPsXdp5A0M65ESbAgiKlKc7sD4d6Z+WbULvUY8FuKHae77yv300PU8ul8JXf88gGz
MPQrERFK1ntKQkyvGPrS6ChCtqucvaEOPjL8anXKQykY+OyxYebMMQQEp6vV/gHVswQUsnOF6YZw
8mUey68sRfMNiBgwdHSJ3O6J0TWaap1g3rKx994miMzlJxomjPcW8asB+UGLCFklN8G4jUX8eD+f
YeyzcTwWtw0qTP++wopF5+pDR2fLmdXdkUQlcsIS1Rl5ZQMTVJCe97X6XVntnBXrlnDs7trpj5Zx
Pt7p6+7QJRQB7J6ndzGE2ZJK21Ns0SX9cRPtUYX34zEEKsVpik7eKf00XySUTocOd+O//FK/MoeU
lwbCjiOGlaR+7UxtDo0U6XsUOovj3xcTMFahgdH1CDeUpu+5TCqq/QxCpTffpYDSPmOBdalAGfSf
LhRGVqe9fiH2XKnqp8QE4aZEqSbqoV+ODFwzIwdTXKfue9FcuBH5K42v2andwXuSK7OiXKTv9h5M
4MDtj5MlHrQbrWpxeSQVipx9Lsd4jXGhdSu+wa+sUyuuj5WFBUf0udWd53kVi8ZgXUAAGRvqEcw8
et3jMPTsUE4AoY4l2NPxlOiapXhCAUdlOHiruZ+mTAnstRxz2jpa5C/rVYnwhawupv4aJAzcDDe9
Dsx4SgasFNxOPb7xpjSE0seTZQn0qmIBMsobLfJgQZF+5qAsNaJ+HUPM/YMvV/bL/j2VFftUOcrm
+cOAtz3YL7B6cZtTln3+LROmvtNXliVKSJ3jXmwCXScswMTyhyOCxZ3/SsbJ1cZbC3xJ3VXmS0qU
0Og5Um1Cf4xfAROSBNhAQ8JtdNo21RETCCOC9RWAigUJc8pL5G5JMh2WyzpndanBMdSxLrTKwu9m
NhhtrfSzdR8MTUEiWAjhOwa/loca5F1mi1An0jFPQbgBn2OyrLzMHgC58I89R+lNe88tCAu0wkZE
79VNNAc8rIDTuEOooFHKSS4uHNBr9AdvqzcYGJZu9500t+3ZavgTz2nS45ImAwDPxTaKFDwUFfs2
cV+vbWxMyQeFsCl3j6JJ8drFZ/Z6wkES8GxFTEqnT8dHfmeS4d871U8Tq95zIhwHngKj2dxq3Pz0
lb0N9fWOm478cYaw2bEzD2wo0vm3aOWnEdTrXwGS8p5mTvOO9AHx64CTYEAWnUYzL+GUXyB4Cks7
9m3Y9gqfHEZQwE9n3NWceWhoR5rRYOGuQlUiiAOcg34FwPuL1KCOjViFmL0MmaJzNHMLRoHKWn6h
gy4eWMd8yJt0glMDf0GFZsmSfQKfT3MJOAfRMPfDd0oRfi88QXXi0eDFSvllv8PjVYN1jdSIr0K1
I276hMMqYXVSZZvmKyVysKqcxSL7+2pG2USfSOrosFauvTUZQSXZMIzFa7tZzgcOG+hsb/jzWdE3
SYDHUyWgd61VcL73O7noxxf8oO/tdTR1/wIif/9ZqRWJH4anhMx821/ROjRlqDIgdl4qfadRUMwu
e2mPov9c+0kZAnPA4Ox4HLRSf+iSnViRliAawyC+HFJwWCkNoCt2abpJ56T0/xPIoYtyPL6gOpq3
UdHfxBgW7O0cfrffFkKEPHWP+otOd1pMDEYljbz1yKOcg0GgaXZGUZyhoJLQobUDMHzXS1RU2F8/
QJlsv1yp3br71mvJkR1jdILYKGjs1DHlqYAX54mOwtw7zigeSx9NY5uZw4kcH12pO55xxqMCHibe
d0odBn/1bmuOChCNRQc/cGTHj9LC60NVwQ1D5i0dsPXcyojXFsBneFwEbeJqdidCVURyZHVHb9bC
sTf9c/nC+o/dQBjsjw1z6uz81i5mY9PsIJBjWzL5Kz+mYNQ/MxNnsIa7R5Gl+kbFk09WG6d/nFhU
u60oJPH5llvId8jHH6cssnzhhobxgxsP7/Xkorilnb2Y+3+5JcisPECyAExdlX7d7mUsumTIh/dI
mZtKOFeM/w2r+2DS63OosrlHr7z+rWo5nAZ0JQsh/5J9bSHZejnQ/oXYrLWtMR2PJsYkhtgZUjOh
zGJiYuE0Ebyj1g5lrNcBlpplmjzUtT+UvTEHykZpovqHLZYZ2fnnvTbQHSyQZ6kj12d0X3D3AVUz
CBg4x15ahQFgmjGo8J8qhv0U/q1X9JE17WIchpaUmryOqOn21Gw94uPGlnQfdspn0WFtftPrNxdg
2Obeupx/WNyTcwLIIttVhutzZdAacMwx+V4WwrhZP+yvmJRIN7Ob++MJO8FsS+0G83KQzHvah3XJ
tFeojVs2kDPGEvL9AVe090/Oa5HcAz8FKbP+0i/ne5gW3ivATSGEmbgaaS5pyTgeZ8yJrVLTdZnT
9yrmAzDIXW0ZfYIf0jos/xevL4aury0q/PMlIA9hKT8LlNn+/SUn6Fa4L0GbOlhFYTTyH8aCzSyp
G156S5af+8JUAlt15END5oJlHCpUiAXF618woyIr9zmfk77Q8JHulEnd+nG/Bys00Wl+EEFHr4ZJ
qUTkgox/yGvHjmtXbPzQudo+q4wVsoqfc6ZufFZO7x9CHTOBcpQK5n4H8Q6d5kd49xoK2VW2iTcK
ZmADAcbNGuYFtzRHY5WFKhJ9NQ9gW09tzrM4AvYU+FQXhj21S0XDjoH69M0CImwfPnso2YOhSx9E
AcRGN/yjdX4yIxXIxhw6ed12kiU95gkSlg2pBIPDDu/LLsocikhtOozqjdtPQh0eEUY3jsq+/7Bt
rxudpmapjB49aHOU359AWO5eg4L3mxiyPG6JfAazCVhYdXWWFzI3gLl4oszq8fxQfzSHEq7UMP4M
T5xNRNL4W8KXCsgQhwoWaExYhaPP0oKT2ouexbC5rythX6ztXIgl6GGBExdJTK25W0Q9nmP8c47E
T+klkTsI+VjNGQGgCf8qvox4FZoC1kkptvsGUtBnMbmT5AiyZLbtHApsLf2OI0Fc8DLMiOUUidsy
G1vwGVofZQf7c2EYzAxLZ7MJOnkbPv5i6Z6LW6p5HFUh+NjyfJ1e0P2HFEz+BmdyXqB0NHAoAxHi
haVeiHJT02rYx4s6GanK7bSFVXuM7DyhP6pZZJ2j9p38itn3X3o2B/fTIJgOi6i5PbTEWv9kGT8z
NyLhd+VfzxbPayJNl4yYV0kPcqRuxx00xD6SCkoDQujw1TDiy8y2m34GVpcheg1kimCXLS0VlWob
vFJ2X10H4mUgaQFFoFRsDxcMd9xt1cF5rrBHGxg16cvPb59RjCd4Af3PW+v34inVP7LjxNpmojDV
5nma/1cK4FgcsEm4lDIA0CyoENtP7zjoLKXjjI8gzy3piEO7tEpfyzlUtXad3Bts3Flvp9wI0wD1
vbeceSjS9v9SyLcFB43HbaDZEkS8MGjGh5DXtQNnntXaQe4S+QqhRBOQSBXstfDAT0qaiABkDEua
v7whNdGd7al+xHjhz1QlBHnlKCMpVqXL4RKB2R+CbCrl6gxA91n2IY3Qv8JMM0a2nZTVa00xXr7W
STIQZdYIuOUxKB/5s0Argj4Z6kZoWhNIZ2MelNcghgS2sN5V/3ieensimcAX0GV+RbldmMS3gtrh
BTf6DiK/9+tYs0GU3GgSOhWLP4697EcHNMHNQdNoeyldjO+XYfzHIYz07l+rwAy7dNcPhRIVXuND
Jn7DRO9SXWZDZgo8AQ3wwBHEb1dlGVHUA9xtKllxFEuV21T6w5YLxBGXYvwq1X3XMLnlvA4PnTpo
ze8AWuVCQ4ngnXx4ppL5+cL4eJeCfFEPv9z50q44WRHg1eii2ZYMOArqEjtE3zhVD5mo7jwEuZKZ
63Zg43oZQ2WM8/LVO7FyFXbpOKFAlxu11z5tYB06EVD0uWcizfBsVkxSyFs7tSDuai8Owa/ZJs6N
IKwoOVr0KUxJilKEsCHxi+ya61lg7B277SzrzTKwF/d3H7tcLmcK9M9OwdP+MW28d5+3D4JuTc1g
Kr8zp8AEVodKreKDrMK77myOMXu+czMv68hdzYle2O6PtfcTbtgWEuf2LmqrRMNGyGId4CaLdq/k
dhVTdc/clRs1NZYh59dKEh08vEXQ0gm872sh1f1n1ueg0khMPlF6GuO0bPjNyi+4v5x+EG/0E2/V
yT30Hd7it2MVgqvgn3/e/mNpwGb8MjOd1QqQFtV01R2GY1ZxhgVeTKvuBoDIi54PWvWjHZOaITWc
l2c7PJ6swcH3tdCVaRlDShl8uWUDgv3LHrRTR3FiM4jrNWPs0yUX03y1OdGm4+jXCJiq3DmM0IBL
IxRwI5UXPDZqYh9YP/IR+znpFlNfZkf5wq32wrjVaNEfNPSkdqA1UEqsmnadQe4YYX4lKlMFxV8G
P/PHf/p4h1cnVaYvpE8ImTv90nlcRY59ja+ZDgvgDQ4q2ZgeqJGAWFJHD5yaPtnfdsUzfGNTXunW
Xt8OLTkYN/pRz18R8yNNLttDKLe/7GxlxFxS959e8kj7bKoXWo2cE4txANp7EX1xyDTbDJ57REZ0
TlFw9t86TR/6czvvXL9yVa2TtT0pWPST3MrtFXNC/LIkJOXyWR/pSc9tFDj7iFW1VVYhUYJI6pwv
iUYiY+Ds29MziCzKnA3yXw7rhH0x1m8Evg5ysw3c85gncWZ/qLhUD2o4B8d0IBBy2WNsa8kCamEU
4a9HgYdWV/2ZAwGCPv/E2M9ikQgCfr0rraHQRmpf7OZibeFiKIYHBQ8pvSt3zgeixh2hNEa/kzo9
VhYVeLg8DuRXyxZmy52i3fn8WVz/QwX2+NxS4XWdg+/njGsZyZKo7vUU/F+fQrcqYBpVdQQJ5oan
Lvy52ZY+374pZo6T5XsH7U/8iTjaku+gbWu3AukUqfpd1LMDFK8+Nluhz+11S4ITXeTJl2jks196
c9bmXCP3JVWysxzJTJ6nyjlViNa+VIFPBNDfKgcmX6yyi8vp8kLjmvk69OOnj9OND6HVfcMAU/rR
Xf8JJy16Kt5MV8o3Shti9LgaA6FccrTtzPqv0W9shJ6UX+mCfHO+Xx3+TD6ehR0J5F7NXsOpa2fc
lgrg+9MzxAqCeMCVWSxN6QEagy9PHkJc1JRTkdKz4+Kwx3hmLh9VrhzNhsW5tYbPUY38vELZ25fX
pFyc4Bu5ntuX24UEhl1AwyN3QkiQ8U3/qWUWo9AEPcx4m+1TopxawAPSNQta632Q0PHefMVlsCs1
uwVhRpF0zsOunN10kejm+d6CgHBsmXMaTK9Ab6QiMeya7M1m4MJu7rtXaIr6k3zpZxOfmcJZYPt+
5vNzWUPP12VUDkhnWOKhTyi3Gx6w9ursLEDLI4D8kXYTErrmkTixE63i8zFp8LzcwdkIP05HoOq3
MS3rJqB9KtDPaQV4zBdaz6YT0loSTqvrmcPRAT2GtLG7ZSQFkgvtZNsuzuK0fSsDJ+U++ilP/uXS
ukvthK85Xn/5mQ5jQADjLZLbQQfCm2rBv0kELFP0ZBdAGRUHE1QoBLLGL1/AEHUj7Ptk08vH4BWv
YyGtFHwicWXq6kL9Jal9Osfu/KOokcrUMYEHz4I1a4vv11yegaOlpnjuMtr818rH5Q2I3FE+o/Yk
irNv2r1eyIYJgNbOdZ0UpNlbOAfGS00Bc7VccEXVtEgTtT6NHx6YSQVcln3kPclM6lX048G2Nh/L
SNRbkwjeWCECaJJA9RU1Qy7XPNWzu0aamwB76qbunf3t+mW4Sj0qcXJaKF4FSOcsQMIOLEexIQ++
Y+pp9wgoEYZ0FoQrVzSz1blreO5WUnlGW3TrsSQI2XQ02qdMtlTDnUbPyNs1xso5SEl+d+u8e68h
H8lKreiBl+1Dt5FHhekGrtmII9jW0SYQgGsUwOKlhCiLDMfEpLWetbYtxcp4QA8MkW+9JB9XA6k+
af/wOQL/ASNMHpHlbMil856wGLjoGCrrFMlqYczHzy1PmFxOmORgpsVjnjfue97huRHHwSznckQb
2S8JtWhGCaLcFhfgzgz/x1alHKKfRYMuxfIV5nRmKLPlhu1dJVHp6tmgccykU3q+N2CefxdvhJVf
a2pyvFHXMOZQdW7hlNdmh6Cmg4twCWc5PGge0N4lANZEUd45MlEpf1hVYiGmSvv0T+dOuqHZTLlS
l+ZiHRxoJbNN92F9SOlxZdl9Ge4Q1puLujCNxA9jZ+Ak2XNOB5PIeBLl6H3jh0W9rZE02WRlCfMG
iqS0X4+ElMuPhmco4F1sioQjnCfnt+VJP34DeMD4RpX+5dojIzNfTRStEpewIGQS0n1npEW5WXEV
O9VUCBjxTZd2sPFMSt0Ip4AmgXTtgQAbG1HlMo2hhEQUDVOIk0WTuyLy02F9YPkrwpLfWavI1mdr
+piPLU0ymDuFuFLpU1YxQDY7okUKZVRaz5wHJbJF5s0FqPwjHtnjwVnThUoM5tT24DYALXbrWAPP
teRxoaKHTuoIkLbNfwT4BzrpU+upqblEMfCWOsDbwkAdRJnF3z6IGhx4zEi9XvFSsqMAxk4X/BXN
gvcRJ0BxOClm2FuDWkd5XG0jZLoumprPNa3kTsNRdgH0Selqdh6cKEGi6PKYJki5YWakEIsdfVno
UnktARcIJJzeiaRon4ctVK+0rxrfUQJpmY/Iv3GgASW5wQzLIF3B3FPbIRPAIDTz1NvlpqpVQR4O
qXanKQ82DA4foK6rE1K7ELM4Dh3qGHi35FqGqinj6Ucp6AUtJZy385thdi2Ccou0h8RXWvSrfbx2
z0lBSi/201HKsC7ly0VacJiPVYQtiBjN+2trFLndH8o3SdnDWUaxkIV3qv6Bg6I8ina0Fth1Gz4e
fO9RGwR28Tq2SRMGX5BZ3JmCzNGNB5LK+yKJSFdKvttwYSMdNGY/aVPt9tCV7bnltBdWfY8yJB7d
QjjAjXcru2dRJJpHHre99eXTNLIQB5GsWoObuf4eDSttzCrVOJaD0+hgNwyX6ZbaBGXadq91bnwh
uCwbSxqlXFDosJwQOB/pfFmYAfx1AAxE5aBWdbKG/QVSfoLBl/27Af3U+p8iUJkabb5upBUgLILy
k4CWYp8KWY1AG/tqF2IixRQFS6M+KMp2UffSba2J5/AM5qiYiUy2xb+3YKDXFyMOYm/Ef6BapdXH
gSIvJvgctWKkGPhf+pchRMHrNjNs9o8BRjvSGmNZBTVre6NkjlsYfpYMWP8w9JZYjAzVE46Cs/Ln
IKQOBZXj3zUjFH77ymm1RJxmhR2dOlUqZ5yTyM6Agi99cvBXj1cckEdPS/DC6mN4UHxPQTujSySR
KMqMDhc+7kObyZhae/8RI8pTNhia0n4uEPFpyR72FpqU0IUybvtfyBslE4ub9kOGKCpRfu5dnIVn
dd7AIxTY8tzd/uqtUf2rSFqU7tlhAEr5j3cD4ejxv4+w2YUkgIhugT2Q4u/HYfWsX+GlI8x4E5x8
pn/fWGC0TgN0nM9NAdhxRm0IYWDeAkgr6bLYWS6h9LRBqtspnmYWlj7UJJ1znR3eNm2JDEzxKar5
WHE3uP7LmXJCCWYVVoH8wvGKda3z5gDuGthsoEvnS4leE/To/xdXYMgu9uOyayx6E9lbQlomZRN+
Xv+/T0KE+92HmlvLFqSV38PL+sx3Q44Y60QAG9Nh3PsQ3643y/+07AMEcL4v7lMJj2VAiwNdPnnu
YIaU5UwrLwPlIIUAwX35DU086Qi3R2mDxTSQU1iIKq3iu8571ib8rNRyuWu5eVuE64GBXO9rDF5t
A+imb15YAcXGlGru2sATavectVd+k56XQM+DSDgACV7w537HEfPdxvg7i4ZT+jq+Tt8CRN58LbnQ
EHzHbcbyPZe5Lbwqyy06C6XhW3f3Xv3D+L5Vo6lpqd5Jc5thda1LK4eAxVmvftMJAZ97qKSKNTss
73mZrJEStUf17P/lL+65bNvj5vPOws9SKflXfhlcUh7jO9LNT0UaWKV7PD8mcJoD/xz4nfHirjGH
5KOugj/qe0E+6N+e+NL4W0edowmQT8HRG1GXmsscH9btr6mpy01RSO2qoNOKwWY4HnaCUbdzPvP2
wU6Z4IDrQwKbxZ6AQBvAJwl1E6lj0UC8h34iPOJ9UqAIjeuTvutYnbRqCheR7WCP+LUWepaupTS7
WX9lj/shZSldd1g6lmU9mGKS2qrA+WTMRDlY+wBy1dRR5RSuHU6JzKuOWhdn5cuhxZqZvgzSeYKV
M5ytXXyBQywBt/ZcccJxPybWUu28rlHt1bmBoQzKYzmUrpgvjTVu46A3D0H+hoaeDCzuLIn47n/e
GBZ8ZewBfe9yn3XtmYGvI1M3svRK3jnmbG27oDk/rEi7iOSeg7MaVza2TaDxoMZEh0H+mJn5pUP4
e5CO+8F2zIBBvDnj9Y3XIP6A7U05XS5vhyOn6IelyAsUYLwrHj+jWKP5hYgniAMpxsYHAz+14UU2
Gxld/dS4BwjmF+MuXymPCvoJkShMVZAs36Gda4R3T+M+A9uk7acxLSZk/BWWKeH8m4kgYW9BTdZr
coJQfraGe4ACWDtIeEjmvPXTIAjLLafgn1GzpVC9DQufBh18K778MR1oRdmFZ9LRpoOKDdt6x+5O
XB4CbKmcz0PKmQpy4LZ0x50O0L2jlxcCxSuDcn466qW0nAzeF87iD4yAOhYajNl7Ipf+yUjxoLx6
kfHjJP20jQYkdNkg4l7CQK2uLIum5dgZmL7xDY5zLhM5bcoQShqljjK8JizgE6XO8kPFDyzqCBVO
6+6erOvCrvra63PUt1LBAWCvf78wyMrYLCHPv9rUMXvIeNsMNErrNW4y4XL7EXY955jbhznNZd7K
pz4eNJuR24GWJAJ1ad4IqbpTXUjBugtAvNRVprtVJl1wyssY4FqyHECH4qibzTzjeLFwqagrxCkj
VPWfNJ5ljKZUVL98R5IsKlJ5b7FtO+0Kft2Ru8yeJ1dh3j66pCkQLT35NWKGizJzix03W7zI0Bam
0RGNSVgTMjbghaegKHflbv8aS5YfJRFJoKxP+j9rIQ2YJ9tvAQTiUgXzo9ekbwMMQF+tRbGg8zSL
mtFs1WIMQKCHIzjSDdatoiuAjtyscVk2QLVm01OAWepnYPEbZ5AdUJWSeqJbBkIBSh+m9ZRAfEiv
SVtnovTAuRGwLxvySysYzVfWchothGfKR0F/j6vyaQBuK8jr7eIDdVm//awbcTAx1s5R9Kf/AhYN
CK8r97P8ZRNuL7ogf8hOkZGSmilW/wxVth+9dHpVIflnzfs6nYXogdVZUGm5uhOHr2eckEZzwu9H
PfQoT5CdmIMu65o10Jeg6U1PC8whv8QJA2JECgViRiWrgf5eFf1Z+0qKZWPU3rkMzudUtke7wRTU
BZFdZu2VmnES8ejBUAUNro3TlSv6ZT61zidEveW6z3Vpa4Xnop+9nX927VPH/c3SAvwG4MvKARUU
PnbH4tIuia9RDeO198Mx+mOrUphi9wgoJsPOZ/F6RsL1d8RgLnWKxTk/QeBxrZWtD1jhQbel3KZn
a2xXPMBnREBQnDqyVEISa2GHWo5PmZSZrYhu9laJ4brFj4D+yhKx6na/dAfNyWKv6ZV8HmUpCB0D
Km6yoEzQQxbqiMlFKm8kNdVkJ4bSMhyLDucIQgVD1VIql5ku5zWQL5W4BGUMc9p+R5GMXLE0A/kS
iAXpNcWVBSr/vEpHT55XJz69Ef0W8OU6FRn2Qr9MCq59hGw/DAf1gnvaciUsHxBGfT1aepsCQ5t0
07dMg8LxKTPsc7dCpOFlDG9KqM7VIAw/M+jpd5bD/kA43+XuIE0F1JDXh0nwvMd62UDZYqk2A5WQ
3jAgOT28TsaiAPtv+dIC55qpJDjMCTDvuosJFxRNcjJtBDcRAWXEolqxYTxfD7anfulKufsmr71T
UvOvBnvKxqdIEwdBxrAsJclUY9he8iX7KHVA2MF7DTy6U2SskfY/FlEsbxi51dx2+1O0wSnB8y1K
iZPe36YY4Q58++e2xJMuZ197izEwUUR3g6CoRO7OlDad0FRVjHoGVnR+TjgDT1E0w9+BoDkpWEnP
J/qqe43qpnJdH5SWvIxpYLKTVqI0mBp6zuZxE1+YmM2iTouw4RIJ90TQHy/zALeh4J+IZbKvxaL6
29tbe31GyJiw4FrJ8uQgDcFKLQ4t33vgQYugd8rr+Bw2uguw7QM1bEABxXUyw1Xrz4x5UDQSTjiK
ASzM7GySJOGAkI6CxRBNS8PYGX5YD9ikItY++6YVby4408NiZ2d4RzVbTRtc7hUan9EFon3+f36q
0jAG+wGQwKfaxHCvqSt0Y8PYQnF/FMB5NUO/XE09cnTczGjPMvSKsRBRJ1yFvI/ZY8CouwWxJfrm
rP/Clfd25v30AFK8ducMZS+jBPP9TrgQnObvGUJjtEzTZfaRJiIOlgXrUs/BUYcdeaD98yD5aifw
WdRsnK9K+sU6rczm2FXS6AlkgGpy3DhBJ39W7Xedu5gpyn2fkHItTd5PhSz9xaTUiWUe/j4kiILp
IqY7XL0ZvtCOrIbMCkMJS3FmUmd6pSDH769QU4T0CoHjHX6Ct1w3OMS1XjqXhUo0ndGoTeaYWems
TODvD0/qNt1YF8k2LOX3YOC/o7sJ4GkvxsvpWtaSfc9/dSuBK4CwC9kIKhTJ2PsQU4m/6K8M/BSG
AfQkinrPfcg1FKBlbz2IRmvelWmWXvPoGvcxMBsNPoKVr5Cs/zUbdDSc6h8ClEq5dpCdaCRatcxD
ksQb5V0k1WL4WraUu/OjwgD/nE5K1FfuO8OOS8rnfY7IqN/+cP80YOgB5RS2VIC5Onfx9XU98P38
IcWdrqZReWqibPbNps4S3TZ2/jA1llYtVldBCNRTElyEz3kR7brg2r+S1fry+kdBISCDHMs2KRwH
VAHEbVnjeKyoqShU0gtjb8uWYNJqAVepbBIVbfhW/L5WWsL27wvYK9npMerBhw2OoqZ8KlyAlOXK
YKo185oq1vbds97hZbHiU2QNbZp4JIIIRukHzupR22juhCPevUdG8m/b7ylzOoczODkoNGBJasX+
k/J225AW7EX9maUDDTgpbJ/7u6LCMO230dl7V4nHmp0d8ubzQoqeA9ijASi1mn0hyMQHI4b+6Mle
Uz4nt1LYsQzYIOYQfGxBAhUsMSlsiJvfCrHVBUw0//8cMKoYc3mQ8RtXglvjgxN/ibXNcpibwKAg
5IDBaGv8Jn7vnrYL9LOzS1iB28bRu4V/mqh1kQ2Pii+PAsd8lQKNfG0xin1TffNYx5e2qs/nrX17
OqmU4VKUn2HSMRI5S027ABS6lccRI/P57Bbz/obLqSuEuIhlDovgLoG/0upFuiwnZeI7AQSzMM59
9Om8BxzfkuFFIk1mOnUe2kxVi8c6Z/zEQTYFO8jeyOj2ccR/kzxEaSIvWwbOs3IL3pZAFKNoc3yj
Ie0USwYhLrqUKpqvIx9CtL7Y49AM4T7f86aVD5/2naUhGoobIAG6x0GvxKdzpkTfRdt5p6WyKsJz
pQGRX4EyhzNOk36DoLwyk4iwlw5HXmhP7H33TAptfD/B1oZnEKAyh4VFf6OsyXfZvTRyvVB3R8Iu
IEy5Rbj4d51dXLYBx+FQ5PYDAKs+sA20d6Yc0Tw7Lcs00q5fdNbviuNHtuRNkYVOPc98v/Wbrcz1
QN8sYNM4b8vIIdIaMHxifQS/C9OxXzbH8rL0N3EogKwDfS8XX0YotCDb5RyH2ZtSLp4M2kjjunWD
uwmQ1VTZGE6i9Gn96MO4cpTJNPhT2lIi1r4/HyQeoLwMkC2C6ZMMIKiF/lF7sNLEVxDLKQrYpJyC
BaCH0a8gzqlQ57uri3BzMNMZANlSikqMFwoUpSHPdVcudVKf7JE5U8FDiyH+VBmDY12cNXPPRo2n
K0kQTCmvF+FbbjA9Z1mLcEnm2QA/uZkMlQEirpkylzDE+d3FasZ8iowXp08q6/hjXCq+xiMUXvTy
lXP+zeCntA8SCDKoWAlf9KIKZDQ+gVNz074WF2q3sZ6Ehiifu1JgwXUaCvJ5rZ0+7xG2wrsiEZMm
IMq9/9JzeFMOlSytIkZViE/sP8zSXTRs6VZIaZlrhbQKjbRLmz9fUlXTMAMs3Wo70SmP5qHIt3Q8
+qIwgxkc+g06KOAjvbwueMI7CDYgsva7jatKNZmL4XpVXpaTpwmaFb9xpc+1kYalzEsJvqmQx+cM
CJES4rkObFvhTZ/DOdO5K8DAbi1PkR/oVjhKdHcQqo6Kw819fmYox2GqysHYhfmdEsPsQ226oETc
DMjJlepKpR3pM1y/+eBmh1ON8qieGIwOk5PwbZctJXJMjV9oYM8rOwhJTVznDdvfNBfGXVVAvbHy
ujWCdc6CzOJkrtqrJxCjZhqXfhatD1CTEKZJOowo9NH9FJjRd7q3wSVumq87U0QPce+azh47Q9fl
jpYUx6L+lGl/x9bqvjnLFyUZCKWaDWKVYP00//mhx5941jqsH5XQNnKtcQvSpvYA5Ki6iaR5PSOJ
3gFIUHp3oyRBpYkbQXAcyVGtF8Wk33OwN0vStp6LjRADHAzGIpU3PS4WJdZETChKE+3UZ6Os9tap
CLZ2xeVu7jKPyh0TzZ+JGWwbZPl4//6fLRu/+troUvIGrDa2LbengOWN/Wm+8X6pHTTNhme5WHDV
jWbe15l9QRLDws0WzxmnHRnl4xCda/M3eKc0crIACdZry0b9nyJbYfLnHIXy68pJu1sPNZbURHTO
DYBtDsh72ZcuLCDuD9Q8JqEvcQVijmiSyBjZA4x+bYeJs6SvF/SaL+xvq/+9+vzDFCTwuRb05Jcm
BUtoONeTueWvx2s6rksG8SW28WXXk5yDpIOuV1b8Of0hjnhrVEiS/xRrL2mKiLNFFqcrLJPWmH0j
5X/XQJslPGTpx8Tp+uHrE7teBwtO+a9dAhwM7EiTKEgn8Kr/VEhkQ+mQBj5NyHFSRj23zcEy4gcD
N2Mb/BCnaSc38Rw9TzgUvacSvOkbDc6bnhMsO0zzYuAuPr9ApoWOSKHU9/awlCmJr0jQdSOez5LL
4eh5qAVv+dNfBqg+rICdFZy5uoX7QxHdfF/1Nzi8uoM+KriyUBkbUZcFTxSLj0vm2NqgRa0xALkd
vURGrS7laGtCOSvXe+84jWhZdnizLvoJN7Nw3+RIyM4234mA1yX6d7pV2HusD+QnvL7w22DoePy6
zEMtRXjfAnLVQ+8DNUbFaqci+om8BP6fPJ3F1MnuYI38TezpFylMcF5bXVKHJrG+53vdEms9tQpa
TRVVRdlxPtHaHgBeDXCimbXw//7NvhKYRc3FntENLDpZcTZfjANGdOiI63LbdG3VARVo4fvgbS8L
ZTnEz06m4TnlmhbibmeJLQgIMuSkjiWgXEiilV8j7NVLE5eBkvt7Xof1z+gjwcYzrJ9+B+D4a8aL
qtrysfRGmQlWc+RNAUUt3RIMH5ipWS4UnJ8kcoegfC8qh9Z9YSbvsR1wyRmCbN1I7pdS99mc8Xop
Haxf1fYcnV9YXQd7HQiuQMECrLChLaEmTScXjddQ885eRq9N3D/WmT8z90oGNrR7V6wBrTQmY0fN
LY/hEj0aEF77xIAYiS3f+cxpZ0dEE/hpBjNuozcoQ+J6XXhVfGdChVJ18HsxISOjvrNJUfHobEjj
MlTGywu+MXgX3B5UWNmH35VKTTb4VB8joDBo2RGMFEeVPfhhXXU1LO0YFSbv2YXzlBHLtyhM5VMb
4UieYKSKFmTguS2HYiHND6578HCbehyfru7hjYfXlBC5aIYlaN65wl0i+KBICXZlL+g/jgWpJFtD
zhsTMjEHXeh/4Do12/qXPnt59ziM0N8aSCjI98zPPZ+Vh3VdWNwS++g1+S/E5b0gELMBJ3mobmVv
S9U+tWhLsRY5dZcmv2elbOSv+K81Usv0zK8UXI9lKlBSqheH4wcEYTHJQwHaoKOXDTKiY2bS3S2k
VQeOxjCJoYIVPNFHOuNwMOC26AlvZ+uzgtyDzGxdpl79UZPJabbHo+eD6eFFHHOf2c75ei636x/Z
Kq8JWJHlNMXgG7cpX+ByVv4SkFCuBqcHdPRUvkM5LwpZMyfelJd1CcycXgJQQyWKmeBUrsw8ZbIg
z1BIdvRC7f18xegiJ0sZu7JqnFTH+q7EghzbsmjwhAaGTEX77z7Zo/PpCWGLXUQULwYWOShnES8x
pUPvfRpwJqt4xHj5U+/m+Bm3jZcnPg2eNmXGcqjA0jHNhHkaEdaIMf/Ky7uVm9Pd1OMNIZpUt7+2
QHigczTlSMaD0ygyhY/EZxOBMTPVy0WXBKaNFC4wYejepNVudp8SxRE+Ggrzk5qHpc2rF1loYbeo
fC1FlnPUCWwmYsCGMWU3mWe7K8Z21P/eSqzA7zA2SGNBvAMq7R+6PIxv7gSBnnolvNUppa4x6157
K4LR7IkbiLQXLOhjUbDhRclxJHsaRY0v/aW2ChYzre17p1IJJw2W26glRx2KELFuy/qiX67K878k
ad9hcmAeB8is8kqNNZJnMOrByfoezNPCjuY+Fq0q5DI3HYjFOf3QrTMYXdRrAGVl2fh/x1Kc72ey
kEVoxNrSRSjJISVfLEX/sSr6mZ0bE7o3l1y7GyQHRVQTdu+W3Ej5yEIFlEokz40xrNR7X55tJUaq
3RIRXdHyCc1/XOWh6dE4N106XvbM0tS2Cls+msJewrE8EkEY5Lmd0V3cU2jUR4wS/TuYwDVdS4pj
J8yNXA1qfJpTWa5aFiST9T6UAeOoGUPiouSQJhLno/nhqDuc7USRrjyW/y7UCAeGkvygxceRLR6q
o8nuWMIb7TaapeKIMgWaMesGanK6mDheSU0pLmqFfdLvw+A6LwC3cmjkiU+Is82eHH+rej8BzLlf
bfEBAvJERcZdbQbdJeDL08BACvzn0sMzc6TBiwjjtMQYffMZhF5uQaBpJJ+HkVXskUmxn7ntWwO8
lapfsTVSnmrQ4zPOXooV3I3aBUTwQEDk5IvINDTiWQYDutJ/p8dD6G/a5tBZLgtrVtG0GTFCzEhI
s0TlY44InRxXJcnd8F1HKOrMGnV0HcXTH4smgYnaQg87HQd0N+uiQU7DYUnEh+nNgJ0Vkc3L28tB
UjqiTsnr2WcphCve5M+G9ONi1vIRLW6gmrAbjGJBWloaFhDQI2OJKK15ZKmGdxZu8ZkjeO2qnt3R
ipUF/uPbokXWm+gMjqHNAB3LT9ekwGcs2w05iMxf9Ov9IVezptcbnA3aAfmDYc/flnThA3VnD1Bg
G8xrlN6+38lSWOvn7wCcJXeH3fcBY2/VhdrUBw6ZvWFIv3kbw6iPhiv8qvMhivFO+bhyndcKjIMD
hPQVBrjGARJxwTcjcgsI9+LSeRzdpfSJq+C45PpmSrWp/xCjpZx1rXDQjPhozcGPHoUQtnY5UVgm
A0WTFYLSHCbuRX7vB6vQrqkuETOOceOmfsdqL06vHuyy5Rd8Drl7PHOGmcDuQ4IK7+K2VwiwafWa
rEu1QWAxnLhMdMA28uIId9J6ddCL6pZt0IUrQa0xnUzdoH3vOyrV5EqvItHz2hRgpxUEVIeX09fX
U7YSzCmcfxtftrvqaOtzJTnNW/K6GuT300PXivd9FO57bropeydOTyoH8Ak/Rx5ucS5afsopwPkD
YBQ7tjSvXdV9k33Et2g/COJf7F6J0lkIp+SIIIcigtn36/mESDrxDwH3AF+RMQXcVsmbHeGk0eIz
VJfXuTF6DRJXvVPIaO1HYCpjybXrreiKzecuH96GSzVO585+MTZOPEuImFMlAvSi759phu6avGyr
9fkGOEbNF/Et+OZUZGGnoOJY/vBLWTU/1gUJ5G3t9kBxppxaoAtRH5cue0XvqLW50fNqwzXotmJq
kwlL72G21kEZwxlIX9iFikAPebWe8K/AVvLh22qd5DTsOYsqW4GZNQ3d6QmGkL8agew1frmgNuK2
3gQVAR8pQcg5vOEkE8+b37zma1k+iQAJ9kQofynF2nuDLU1s+rQi8DTWiNKpikHFPip9oKomm2+t
nYTcZz8Z6XQEGzswGFQncQlbJY/r9Cg6CwTPeKSRBkXOOIrc3/cYEWAUeabfk6wZs00UywCUx4wn
sWrbuFS1PaD/3Ni9fgiNgLSsqHmaSF0iAOttPbmSqDsGoedtMImYBVU0BJ1jR9qEv7XtLGaSZtOf
MtldeqtUPqEN4pgXCYNa1At11b4eRcUoPw4ObnPs9NWEBkenCXaE2gzlmwSXWNBfMq4E6vZD/bVJ
RGebcbkjOqp27kD2n0aN3P3cu+t4KFoBhayWK4CL8KFhdjIyZUsfMUmVCpiRHP6IxJZZj5LgCB2U
HtAtvpmB5GjEhvXFBDkS9NV6zOYiIkb4kgtmIeVvNP6XgsKiVlyhnAgamaJW/3IunJ3T+AfwlWmy
A1fl9yKht9dJJn1p8u8BN6433kDNGGItG54+0f1DDI/JwbvUOrKJgMR+cRyVvfy+Hn9hHXjOOXUm
yjY23tej3Hu3SbngW8pcM5lEh+SQWjFS9jPGVQao1RmRRaVJrZ2r7qokXdKKV1kNFygTDDWlzHTh
1Fr5cjDVjXMd58LnYqBTW0QI9r8elYuBrdQC+ip/1E9uIBNXKC5G0OBROdvegzqYyln8CYl+GBfI
I8BKDHPZV5nZ5/fGv7a73bpZtj9s+xlbFql46nDUeghZWYfP0ic0UnbiuNt4V3X+2ZOXvR2GFYBH
Vlns9l87J9MfkQixXSM2lTyPAg+jkZTdTBbuIvML/0+R1EaYz3YM8UdfzHSuoEq2Gf1dPiSMzlDd
QfT+oHfaBXA89beAX8/fdN3NtJGp6unJY7jLLYeYxvlCR9eMQZATzyHpW70es8gVrQs9/lZrGjFP
kh2SwRCMZ168TigAPPWbp8FcgRzMkbS20R0eFKS46vfsNHKdkeLO2fDfvWBGNXC15D7RRcn/M0Dq
HPo92XJo1NwOFM6oX+SPCZ5GTXoBMTWZKvqVhkyxRS1FuG+nR7GijFk86b4OYgcpJtA1Zw81megi
uNKAEwFL9kibLd/4sY5ZoP/5mSKxfoJaYXpCxtF4vWuyEMAJ7VhN6N0wEgkQ3SPWrXziJPxCtFlc
FxOh2gVwk45ku7DddFy6a8SjT6ygukWugRYN2RFWv4NMn2umu+p0dseSMWVwPnAzhKGua3CLtdFs
liGgEwI/kavL/Z/Hz57w5HvaAf/XNZ5WQDFj9Xi6Os4v7zUdSswpt2xSVTjALoaGY41YrUpL2iCY
wHg+kB8N6CyKOacMC2nzSiAVdgwsRUkHRa+nEn8djHN+eYU2+gYd/ajU3YPgh33YWAAMFCZZCTmM
t5miMq+AJpkD+08wuxQN+0daFU6MbwX5ma/+R9/bxjLRm9rxKf6LpKqK75tDorbN1Czskfx7HZ0K
4pYjaBs0fFuTC6FXAYaM/OJZ1RuRN+VPbfwx6NmeuEBhZQcHq2f16R+XviwPU9HFOUYpoAcu0Bop
H//g8fwnPptljfoC84ZpdunSjeA3Kdzo0fZWYTMGPHVElxWSkYMSbsye7VANvFCGH7B61p8HKePs
F/jObryqZeS8qJPRNlWnzcCcY2Fbvbq0k1FQuHYCObTdxSzsfGOPahoCAaGV7iPImrCJocP8479E
3e1QiAkg8zzy2OY/5sjmljSJy9qacP4I+6BxzfQe8EjlIH4V8HDFQ85EHYeowWcdHkd8M36wY+jE
TqNmmNWbw1MWKCU+wfKICIZnKfaX3zFcKFvuw/l/dVlYYf7lQ+k/J/32qC0H/liOItgRkTJd1AEY
ydNwozZmMOvHhFRaK8Bqxu7FhKr4l4pjvyCttsSN16ZKIUaO56lnwU1eStkjPQIi2sZGmqUXlLDx
sYFnVkwdjlrGF50EqLk0wXD1yxtpa+F+uyh83MpJio9FEqtwngV6EoXDqzycVu0Wok/0xtwN0BTj
MNzQaT2sICAwmPSlLo8oW6LH1v2D2W4yRJMMQGPlg746BHb+xwiimyx7P3GGfnRgafrVE7RZp+EJ
wiYkZXBpyfv4ILr3ie2LRo/m/VzNbH9+kz0gCWfJJ60SACReOoHEawQYf7sEwM+f8O7tR3J7CazX
+xEp4yjmABGqh7/1LYyk5Y3qwGuEyCwM/pJx5DCadMT7OVBy3IN3GGgvwd87JRmx/cw11fk0FB4Q
yYZeqad3qXjPylIn9agzlNP0TLHZ5Zjo6BkNzQsOrwRU0sZITca6Vg1AYU0KT3+Pu0KvvNITZxgA
YudkIRZHSW+bLyrmXztprxnW+Nz06yrqe940tSIMKy0YQcv2JFUJIGDzU0atAerusAKLlJ3UIQB5
9uaLSLEZBzoZmVw6AFZCH3fSq+KnuPZOkZYi6zd36EKMqs6N+u9q3YkcfjlWU9Sadak5/92CWL38
xtjw5ypaeIz69q+yOy3zXFvy0CJWLurlVyJ0L5BT4qBX6JOgx7NrcLMYf15iAWt5KLQ7JMJuS2uv
NAUP+dhss7n/8B5sZkqr0T6c6aoTmhKDPwLOpL9fyeI6szlD9r6AYSm+xO4tM2dSeC19XnfQo9wH
DedaLpuh+7OC7SD1lO9iW2NzvJsSN2tuUgO3ocEtb2ep5e8/XQPYxv/7mfTWsF/HWOJhBFxbK1+9
U2sBYZRJimPJb+DfMbzVt0i+TOfGlDY/w7R6pmPcB/RCIRqp6wWwcpt1H9+XYLApxDHB7Uv/JIJi
4jumB0OVRZtd/queJdCr+pgI57zjNrr2wVyPKTiyq6jl8muhA3BaA/kE8y2ZpHvtH9CPfWZlItOI
CgasJHkMgl7VZU8R7rXccCU6qcTJtYy3rbtVXFuOgaAONKH+2LCmz71gVSUkIbgUwS/PZAtgBI1e
xXM1xf2Ty8eTs6rXdVJEhNnppSPLKnacUHxXwtoJlXmp6wmtZDS8dik0U2Duq3XnFT4PjnB1f36Z
NMVwTc3wPO/lAj9WFcqZG6u1+bCDpfXmB21Hkrz7szpfTdt+U7UFtkPqL8g1c5ubFzrmm4q9eE+n
Y1M2/Kl8jiEsPjatRnFWgKOF0s9VM+aINxZgDsJprN1l3thZkiah7izWYfhZmNr1NyUlu5pgZtq8
eqmN0x7Us05AEX2Kgz5CBQEF6Z0lo68rU3MAYierYTXX+vorM5AgBXZgyO0st/6wfBN2diM11BaP
hEM+7Gz92MtJPW4m0kWG+hXPdQlI7E8/sTQxMhZMx4fpykBotmN4xbD03sb2u5+6XvhiEZgqSTy/
vmJ3pfFxp6kGVQ4LWj7+jKLpT+te17k92dLZBLfuNGP3p5DLCsbw5BZMzoo1c1kJgjl7EwBmrnN9
QFItEfS+cfueDBHqJL05X2oeVl4mguvd35+KRVrLCpe9xUw2fQJdtNydFKR5AIUzECVslt/jTy6R
YgbbYfYdK3AheDg/IKcquglKkW1a+D+GNotcCdhHCqgmlgi4sVfbxLoGiXI/6Gshq4xmZcWUceWY
7PPNa1YbOxxu9yKKD8cVpaKyE+G8JbkJNd9sxQbL/gBClkoMJpqOYCO19N7iI6mmUuNiOX+p02Ew
MZ8nFesIViSGHEjWjJ18hFcYF6AlzXIpo/3M2ZzPT4zX2sQSW5LGcP1JsGUmeJawKYDFazN38CxN
mhd2CDZb76UwDwTlw4BtoGdTmi/fjuVsKfYeh9b+ww0gQXAZDSMt85gZoTzpK0HNFXADaGxob26g
shvrN2yDUeGbqZsvvOKe1R1xT90W8SJ7Hp+tpDE+wMQwEIDnlovHWBI7w1XMOiGLWSMJlCEzrV8Y
63L5qEbXlEZHxQdtJZDlptTtAAu3PTrBDfmqyCk8M2K9wjinmlVzaysg3tb8TkuFMkrpIYH4zX6j
97B6qw0Gq+Zeaoqy6SW1kvzHj9D7in6V/WgU+so2dEkrhsfRS294bCOfQIvRzfIXFCCpoelJHUpp
2y/AzCUgV4D5yvDIxdRwqXIdvUjQbPUnsF29iyvxsRgWLkeNHJ553L9lmGDUK2wYkgWpRgsLaEJZ
FKLbmmEJ65ANnfGyKybSMU0czsWBPT6PQLQrivFlNkN7illyctH0BXWrOnF5L7i0RpZc0/xhOvvH
TXz2b7XQgkp5BCUUXT0KMY8B0cQR8Y3gJ/98wpuwM7wWz85qxLUlqpdfXRa6476m9G7J5whTXT9p
89kHBp90n3Ch4L8o+H94YqqPUD+wkCWLhtGfKnUA63xBuiv4R60QGZt+c1SkUoYn9RxwDDoNc2Fe
d+RdyOeT+J+NVrAVAk8cibnLgmevRV+GFgxBUg/63nDq50IlGPyqOFalwwGP63Cd3LcjblK9vsQk
aPLnt+ZDIDP/dNQpB7ng5hgY2lsqAGR/viC2AML7Hzls06fWFKDHa/W2W2Sw87k7OOuikqsae/1f
0/0LHnFQ8BK6KPTECg62x/lLbgCV+AfNYVI0Qkc1ULW9URSI18W/jN0M646zk8ORNXnqocVbWTUU
3Oe/tZ7uA+Ck0FMWFtfgMaJLl0fqUabmra2bybaAPfXevkn9quDFytyPcsRWVYO001v4X1oNsMnS
sOyZf6nGCQBk9Dvm1GMrptvAeS1NWkn5392Npm+la6IrVS7uFzDkldIr5v0IItQbCLQR1Ufl19ex
0l2WRCDqOv7Vb8FVzOmhE63EvW7EV2MBy8ymV6yMFcfNwKse0kI6r9qBkBhh2KjIGjo36vv8mumF
yishDodvs+sAH5immwtc3S0+5lpdu4x5U4xpN/hAmHmZaG9AkH1A+lPPdYdd+PaoEJh+HYpJHuRS
NpcFHMonxNgVN7kkR0kSEtTIFwV46fDsiCTECpT9+HCfBP1kNnR3NnpEGjLuKmNaP4N3cZOgaeIG
a10QIv1ADwg/ZjKYSJbvEnNiqxGcw8QTgXaaDZ7PlzNcAPIJkWXLO5s6A2D1+/FKMTyT560YSJEr
SuBuS3X4Ru6OtdsgQhRoSITgPf5nEwbSzVkHOpsVDoRl7284Vpgq9aohBsL0VXnSz94ClxK+nazV
sPlscON7E5wNgwlcKv9vt5AID7ClXcm3pAj9OK4TEGQoR3kGVFhAx6EHlTRicK+cyvIzDdy1U30E
pPUBK0gNNIUNX3uFBScmQ/NUfymFZuW/mSD5fOzV127VuaB8IgFoWa/GAbrWLn6kShOhqF8mROnx
I+w3mNzHhnJ69dVjaY1LyoxHrnNXoh3YQgXasG1cF51Y4o9ktZhlAhy98cjjTj8rz18LnE9x5ScZ
vM3CMY2pXtCL/YB1jdwifOVOo6/URCMkXBI+09hJrEu4SE+M3BADZhskNHOJYFdpp29hpQZOaFZT
Khbuz88pbKl2j/U8MhJzGtz/1URHOzyK3PHc9LdWy2ACL8TieQpnz9jOIqmQZhLxjO+nBOpxKS55
TJqWuhLzffIvD3R+5lXSAjMkYm3jrC0zhOI9bXKhyDLx40WayPQqYCF/5T43xtdJPRDM8bp1/+vN
AHqvZO9UypcV3t2DkNacDC4EIWAIsDdN1sHS+q/xPRs8/x3Dd9oMqrX061ECCgGPtsO0W1jGVGih
FCyEFP/r7pejtKyGfAQ6TS66mmzbKRWIrs+LYaoEp6wlFOp0Sy8mvhq1zA6WpfmQKFE7PPjZ/YUC
H6BK8sVseRl3tZ1l16OjsXNgHDM9fgqfbH/81KPeKvKQXeG5otrHSR6Jz9scK9vXuaICr55Gzr5f
nJQvs/ZAVO5n9vRRxzlMPrXy3RpDjmww/gBcXs2CJmSem5K9iH0ydMGX0FwUOsYNLzWNOO2AUspW
cdCq+VUsBC1IOf6ZM3UutikZCTDRezI1MBb+hpwa1y0kVPBDzCKoEiv++NuUIRMQ9D40JBWYri6V
fRRwCoM7bVxSq63l9PVLyC0qFUnBsVSxKF353bSPPUHC4WbskE37HHGiiRYJxSPThUV/krA/lvSo
NbpnNJkPrS+1caDO+UmNPbMWdhv1UeU72k/Xhj5tL1FZi3MFvhGDjHYSB5oP92+R8Q+5kq1jpqDq
xtZCmvqxGPTiC6aKNRLfGMkRP8rdpmKm1PFIv1t/v+jVsSqVkhjbrqQSu9iSS5jyOz3TBv5wtRXu
DftD/leVlFzHM8SX615Il6QJ8tmKUCxmY8rQQhwWQZAL4TewzYUk/09l7LeYqT5TO2yzRJRO/0A1
TY7SC8dztuu31VNbQ5rJBcCcAvlIxGfj8deoZ17OE0vWD0MVJ+FVr1pOULsXz+oNJlA9ZoWWdR1O
+SHPVHjioYGJDbBdNY4a5NuS/duCa/67UxB3Ex1yOjS5JuhwcoVqJWwVzKXPE5tASCwAxPLp880O
PsnCvYcMnT/0DE0lc0cdswmzFkTqPr2JvjUT/Uk2m5OrcmlwQD8l6/cWCJeKmUNneu/PLPgqB7Ih
TiAvnf1hCn1YDnudn6df3VYF0eJWydNGsD/tj+yRxyyVB2arGXstO8+NNAwewZOyY2hMmvSW/5Oh
GNu09amZl33LsOoZgWs0E2b/iEDXLQkRtcXfWK3YLq5vNf3/tjWNeGtmpy+xqHmZIVs0dzvXdp9h
yLoEoTFqkvQUlhlVzaZzdx/FWbHQsyHGhRPSELvPATbIKGKc7HFKxacmOnGytW3QcLjB8+MAXK9H
qLKdMjQPpc6pgdIL1OTwO2YWrtD7sHADIlpZo104rGJm+JN7bHypiYqQJSQFKs2AjPFrrVk+aN7y
xm+js5AZxunMf704S5J3kZv0A0Rt9PWgJYEmZeH3q3zH2ZFGRRg6o2OSBFQWLfI4agSNWgOCWz9C
zbqtV7Wx/vjEvqGFfbqpHkwpAnSohkmEgAb5oiTknuUhDb50Wgb9w8N5VXVS+S/glTsw5kcU5H42
Ihmhz9kKemzlRMkTTzWp/X14jnpBhJ4UvbXvJ+vlatBi9KUkO/hwNwOZmeElYVfiXkjuho802BIn
DFDgdtqzWkuuU6NDdjlwjiMZFff/vzhzjQQQGxSU9AQObP4A9lKLqE/Y9t+CwOVVT/gRPQHLXNuu
ZoHEbID9i5A5zEJC2mpyTPMQYmc0jCUOi8HdbmvnrGKoL3R+G6DduJBs8Py8P44j+WXWJbJbwlN2
uoU0OHxgLLHWdGOmLrbLknDQ7GDhNThyqBx/ez82i/kWg/ofLmpFDDUYlaBlV7E6MflUp6aNXcPJ
8wsGaDEgEnN1vYGZnjpDN3S/JZ237EsMVNDBLvSGKQ/g/FkP6RpBAZI3rWGi7uXQG1imCI/BVSrQ
bz0Xg9CklSP9zDxhcQN4k0z8II+cZs1iEhar1DwTYgb9jA0oKsvC9yLBovOuoaXocc448asBIg/i
niuxJg34ptG7Il5uIvX8A4rIUr7o+5Tsy/SuTReoGZ13Rr5f3Q8VfqcWCxDVdpJpj1OKaX+xatmS
nLYcMhCWBE/KxzLpdfbEBohtYJqAaFupY1Zgv6kpg0a+DCf9b4N/A/H4tFSxry4MoyLyGPzFN+39
A3sQxk2Atxd9ysLFcFRhSLdYewP1ElX8yV7va8sBQddA2d6qBSzs1yOFWyAZXtF2dAxrP+kdl3e5
WLlXpHQe938FANpf7p12PuiRbeMe9UOmCwc3Iy77TPOJCPbC0MNfI+nCCjN1ErRCuxbfhyEAG4Wq
/T7czsjxLaPbyE3jLj8yOqcAp4m9MQfN6fE94LOQWHQ4Aklf36YMW8TDd+5vACNHNloUyVmx7Kdq
FBhmqR8s0UjgFWN2KKEf7a7iMapgRFXNq4xES+R8wTiQSqKeKE2YRJ2vv1AbiEbgMaOCOghQbKIM
rF69laaszqV1yJ67Ud3dixeOS8UBdv9aTLotfVvMwNAghwP/D/Uuweavpa21faNh2Txj8lhPIvU4
xHhi00ORZTDz7NHUQiNaa4Z27pRm9WqhA7QshBS76b04I5FvMTNgmFdGyLSDdY19TSr+iUxb8/ps
UY1AGAL32qgAAMT4KCdj2GJFWT9hYTuCzPi/ILTvyCYe3mPZ2gW/ioC1LNzI+mJZR7i7moJ1/CH4
wlvX3Yc/mGhr298isFMV7ak6pn7z5EW8kQxYRov/HksAH+XtLESCYz3zKZRz6agxHTo10UdgmFc9
p3J4AjTFhbYTYIX/KxeYKTTSmQ8hGB2IxDH+53ZA9RYwfDJOHRA0EJfkI2TCR9vmPrNHnbFhRR1c
0fvx+naVZpQzCk1ids5BGyRaoMJGhlD4oHZ//dgL847gZMe5peDjhcxhvtoBPTl2LbhvNAgepogB
8s9AmUQg+VMa0mcQX3QcosLgG/btmZECgTRvjF6FadzJhP+p24QweAB5eqiry+J+o1lkbFriaRvQ
9p+Rht9q2WE5WZBVjgxNznipBSdY/KcKbRIrOGdikkhwWXhTInvyKXdXnh9lnKfWoxTsTt8snlKo
BvzjfLG2MMvmtE/ccegPK+pIQHqk3xSJ0sZEpFaXN22gL9W0/YGFYryYxc8WzTfMSgqNr8KscKPv
RMpzRsRxzWIf9vnmQiQQtxaqfXKN+ohqL6kMVZOTeQateShwvSoOnXC4VuCGbQ63ldvZKdALiFgI
WIKRrXA8HwhnEBECHtGfUQsXgm84GC1iwcU+1MWhoj9KLqP6D+KqYRWXmGIq6XQ+tWD9JomfMcC9
5efbzx2lPvmRvCywkg6iFH5s8BtdHvseky/9/+++7mPbTpIc1n5S3x+LIpNNPZqryk8FaUvKm88E
qRksH4hoo/Bhf2ufH7eERSO04fotSwwEAWjm3+SKG0Dr/SHCcAwR78zoaPhf1Ge4sLSk/09Fdu4t
7o7g8Tzmjdl3XsBZe28cmTeLZ+KjIfDWoG/h5GAeKrPSEx0WBflYFzBr7WgQ62b2Z2M0YChQbkda
ek0qAs4muVRLASy7ByaTp9eajKAFKdsqgHJGjKCsab2xTGtF/dDv2O16l+rRbtBG05F4wzyHYd5d
orD/rDvDv8/XalliAabDtRB3WIkbz7UCzvF3At4iKHPFb4A6CGsRpXHs/rQpgym0UWiowycyKeG3
T2q927YtUMnXTghQHv2qH7t4eVZWh3sgHZBKAmx49e8nB7YqMjZgU7HM3EAp3Shn8W/XPYBHK6C4
j//Gwg7wAMuRQzJ7V9KcetGC8rwlx7QjigHRDc1XhR4EWxaB34beKf5B/UvUwB1fP4eQeLEIEXiF
9i1D3lzd+K6ez5AqFmFc5VvKTmalWtj6OYzrt8tA8Zch+Agtj8SIy6Tknx8BtUdZBa98+mdk7fDL
oJyHZjojtZ+HW5hkV3QYXu25jZviyoHhzemBJcb3ode9FQBhjqozPZ6LTZIiI1WUFeoRlYvcb1K7
EavDs7qzr5afDt9UQNcRptq0UdU80dfWLtc2LBReFwQpS8ogNeDaEG1Ihg3opiEvfPN3WkacdDxF
qzfZjxKf2kO6xt9cKAAf/SCCUqpQG1lHmZJ+i9MIQYmjw/Q9Q3OtXFUsUYCW5Re5vxKto7NydFi5
DwHrWWubTSa1YSTezXj8ICWbxLx7tW5l6y7rGijalMzQ/2F1nwV2gu5rM8tcogLu/J0fNf5+3LbF
YnN+CLjEHtualTYd2Ty37RpJll/rUXwu97TuapAckYuOjBcvF39n/1uBPIqH4NvyT0jXCFrlvqUk
MxTg12mA8znkllh6ve9TMjnWGZGVO7rID8nxQ/p9LU/Kr9io9VODoqpaFtrmVyClObhRro6hDmkH
J/Ocx3PeWis3cdFzfo+phgsbRhmZjUGP3X6vG1KQfEA6p5gCTo9L1ARK1aIVSfVedYi1FO5fcSuE
ZoVXwvBYWCoSIWQZC+bcp5gWxUgmenMiHiKo//gb/IUAYj1NyTxjKcQ3B4MXUodWldwYkKF42uPO
/afrSTh5zoPIac8UzUCpzqyfXIZCBQQ5zWWw72pOCVubW6Sfu8ru5ko5E0nfiVFn1jFB+fy3HPTl
qBl3nE6Db2jMa8aI7MRXXnzIfk8WG9wfytTd3RKhxihCZv+dDycwQ5JmXY269fGXOyVm9Mm8YuX9
PG4S20KGSnMYn0hSs+TB3LLWPdmga8DBFjma+mJPSPalooyGpLDoPPOzUsJ5rJJgeScN8lMSzhuI
uZqMxw10Qaw1pWOZEf9Vx7IdolLumuSmuz6ZXWzuFOtKQ3B9VZeM9nM9AUYDbCCUycsBz4OKktqH
rt7UM7urnyRYqiVaSOfoPDh/vX26K2Ng7MnfzimS7AOb/l+C5hrorPReeAalaEEvO9f8F9OJqFRw
QprByPvmLvm9F/2y9a0+jY5E2qCh2WY4hHOcNFm+HW2ZvAWPIQ+Sl6DGiyrEmLl37ZzRtbUjN1WN
MRw1PIzzLndljsbAmbBz3TyVnRGB7394C+hr5FAp409gr5Wq4rhK8yfsEigz49jTfdMhMLVWNiFj
VsDjR6kOw1hmuQY2WtHzCG080KGR48oICxygQiLbR8GQCRExH7/orQJjbu+wA6TJVmBH7klaBO76
hFREXLeKsvVWIUxMrJ/C4tqPq0poMRm8UW6Qrp7Iz8XbJhU+QhuIh5uBKkGAxy5OoAWSPacpgILx
fMiKuEtTY+EsNImfEc6cU8itCaxtkVZsn74M1qvhNQ1XQJg+absNM4asVr86IijSkSfd+emMOszV
Rrqi6pMgFiOkliZLL46wheqQ2RA0h9K8m8YNvpM0RCCbg7X5YXT66QaOPmx3Ix1yRWlWYOwG857J
gPCEZnHA8IdGBvfcs5kBf65eEPzAqlVwD8paJ6Jmi/QXaVqMPmNFhaOxnMBk1VJnEedpxMwqBkxd
WVxdq9ARtJB08SU7g4hzFUYcNwVm+NoVrxUtdEH2vCODkXa0RvFuePrlpNKUrxuNgSqmDZ+uamh7
nzzqEZ7nr5D2QAPUQaMjt1WeztOkI5ICtnoyxbkAGUyqANucAWd38IutGnEWMoqCOe8inSyBCLK5
ZyFGw6oDdO3CkW13ohBlgfcaIyYhTEqV6xNQF0pP6SR+xp/Ekpw9G81XbSNbTebXBapYXWwgrSlg
vfZIGvr1cauzJozZv/eMIPgoFKo5Va/KtRJZt/py0jQvHiPpW2za19xcU3nunMMBJq6qf2oCoiNH
jovMORjBG51bOKgExJEZSf4ivcUhvcr7f7pZHLJ7uTY/XAs92ncZ3v5rY+v/QkdIUdrkz1KkNpbP
uAeEWrLscsRD0S9AMuGixNRXJl/HcLvtCtd0pRy0usuaP6CZ3udqR/5Sx7KcJGNvVxLpzyDUPrw4
4qReOEuapO0G1b9UBgaiiN2PJ55TNPyY1BqSVpLE5/C7TTgKZY19Fl3yvtAWkd8AXdj0uX4Uvh0Z
kfAxFUzbnY+4inMSN4VQtlDR4xFlNjH73ZIth5wZ3/M9dYyWtzI8eH4x91oaJZWVSbYx7ECewSEX
mwxWcbMh/KaS8mwlG7U/bU8Dv7F/T5PvgrSWKLpzr7RSs+NeLOIs4fME6JesUeMeB+7lqjhi7niK
FscMYAntKO3GF1hn8aLJkAz/ygEBy6LiWFfcd4iuGEWL1IGjYn+QgheOJHDGWKtmI08bG7dO7jSm
S4xzRRTkLVwsvbC17BMPnulCGZ6TfG8gbIa7xBFWGOrIyJCQXvI15ePfHpv/R8hh9Eo7PMNqm1pX
AjpOSZPfszufqInrdGaajxPz+pYUWTJtsCxq7+6tvSrsD+XCsoo/hGKRJzNyBhMfMuHyAz61xQqq
a9Tl3FbZegmx1i1ZPnptIz0Bygdo4uVU8IkNV8uA1LJA7uamW3h77tqCyym6lj4o02b0ehkZtl/o
MuejgiquISrK84Nyw6Y9P+778eRU++kMauoen3YNLIoyBQdyQYd2Lne7Bbu0UF7h9XwOyXm2hcGW
Pj7SxZq7jZwkuFULlrifpQrJzvaIFYzVgJQaJ4pweHiZOgA6Bh/Aj3X9akoZeoWWLKEItskBbOdR
AM17xeIokEV54TW4P3shhzTuNWQPcPfNrfTQX70K5Ot+1jShOE0wlWw9DP2iPT94xiqCUewn19Uj
b4kvzpiiYmTkD256DpJtUdEXNrUIq28CJsnLgdRNxEjvrR4Ug6kYgP9OqinbMSQ6GBdqQ9k/H4Wf
6yuzMx3H6ie+uflWlmJUBxg07KK/e4RSl0DLvY3sZit/0ciG9vJci0v42jPetF8qu4nQdKxeYh8q
3q4gQu/MX+4x4HvFScuJ6FGaBxrA/Muo1C+Y/0pqRtqw/50PsmYJ741jmerqP2qcQ80zyrkehcNO
PgH46UGOYS4+Nj9X0vLf4TXfXrbB//tzaCwKxDd+gTnouQxVnggUpxq8Y68/nvAZBLbRqFdzlEb0
SDN2BxENBcp21FlMGiG3W41t7rF+5ZuSvWg9itMIk5/3/Iw5mZBtPqGpzDe9+Vb30340Gz33b/Mf
2Npsll1/6GA0nzVBgT84M1eiRyj8laVQ3OQUN48rrKuGZ78YdcylphcQ8nhRvP2BCGPBY8AEtQTy
lpeSSXqlsxahA46YaP6OUR03bqp6IHtvzvsR+HfuvcFRfIOHj2SPE0dluv3O4bRh33uRZSm0Qdof
Vk78CCswGdqcDLXvvL3fOxHkIPIKPG6reNXEmWI/OoS3yfXqJGH8kFP1GbwX6Kt7vyyET01Cngzz
Z5f/WPqargjhRoBKSI1VuhuM+AKC3C6npN+jG+Z3M9FCG2LurHFAeIuBJHhTLB3sIecohDj7ddic
zf+7mchhmoazVRZnD9gEZ4JZ8NPGO60Zyy00Cip0UtJcAGfV1iqjCkL97cnLsZ/OZ1gs/S7qhV4l
u2PL86LL/yad0YlvJmo48F2g9cdxvnedLJRmVYecdW8QYFMrBLmvudHqoWtU2zd1Km8nnVOm4miA
RCnq2QBHkjT8q7gn4Y4+HxBQmWcsWWyrfjxCKoNcTi6LNwRbBzkpikJShWMHEpObYtGlDcIV7tlp
9KEyy1UbUzRvuvfdV4QuPW4fbckYH/3Uyw/w0wCkymCjtt8aOQeqt//bkk0GPdHm84zux+9uyLx8
wUjhL13LOWGWNS7R17aGG3dxqmFmp3AJmguCf+srGdj9iYe/1oG2dikHLFGlrURKNxUB2il3GcLo
JqD3A9sSws+ZwyKwlSrCmrnt00djjhWy8Ett6q3PmBMSAJ5hRGfD6QOz9BQtR6OVUZXAimdyJOVn
CX70H2v61s2ScUU8UxLfVrV3T7M4BZdnW7R6V7hCsuTr8XaRj3NWklyk2YE1QO5uLTbIRJ2XK6Qs
UbzIPYiGaGMYakch4D2zra2RVBJswZk3jCFf4F6u+r74h3jjk8cKS6XQ1VdkmEo/jFExADkg4wqk
NYYvzPm/8FPRdvQ8WavVyWX6QozTdNsYyOfWDotNPAV3MSSd6zTxE4xqhz60c1hfVudKFnziqTXE
Cw/etmvzxkFJMStzrrg2P0DdJrydMowQLPDyp6w+8e6LS1mbphHz2I2Lr/lukobm1z9mpyIHqfZ8
BQhTO//LIXAPlc/dzXTsXrslrrl680w4c5auqBh6dvtWoMF5i2S/k+ihDjOL5lqAnM57+IG29tN5
VyV8etz7uAgTcWRl8xptr7S+zNTi9CdGoWmGh/t9ZHjX3WUj9kTTc/UG6Huff07uBN2hmraAOwTX
/OmVLCKoLyXkUBCnAsj6lzCE2tkmb4pVWs58GJnTuuKl3gF7cU+kM5xsUfUwo19efv/or5ot6rYE
0M2xagsA9YWsuVN/+1J55nf54ILeoHdGOF+fntvm0zLZh4XDhw5S5RUOA6WjXRnVUE8ov2gBEy65
hrJjbdtjuVoyGzvuKsUgiQ6kvRAbzio6wryxMRlHiSOhUcOcizQ63alABPLbNK+Aslo/ZuNEewlc
eHDPBt3LEBgCBLnM42C4oKETWTmmQ1bV/wyJGieIgkSee63uXXSvl0HDkJvX40Zm6Xod0x78f6FH
q9ekRhTigfOS5vR4Laz5L0OmfH7svdq1FMMf8RcypTfsJ3t/knOlEwkgbikt8Wbu5ZPJcEXU2LRQ
BC56TQ3ESKJtEbg2xKiVwY8C6OlkgW7SNiWTsXpIyA3CmD6YmQ8xFHze/kKNVIICW53AZm66kQFT
sswmDVDj+5RczYYsS4zoQqBUFnrSVTrBzagUzdGR47soEUA4vovseA6ka3vbFbuI//+x9YG0e2od
jaLqEpqbXr93xX0NAsPCivJUgYDsXPpriWhMwxTPT5wQClxAOCUBJjrO7tXn3NNt3PvX6H6ht0aX
V87ucDl/olhPjDb0h4rHFwurlwIuMinvKZie1f3ebYoTevxOL9IGu/1k9mYglqUnaUIhROGuSq3s
PjCkL9C/WKgunNF0tm8xiMVQUs5wRrNQHRz8EXrUJtp5PuD7aHFnWav4vXu7JMtSY/N9wSyAg6se
EIcDSEoPJrkxCtY5x6Yh7qEg5fnrACNIoyFluvscygbg5+U9d+rAKR+HjW5xnkEbi5q3qyO/6CGL
q5bgzF9U0b9tZO32iZJfxcMC9loYXczb/ok80nq8ffQZxMKSG001s7NiBlDbJ2TpP8lFmmRsVTUg
XFpWEEVB2mgh6aLa9K0VfKBfu8y8Nul7QokKiHTo2ipfEbXmFvVZgbRDQ9ps3fnL/mMrL1yQ3ZJA
K7ANBCYKVWAcmEUroMWtLK+FxIxrmWUawiazlv7wnBU5rzFLnxbL7XB/SnbAPadwGwaXuWZloLYZ
4W7UK3Wd6VboVOc0MK1/hPGFEV+MHNKiqsakGsksSIW7ZqakNW7M59jWKL+t0qbbK4pMAN3RBEy0
4BQN4JipqUhYlZwDR9GkRlJMuUDEhPW61ITIU2CVZnY3Bgl0B+QKRlkYHU4sBWYjU9mKeG/BfWVD
APcgnDMtI5LjzULX4h0wby2lYwjl046uF+u0ZijmzxrDOtwBkDAhZTstRTAy4bCjz9CeN5k2cuTq
KT1VkLoF2kd/P4HKFBsS29lTuwlnP9XliT2QLH4mRk/ad5aDZInPrHrBZygNzmGMMbfKKNRx1VuA
qeyRS/MCVJ3/4KxpXiTLRmzUpmOEdH/jMh+zf37A1hmB2jgvlKuWNB2Rt/eiXnFMdrd7MH8flbVD
DtyhDXzIUS3z5UD7IxEsUEBIc5nJXcY+o4Td/s2P+KS3kkG/F3qilinZTYH+oKMGZus/hshHyZ9V
Ek9diNjuqD8KCn3V1Z5o/aLwFHGon42LxeCk0CTlTJBBR/xt8wwr+ndmejSofWT0JEUqr6Sy/9q0
IOUGEZOCVrbsZyU0ye9oh/8+EyRi3bSicwMHOnGo0Kjs0e3knk9wbkgBZmBXLGzhxg/dIBr/BwIo
5Ilipu3CogKT28+0ZL2hhzDcFSZzbR8l8AcbfqJoCYPvvZG/CBmLtfSPiBjEJmAyKQi2vgwzKRK4
h8Zk7e2pfYnB6fujms6zZBTFmemIWlWCUxjH/FN9SVZK9fY8s4DCRhMtnCLL3lBSskLusrtqfdKS
j+jKa39RNDfHlJE4Xs1G9Z5DujPyPWK/sSIW+BnFjzjuD0l6KrqxFBrwHYUVnxs8iNADf8ee6H1O
RioA5cvEQkiAF4/XlQidL1eAy2caas7IMRHFzsW0g5715iLnqWkhf8xOJhTbDTzM+XOC9+fhJbbi
+ZKiYCoApSC011Ru11TZ7UxSohJaY/AuwWhIo6XYJrT5mVi/JiJG3/vU8kHA7ixLZlpzZ5EcwiuF
A1owcXbLPhE0oLq+LOepEOdvwtT8o9OcyWU5m/n/VQrsXQbASES5S5bWvyq4X3YpC4CGWchyK6j0
MKgb2qRwN/x/FGAwSQofXI+cAssNtW5JjICbraxeGe1AM+Dt3qyXeybMFuoY7yPDQd8p0F0efdCF
xCxhQCI5d0z/s+721+O6DTiEkYGX/miZnpfDq/YkqXeOjO9a1yaiJIiL1nWdch7HJEHshv7qTD5K
bX4uG/moPl7Mix+AsJjiO971VVLuLFzx4EIdJ1RUJl9zwy+oEAEtHHay9SzwFsMNyuAO/FOpZpru
Rsk2Bh1Y0TbjEG9ioftQJj6eJ+cWqVUTOnu2HNrWDLBP7yzMns9PsPryemlrg15ZTm1rugSyucFb
tkL3ZwQJRyU8aMtW9SnGcK5QFuAWRSJN11/7NwnIs+Ud3u25vIizUuoQxYBGjjI6KVa57NiEFJYF
YZvmA9tJgKzIVSGpKxevWtv1AYbPPGPN5FZGySZlBynN3uUkBFVPvgIgrgK/ulKsPtAVhrCZnSrZ
Erpg3He4nD8tPDYp3seblEkiLJNTh9NDHF9NtqutE/z+jZuWqKr4BdBu1tBF0AxHc3ZeKhEeITSN
jP2LNyqJcIsdeqWwtARKs4sHrXWjdJoirj9/3CmVJOx327ayj18A2E0uKP/fYFMJ5M0p4CcoTumD
B1V7lTLeVetZ79sXq1u1A85APt6xXIjPVYnNCZp0JG+CSr30Fui82hdN6JHVZCXKQpQGblEjmC0o
3MI6tc86u3kelAFf+J/HxAAS/DmEj2YR44AOqyHCc87qoYE/6eHbCObi4qfG3hBMi8gpFjOQNoDs
PW4ytwkfth7mW9i6NZIl+sbFq2PNcJzvmJ+GhcOdMnVHkv8UdDc8xkQeDR2BElRltG643HXlPVxk
41HbwZ6Ixk8B97687gPadLzOBbcgW4urfoc6KvrxLx7Rj+hVD71DQCovYPuXkYSboXPOIa8tKoFm
QY94cT0qCA24G2wtoE54FgN0+u6pu9liQxYfjzgKADMCczbB+10h/1XdW0bDE4cY6+7OWEu9d8jd
Z3UG6fWfij+XzW/7qDHF/KAmex0KKedzx+lopnTQrjXGv/RH2Qr75DAw5fGiF8UDqixhL8qlBZPg
KBnFoYpXZo6lhyRNukVqb6XR1lPy+yGjzns5VklIQgSpd1Z3zo8NCLFXXMWKzm+Q6l4XN1pWTx0q
jDI6r3+eOl+PbCdECeSeRKl9dAs/04xX7m04Wb0vDraIJRpJWoXSO6HEEW+ohn5HArWhKvYzkGmk
w/UWL7sa0T1tt2fRgC6nnFt3OgW6lC9aXtn5/WNl1s78TfGxOW4KA7sSFXfJkLdLsMOuChQUz3vZ
DrCOB4z/buqlSuNAup51WBDYNaAcKPAXK/PytbDuX1y5TGUH37vH7komB6tHKpJO7N72Z7LK5Rbp
MGtwFhuufoncbrniUmjKcVm2GWlMsllsQn/88R1ObzIWxdBeggD6KkRMWKXpPyXKebJ/xrQ3ZZcr
PVsskXtZBPnOFwwcfN96/kMCLKUr63Z0g3c8AdMStxeQvzid7gfMqxpRC1HYIvFu9y1v4Awmyozk
7Wr/ODlTrfJgLqL3lAI08FF590ZvdVgYmLmOcZT5Q0usqhM58FwDTIVArA/nSd2BpTFFr2BCTBiZ
yRTowd6Btw69VQDYtzD53PYzKdR2WyCcueqSkgRRs8jVlVDWJaRmNTqzcte+zZGPkx6sENi/YCFQ
wkeQw0R7ybqMsRNpZ80HeITSzfUUY/cPxV31K7DEzx+qUt1TPitiVqRRlr2hW9eNIKbcvQTCE90X
ngTqS0s/9q1i3Lb61msr7NVtOTqgs9r4bMJbjpX38bB3bx2JWdD9lp7tqrCkuX2LLZVG501S2yiG
fwB5iK5XMdYfgxBWcAGllregpdvX0kmad4V0N4SZwbS7qkTitsuwh7PXM4+XTLtks3ugA/71s230
oucy5x/MMU155MnIOJ6/v5TF0OwaeQ5Z6Jx1fCtmBtZ9F6u+b8RERQ0qcryhkazQhcbsZZoas3PT
yx2+WSj/FeEX3cIraSXbVCTE9VI6fV+pW7PhCDC+5S/zJwUMXsEuECqoq98GimrZctlPnp/lycuy
8PKjVQXC5UsqQlD3s5bK/O0n7i5obzgVG/au7aSvsIUdZ+/gtjlZU4ibIsxIwKNZDluyI+5DKuP4
4H4jcNO84LrwfpEFXCp4UTNdcqmzNQuZ1EnfKaT3dF/wcSiqDjQFrZxfA/VI88wnWRRT4iS/5wMO
XszXRqqUFRvx9whpeHpr23iwpS8vHNkCvn5JpEph9u9WOjCcyfNL3w2P1GIO3w+IjveDG+m1DaUL
ZIixnhoaS74ikkNshUnJnDcFS4YU+fKb4K0xQjwQgMAoneWbWfZ9Ga80wVXd0biC06nt6JmkrwTB
DMLcdQD/r9lpCBn9VynoH1mRbzUgWkNAXNuOzVyt1Wp44m0CAv1LdK1doRIQESXtScaq2E6AoCCU
XnJVavPqy+0gxuRW45sGn4pIr8Vnj8EgTmC133JIEiAfs9p/8RZofRAm5oxXAqQzDyALX8p7b/IG
UdGplbgPMArbtaMJItHJZpoTQsi0LG///pMh2HeLC2PkJbQG4cNPHnPmq04R+EUNgiHGl4EwK6Mc
DVhMpQUJ2pKUTR5b7Hy5OYyRPIo4z6+sSL0oS1CEQSicKv0dp1XA1Osu1t94+zZvWyQveleW+L9F
IOVnIdgiP6ky+0tYudolHxo7sgOOrSpyOXsJ0O1ufzfc/gxEDYiDN55f12P3zImzeSaA4MomnMl/
C1tlX7EK731v4f6Rt6npFUUKlYGkByD0bcb8tU5NuxJASn6atbiLa5HWYm+EQj1ygTVWIRRkpaOx
SXiLWjEsv3rKaPf+oV2xkyP+Yks20qgqnhpPTSRB+Ugo9ag0sZKVCEQ19Fs7CeSpQr47AbMyD7Dl
JbAGeYFzpXT8LH9e+CGP1MIhiVGY/x7ntR0egjyWVLKmpvzZgp17K8ZV9jC5sGVpeyjlwxmsz2Tm
v82/u914E31khI3IhoiaTbnFqYhTbp4hE4oiBNEOtRGxoKWpE9tl9pCfcIZUs44uKsbEdeROvy7y
eaGjeh/KjksvZsMxWT1hL454GW2l2Vueu6AXtJXTBTuoD7FLrM7YkQY6fasuQOCOhLqt7WtObapB
ii6hKoht8AncLeaukD6l12d+uf2fMY1j4ocjqF6cYOrC2JFRFUkbIQpSiVjvriYSnbaA8yMUiyWX
b/lKGrxEWIW2cMdmpJpbuOsuMxcMCcrVo7qQU1s0aQ5sAoY426pA/xN/sqw7lDCs0EKI+chf6C2l
2de2zpuZSS40HfB5I7aBuTDStVQegOhwrGqvQpksd4IcPA/jLngwWiRy6FYA3ESCwHBQIVTWU4FV
86qBuGtmAEnn5FHyOD1qgmHG0dGvUCXVu9n7sCQiVGkeTpOWv1Fz9WqoDvoyDNgg+SgLN2p0SrAl
9XdF4KhWmK63Osov1Vf3M834zO37/YYdE28wk4DWII7rot5TLnmjycSIjP1wNes9mZRdVsxkPYi0
LQhcaPgrB68R5yoPRHMEy3QrsaAS16Y+sG1NVmm4yoJOr1J/fprIkD6v4fDQJTB1XC7UbUZvAGpp
10OlOvzGIQvjWBvwO3o6XcIylBNjAElMGOAB+sBgk2aIozYuUx0iZJEJjFYNvjcWGQWHdBUCzH/a
q3hL9cC6JXLIT4kz+F8YLTEWtAirp2gy7FZwO7L4U3FwVUOH90rpwZRLNgSOTXlhtDL/Uw6W3G1y
/gdGTNJCdgE3IkR2Q2tqg23HqW3R3m5RGEXSrgIBa3PZQzqMRXQ+DeNbl7AZ44k49IBouCM/eZRz
tuYdx9o+lEjSth+khTsVnu6cLiz0qo4uD5VdNv7zTx0szUHYl+X5RoD2RRxwB3HRsuVsY2oIZjeN
JgWyEEfcI28UiNBAn0lkAzRCcNJsiANIpZsUOEVoisTJVh6AMv9PhFGwGmOpv6Tv23yi+FxbCqqK
tL+TB94f4MCuRSPSO/DSC1H2VWI59G09pmbkoG5XIpi6Wri+dHchHcP4Ku9qIXF5Mu7WX+1dQwoS
DR3EWSJyVivzYijKTNNuqEhi210tuNoQW53RkiGl8ZqybuWXY0bwGgHal9P05XjsbBTGO1sPvp6o
/ol0SO1CamjscBxId50vDgQORZDgJMcD8l7vi/C//Q/j1b4D+asTreIv7GB5AYRwCR7BzpaIcyBe
A4HFbN16p5EqISj1iuxWZ6kyAsIFMu7tS4EPsM+xKYp+sr/GG/ufshkTh0UraIGMfQ535t5AplN7
dqK7efixv3Ml6kJsEXcHHfcE0aL2fS7wZntP8WZtnFBO5vtYeN5cpK2fw49nhsuV8S3RUpuWi6Nc
Bll3QWMRkbm5ofPDOPPEw21IWqmLS3JFQKmS6uloWlyU/W6qFv3TGqk5NrY5873WD+UyyBR08bXa
Z/xgVMbBCB3Y+jxN6/jK2k7vxxP7/DN6RWDSq6zwWDx/Y7isd2chyXjmGfFhL0P5aUgZ4ojTtMoC
V99gMiW/wAukaSusQd7qnzcdroAaDe1km/7nXu6zT69yE4NGXmLL4TZNVvaZ8zNXYevbAA7Sm/+q
Ll1ae2hZHrZbVZCJSUNvIrjw7vsOqAYbt5ePorB+1IQQQfmYATuoQDRzBcRaOdLum3BZpuwqG/+6
wKaUSDeZcj1IcvdwWz1Q7hKAWVEEmRmkq2qFTkoiVPBJmtIIBnsmKLBxn4KWUhayxjyj3JCINmaV
OLmu7YyaaJGWpWoCkrbCumfZyBzMC7erUaAT1p19HTcQMkB3Gb2KDMgP4CkrDFW1jr385zaVG0tw
1j5Q4TpvugckSGZQlEMveZtgmnoD8iJyJXnabYrOIo5wXh2Dv/5Ay4+k3esVYQkqrWZqk0RHQ+EF
Wmdu/ql7ZNbe8ZdBQjMpbOb9OUTy3OZ8G8SQ7ny3TJ3RLYTuSqW//Q4LcFXJUKihx2bc56iRRD/P
+wdvTUDyMss09H+izJPQ6oLTq1wM3GUqVD33S+r1882HLEE9w8W3AIoCShdCv8Tw9OPltFJpfa+9
38tZs9mCYMAOXBzydX/rxXxuDyZ6DoFXC9IxvaebsOr4PxvQl4oSL/MHB1ZccoQM5o8sUK/bldM+
3csMmOpxZLLNzEiU0Rt5kKdGWwTWEylzJb58XL3GHh7kWuFhX2RTP0BjdwS6qhu1QHJE3OV8NJw+
/pzbniLzwqbrovaAtH31VJyXPAT0OB4CwEF+p7Iml15ZjRaBADc+55wsYYTGn8Cq0zTtHOdIsjHb
OxpzR9GFeTJiWovuZuu79Jon6Kz+U5wwNeswd4opML043vkBjnpADAHhnlqpKVOZiLGQorqYmu4I
8siKg9oBNZqdTXNXpKeFKf1baziXzOuMHF4dCEyCX6kWRpOIOlO3jPc/trvJbIzNadnHALhZF1Yz
IJcA509sQE3A9PWKU/V+Dueo/WU/mpWlPe4RjB56hqGYNSIzc0oUQx/ATYvsW+gRphQD1H/2kkV/
4ChW5ggz468cOePKLvUb1tgdrPONViInpDVQ4Z3pzvzSaKIIGZbUNDAJOP8eHdt/I6zzlkWnyRkm
8AiQS562AF0YA46nyg+wfr+8iUKm/U7JNl2jnpFZ50mY2v+p4ywuzVevThzsge3RUfJ9Q7SmnBZz
9SlM2csfnWlNUkUi67ys2hoDewIoMgVZtSP1Uv/66PWoks39tVRaZ5yGNpEhfFx+Zh6DcQbXdO8N
StMl7o7TYyV+285uhrz6QlpQz5FvQakaCxM1zItCd0GO2vbbjOyKtgFssUkOz/ajkm/piSRbC/2H
vJrbuA4nqkRYSGIIk5hnxVnGcmfzgpmVaDLQsOxTuTuaJavjWgI+N4kNESXmsWlWIA/aA+aU9uil
vezGGMIM/P+DPGr+mqdWtB96xfVi7NUKM8CMlt1HFpaG00+8LLckMACJMP2YETaYxlm0Kh9k32bi
SoinN2vRHeKQ/snjNQcTqnwCnPPc2MsaM7K4Q25LpsrNN6490Vko2YcwmSQvBzXxblzYKCRjFFe+
MHgHojzSC7NjDIwvLTwFtpcXm52g+zCZSCxg+qdUwqeSGxiOj/agouU8fBXrLVStJF2dwb/LLlC9
g6fHL6/y1un3dx2WijA7JsSKlytiacMF6ZVLr0RPUUia72rXX8J5u4Jrel9FOTaFGPKYUYgkKkxw
OOdy86EdFAGySGXMAkOhMVIFXVCkUD7r77TsGCsrCNImE3eBg0PY3gji3mNnI/kKDMV1TmOq/M5m
gg6p78zgzb67wIDASYNAiX5Kr5ax8prYG1JPGZRurGr6GjF8cGxQOkEGAr7mR4RrQFGtN9n4kM6d
wCcf35nPg5/gYpPamfiaip9uCB7LKC83XV3kfp62KEWpVc1d3bQTdYbc5zwElKEnxBwM5OaL4Ect
BPhFEHo4cZpQ4OoiPVcltG6G1csqAc3IBwvWPy8ZPoUWsdKsigsiKR/vGt4vlq/llq8hyzwGMSwn
DkRfkSjgor6AWfVh+sqK+Bh9QBJLAoUrKI+SEoZkpoqpW6oAJ8M36yFedg0tO1rDxwEvtnGh/J36
Pz6bv1rylk+Qr2FUR8v/81RDLAX1UW4QcTPWoCDcytZmo1XRuYYK2nq+QtXlm2kAzAApizHyHcnF
ftP26I/CYp7K3EZ0vachOQKoBUYYcb6XluIN7QQ828lIKNa3r9Api0uxSQzPf1RGhNtf2PWf/uTY
yNoP8FW7toga/hfwqb3K6kR/w1EMJjpeHyn1RZTeyRtYtK4c1JFIbb4TZHDeeF2oeD+r/BrbFRIe
ljwGalO09kWnlHb51OZuKB3YOnNUDltTOW36a3KhT/Ng4kx5EF1iYkfkNwDE2vbWC/EcDL9+/bYe
jtwCaxFW3jJ5l1+GbIZ2730NfiFkAcn880GGe4eJfKNp8oBvbl63Bzdfl16x6Weqhxj+orbmU1Fh
Tg5ZIZnbwZWHM66a4+4Jlvs0Qyve/Kv4Lgdf7Pm5j+H9ay4MHWRTDhqFyX4lMs7oKFhu3X6gq1S5
avAhJv3EPKnSzq3WtEqP6Mz0I5kFQyaOujA4r+tjniS41hNQK4q2qD4+GuhpCplIlcGcXdMg8yeI
WB9R23uPMbzslEI8QceI7HkINHaAcPx1Ce6hhI/l2WCWB26ZfhhMY626lJBD5Ei3EbPga9Og3+m+
h3Th8OLN2Pel/s+sQZptEWk599nDaaYUXwH7MzZ0/clv1102z41R3V8FvXOuxWK80v3I/yc9HULD
nv7RiDPaCdpOO0ZSPm/GUshe5ECo+73wfS93Bkzt4hBHBmZ9Sv0vM9O5H8xmbH0VxuggMqEb1ehr
j7uVhGojrbTnlXDlaLo/S19BVYTHZaFReVqrt07FY9QMtyh2JlVTIQuUesNykaLNXN056+LobTbR
HO9yu0F9WlnpSNRap1YhmoPTKFRu6t/Z+TZuAIHwA/l/BNMqiTGtSICoUqqIvkZ7+KrP88m7vkb5
nMzVnHDmKInKpR5BMs8J7nxjulNPgBtRXqx94gWk0H1lEFAKB1CsUPBjBvZH/bp31/NDW1mHddyA
u+PHOij6hnB3cQAAhf8EVugBqne3j2JPYv+MNX45TVDfEuYnWVHNUkM9H+5yW0O4HPMepDnl3Thl
FHA2hmeh2PfCkYKaYlajuuJO/w+TO+8K/gJqKjcMWw36/eNICCPq3OROjrl29eSZRp5gvQtPFax8
B4l3HRUXRL0OROqdwBl74Q3GKJ+MOCTptEartGEsQe4vWEZb33EYU62J617nJ7Zf2upMBBiSvQDb
4N2JbU4xEmQDmnlQn5ugB0FFRUw6GP8MSRUfgYnqfz9L4FHp2ESVhh7zW9x+LcVH1mfFeVguv3tl
L77oSKjkUFUzu0Jc4YYpJBGfsk1xfyAddQoYOB6xT4jXZhba0RjPudfIM0aVnFxB1JJoAw46NQBn
j6lJebeC9PuLoxoNlkPurYx1bmb6A4SlX0KN1WXBozpoWgPFr/eCIsdxZBVyRl/xpxJqDZitku4K
NXd6KS/L8YRshW2oKVtC/TNYWbc20kyeB1HsWOa944PFrgwpTNvTavZkmWnvi5fbeKFJfa/j9emv
LvMBNe1LfDUeBUP/CCfHxxwegG/8mTVo/Uy3cnN9jVjxp6fNsskF41rrV6STZpw+FhqDXvqQ0iAv
ScQ3nKWBbfeOzSKJ4NiUqQppNrQcw4JVw7+nISFtSRFqRUc3LnhKF0PgzDNwSxHLsJy7NGebtufQ
/28MUW7SgL98s9iSStYHC31vJxy2+bQv68Ng+CmpluPxjQz5t8fLUZ817NUoqkxvlK9LFFUrJEmA
hD8ITXq8x3hw/gp96O8U/rP+ZKFVv6jC07uGfvpfFiEVxsNvRuMfI2TCp7CLXOj2q2/gocD8N7wb
HUZnDj4ZCQeDigCn6kMFDcDKNvMidSich72Q954RyzxpsYnSZTk2ryIJBxNOlpgmhP2kpX/e/STl
R1tS52K8Ev2HB5+Z3NHFKqn5Fi5iWxhqe+fIrdIeBr6zBex7o0NGmYsjyZWu9lHG6Hv89maqZwph
KQxL3ozP8lfNfOgPqNL5E+UajuPKTODE3XZdwUNrSxHZHFQPdiuLD5dZLcskk/XQ2QsGTfhuoFTF
PDqrvVFT9qks7BB7sps7w95XiRCgLOSdBsgYiaobYwt64Ivh/pYdr99tJMnBx3R3/U09CNoRyMsN
di4lF0Al6yI5lP84ObEAFmU2FPIkX8JuFYeNbCR3JaPG/50MQt25L3dITFqrTOoROupBLJJaZKvA
/P34qg7y46I1cEkN5YeDaZfMBk/vwjJUtfCpKuLSX9AB1YuJp5zMfvENt/+ek/LDL8Mz/RmawiNU
baBDZ7mTsWBt1FWSpLE9aSSJ1lFnk5lyC9uQtLurb3nloy/fY4+xqxc+7Vx439xSdKdG2cvpn6se
8/iHhJoPkOaPHZd/51I5fa+gPGYLEpM8UcQbfn23G/vcxCBqkJr0p8W22/vHm43aIckjLnNoh4ie
7M2XDvqMcTFU9sJa2j/gKG2DBb0KgasduAxoGMgc8lHFEaOuaI61hz9pdGm9qAS1Etn9qamCP0BG
9gti8zKpU7ESrEsrwq6D6FycbSynhcFCGddltSSprqWoZhPhieDTUXKWV4tu9gdWkz11lXS1HuOK
QcLqSggg0M6hKi2xpGn8M7TlqgzJpS761e97YYuWTWfY2HUJf9sxIsT8rGVhkCB9y/+Y/Hi5tHy/
c1SLGmJ3wGOfOMiRmHcAchkkZC9pZ1kffFXsqwiJgbXLXSBmiSucykB0oCFxDOzZHkJMqx8wbSd3
nPd8y+CGSp2IezDAogWWwiXJ4ACbfYr+XN2b/3R2VxjBnXiDNciuUWObcTskn26/VUK5Xp3qxjlG
22U2SP3bS8TKGWYl6QZJFWvMCL5aF/lPwb4tMupETsNgejMBUP/lsE4PUBP10k+p8N0G4AMNskZp
eU/AmDyQTjmmkqENJy7btNP/+qRvG5uECDaihygA0NDhXD4WwaJdU4SE3Bd0ORpLKGee8gxva6aT
mFXFd7wO9wvtl3Z7di1nP6LK/SPYa57ftmVW48rT9j+lUxqGoWPqi6rWj7mATPBAKCRl/1ItCFej
bdDV3VHlktHduhijo2ncfCnCPbR3fX+Z+KFVgD14yy9lFvFnWJ04Z8mm2+D8iXw7sBxYkb1udGRG
BS1HW29d5qaW1L2EdsLTeFBy5pYMJba/uRRE0Ozu9hN/6q0wutimFPoPNu0E/sB/GtXS0S7oCLZH
wKFgza2U1QsWt1NO7J3Jc59NwEV3g6Bnmz1o3kACrbYqF/1mQ02/t3RoaQhCttnKQa2EecCQKqcQ
4CuOQbG4tE79uaBcmswpLtLLnjdHGwSq5CT8zqknOn4DvgFzeZcvXxQO6svN0v9REryyqSokSe0G
j+WJQbSV86iJNVrHvGpST3JuOPx2UrEqSun0cxn4yyk/ts/jWJK9NpSSnJE7KXPKB21/HxE8z/H4
XIA0Wtfm5zPEsn5L8wtQEyft7scFIdpmh8kbpvcr4JW9kQH2uC4g4XatQTQ4ym74HrauqxmPZHfw
MTEI1vjVFlQ0/Tp4H9LGSKYxLm2qnTQlHyp38no/Z2Rxc28mU13bCrF4NaK45HkeeJsT+f+WosR5
fTcq45h9szgfBTMi7onC1wgr98Ved3WenovcTAE2ulzOMN3GBJsPJtsCQTVOyit+AFPIyVc6OPRD
3E0rEyFfqavpkQiQS9gTXL6mOhUqSJGOdxhtpvEz2G2J80Em5uG+m6xVR/YlUODlizs1W3F4xXmD
OWkwYAXYk3pmph9uwaITKCUKiGY1ZLsOMAhKnhw0SKO+v2WMyxsWXYb3kzRO2spkto73etuJQUlB
rZ1I9wxmt3gWLraR6sCLz9sHguQEjTfDxN89H6Bxf2CzZDZt+cwV0thxT1mHBqSZnfYBsnHTGQ6W
M7EIqn62ZFUEEvflGr1+PZ4Yi8eTJqvNbUFEnXPo9FJXJGx4D4fgV1Roc333mpdnnynxKZQrs1Rr
DiKWgeWFXRLvvIxDhkAG4kxarfAn6camZinbYM+M3SeVr6viIncNXxHmprDML3CCfdu6RNSQP3+n
6Rko+iBuHDnYgaL/VUBUiaJ8i1NGGYJF5hssEqzX5iWowmVyaC+/tW3DR1r1p18PoXGPzigv0aqa
brHED/NKgWjlwjdw+Qh+RJ8qvA8g6AXsGROpHbVIJ3s7CTMqMIO7h5Q7wCJTX9rDimNOaOLFPqOF
rbKit6u3EgJLdpqhrm4PGLu3ogJ7s6E5T4B/AD8kmMFkbxJ+PyyyatySCluvfvpoR0JCHEyFa5Zf
RYimWyzq/2e6hV8qPK6JXYUaM6N7MtWY9Ob70JLL2uVux7IhDJWROByQWWs5Hoy7Ee/WPEoBH9IH
QxIzYSxQ03eHpBX9JH2wRwxuBP4XBEvaVoX/aFYqohRgbzQduQtXK80waqaY+AE6REs9IoTTDxie
K7XHnKKL221E2KMevooXKoymBfXuNF/juK0Wdb6CRGFhmBC7rjLqayQWy93ApJCFqj+w269aKsN9
nkKs5ZGBRdeMPk1hN4PSD6aMuFcGlUpmUFn5K8o1R4pivpl5LRese2553NpE12evQKhPO+7oYQcV
3Gbi+P39tn7Z0wWcThoeZ3DbdrcXDZB6QbPUlvL+4HgvfhKEPylavtbe/reMUqcf25fEPc5/Ctcu
yK+G5xLPGiwWbY1FjID382ZpOGtIAEkdfE++eVwLOngkS8YtU3qZgZub25mZJZRbM6oaQAVw5ZPy
MtFtKkKHQWXEJbIACgUI31SzVjVemS/VXfl5W26qm03HHUSsvUmCA4mq0XN4kXR9FmZD1pzfOnd4
AbPo3Lgp+2VKGCm7oL+mbJ3ZODq40sljxJ5albQ1coKJcWjDG2x5v60BzdKQ97zNPPie+ZXYd8PW
Cq+JOp6/4bacu73PlNXwdcXHaq1LtFR9mJRhby9xTQe0a1Vs+2TLTlS6w62AUdQ0zE1HwL1rZjH+
qbEEJuZkRFswphepbDGCHLKnKnMuwU4ffd694Enc7pwaGBYeTBuaYO8vjduDiap2oVn3HWWkrW96
e37v5jFA/WjtRjLSPD/rbyHnMcqQZgRB2+NDcQFYHcIplTG5maVHJ2M4dqeHzGtl2F51akMD1koy
bHhvZEJaP72HkvdKsKaD2kK7xtw0C8CTsfExb38gIGzsqdBWSzcbsrjcuMGlMMnfTBaYUanb3t1r
OxSZIp74a0WzNA30DojBBlPZjRIgsghDM6EquMQZ0eauCl9XJL8DgraB9k7m5t8Nzyxo0AbwxmyR
OPkrPF+/dbS1uL/NGiFXBnZu7XI24oUkWbXxllsi9PkaTw2LCXZvdoaaZDHrOOc40cXzCqDsu1D9
W285T9idnvVyb1R7CBzgcCVxpWmPZTLmkfYKf6dX90fRKxRMS09MBYQgUbTETeUO3TwPwQNcWUkN
4Yga1rULLlUMwvv4fsCHZ0OxFNempwfpSM4PgV0QxotgZ5brzX6mAmzaL3I4W//gjojMoBHdCYYE
8QMbXtQrG2yGO5kiGNz/2474qH7YHSsgDMvaB4KvQIjfiFIv4zucfksgihQ0S1dp0OMiELuvHrqg
3OHHM/puKemExam/fJFJH/tVKiHogrb4dUUb9AaDARP130t5mmi2gdKGCpJsr9mhhXbM/pn3PmSy
uLbNOLzlL1fX9YK95LdgBWQ4p/llub9hUdmg5vXi4h6PpJL2s7+iOVUBi3XtqDCXJRf+r54QsxpH
i21+UAFOCA5wRU4OG/f2Q+2PM9d5v1vz7znnqfuYmO3yD4w2rVkQCum03nCC8DmmUAjq+MQZjZh8
3370dAaC6iIR++hWvIxkF1Pe5/ubf9Uh3NaTv2Eb08OCkAXWptwwT9p0Zh8S0cjwnZz9xEb6s60B
BfAqjr5cjmR9QY26k6pULZ1j/7CfJNOT7W4EB89YwPW0WZwsFFcZDycVbF+2RIpLofLlOH4R9Ekg
/l31zQaAjMo4Mk0lOOTMYvNbj1ULmSpAKgvypBMf1ny4h8dWM/IA7OTjP0/tcIXugQ1nalko/14m
aTBa3hjZlf53T96DXjwdFNmjSVVb3k++xD+j8J6xPsowMPx7gibLwnLHJaPcSLhVd/WdY6Oovehk
BWs1qiI1pGrJIkqhSMxdFj5duIt61BmWZ+57kT6/Wynx9o5hUlqT+G46WMMwAXvSxRpdg0VvBdM2
aTt1MSA6eaRVTXqVYpNJU1+l5+xzhpKe9AYIovf88QFvaMXr5okQJMUpcTu+eDkHlV1vnm/+qyVZ
WpZcCy/Ood8UwRnVh8/MeACHGFv4CAN5l3f029ppCRrFxdms9fHz1JxOAo9LwHNe2NsDrS0741Oo
OLL57upkbPm2cvhe/bk9MioV5PxvRyAOdOvfJClZtNXC6Vnay8wKVXf7CwccJDuj0r2w1kPnRWNv
eUGx3u+vOW9fcImHrBSsob8JaQhjo0hs1q1ta8APV5LV4jLZgJ/WY2zgXYOLjiCLmGNiXrg1ogpq
CLlKdoL5yFXBoaDc+Lyb6sBTNUIC2scZghoOCRXUWoy5YMc/DylPo/3iB6YLtxe71q9AlMyKptQ/
I0LYphKWCUHclzTpFTw7VrcEdLjTiZyN2VwUWYemddeAmsFWiarw55Xhil3MQNDqnZTBPFMPuItF
3mpb8rKJHjFzshZu3rDCG4EB8FMpIyBg73jx2ym3NdZK6tKPlEOvPEZWRViqpIMSAFAPe3u0bFyY
HKCjNhgDKxQKvxvc2SDxQAvDpDgaylYcgPsT51BfeZ0xYktUFcAxuEnqehoYixUfLTu0RmFt6SqR
2zb1a3mvhwbgvIpuysrPmMjGPZIZpqCkQ4dizgukBAZvaFiGlaYZobgoKHvVIZrOk7fGT5fINGnz
KuERAmNJCURhfYUsjNVMl68Y0Mh0i/iRYPmavKAr8nl/3RJ0nqIWli5TfT5ljSR75F3d8EOVOC6+
O5wVOUtR8Nowi1fXjlkebyIsK1JcpwodV7TxAwDEqHxx5NeIjadbByn+JzjNaOMTEtoowkf64wH9
L/AIW4wDPtGv/bh65LJC1pF284k3EIaUzyTRm6A1vrBB4z4PUbjWbsUCIFWhlV78K6S64i+PrT8/
pMQzpyWSFICzv0LDeuQBfd+9pmAaYEPVnWLfMbI+9+Tqilzb9VOONQZZcwHNaDtNY8Amf8tBPZFY
HcqmPAwyVuQqdNr2owodimAzti1eIENFuHoIDE/7tt8Npx7dtbjtFMoSrjgHPyoTOW6GIPu6XWxk
wSA8CwaTaId+yPJVOTi8/gtrL2x8xS2OBEmyJfDd1jp7Ka/7unm+FsQL2SJ+JaEqVLWVGwmGJJVh
2NtuiAoBEIg0xZftV6lL1Acd+XALzJ5doStzMH+OVGd1bvMS9q9Qmb71E4yUpbP8ct3AGRXG8swu
2TsAhFIYwXl/ATmslFgDh2S1bYVCm5tm/SWmTYjESD/c0Q2levT8LqhnXa0JIJknLGi3aXaUV7zK
I5sPCup1NcruUeWawOYAOSXsuyW2rMZNxkmX60S+39W5ktKQFFIlwIHDtVoJfJ6KOhJpKO1/lT/u
40eIHshgOBFAVyYu2uPJdpmolZ6oinBzXX+6P5eFb/kxHG5V6Wz/ToDpEyfrCt9FmHi33Z0jBYRw
yJukTT7G5D08loU+oRToYJ/RS6CbM19xREFzJiq0tC7gJmFK22xIWf3ls+Z1BzGgCRjExMbMmrTd
6IiXrzmkYSCSISTWs2E7tpgG0smxo29RTHIQKgXHqMjcyhLe7V8VLhBtnDgRS3aaxyGCL69Ee4tD
UoukSA7xi1GOLajKM+e7hfflIeQDRmReV+5KZuFfDfgr3kmZKXz6KvoJB/oe+ijJqiuATVmPb6Pv
OLIYlciZuCu8cPfh5ccv167HCagcMVm4wTMCMOghS00B8udpDEVRCYLxckOVSgKXHkBodFU/pp4m
427PmibFpWEavX/41K+Hq29ipWa1YA0SkSxNjfQID0S69ghO3vKHKAQOYtlQFbQRQbGEvXN4MYg3
ORSMEx5Mc4BUtmlgPu1KkYSFjC/CoAkU1iZg5Zu/jMfxD5FJjCV4LCK0Kt7HUVQbNHskWAqg1ZI8
Yxy883/kHKOFnR6l3B914UrEbux96oZ2MyQM2q/K/exHONNWsmW4cNdwa0cqM4UB5n3mSk/LpWx+
2gUwnC4WvGFpFtwJmMPMakLpR9CDomKPcrNoLmPnvxMxGvQLgRk2ZusAVe+fuKYnk2uCXTjMQ+Ie
+LkrApZEeGe86FofCtFXGKFCceSffABKikFISoQGyfe07xAB/UykkmFDPK+F3hGQHLTDTUYab1BJ
eUEsIytvVPoBSlLa6dBMnBiQ2WJpRVu+u7A78BTLB8dRJem45VVGfAx8+A8YwRIDjjC/VAOidomY
O3zCS8oeAxoKcrp1uWZHRb9pEh7CQUOQlaqagOjek8ZtJe6rorn8EPB38KRSL9xSniRg2zy8fPRN
F1lAsNXFW2cO5JpYXgPA2LSlxSuQePaHq89G15iMEFS4pnZybxsTQErD/h7Woc8AInfjIMVxcbTZ
LYVmEVGqocHSWV8qVutY4e+Z7px5QTTKon+lyQt4k1r2jxMHKW6ClzEDY1hgqdKjYxYFmECVhImo
86R8Iq2MKQZmwr7NIg6s0iMcbsQT/iZPHDqVLOZXgE2thDFh92Vr2drYBz+wXAdjIxrqrSHKAjIQ
je9XEwQxDiFm2t4e/+47H2sIrnhOH8IXvsimyaIXvzukrgBtC5T/JcbShwbpyuhgt3XR0FvTeOyK
CVh+FQEq/4EMSXJL4vJVeefX64jBHOEZeDVgqnI525zeZbThu+gBGWJTYUikgqSDHRKNArfqZYZ8
e3eX2xcFWs0oBboAF1t6577c/YpuggL51yDl2bQT35wF9TjvOIxEKiRq2snYqWVkjzuOGBMtJsw/
rYx8CS20N4bGTQZqFnjZ/+R2qupOKdyR9VmWjD6/p4Agoj7GdmKQ6dk10tp4+SstZZ5Ehlzxqt5x
SmhoD1opCc7kYamDucPzH1PXsro3tfyf/UOuGk1Sif0DmtXEADscR5UhQCE1GHm8dOgfhgbm2qwG
l1SWcPfCJKbAPSJkgohQv+kBrTOFRKAe+19HRX3oQAu1LiCh1rzbgbKu/yGGjI+8RGEV70vVKlXW
1xq7dCdBiHxxfnju5A7nPJ68Z1gdMeeWszJ7OMpkbk/esKy7KckN92bIomYwfkl1ijM1fuR4sWfl
96/KcMvaBJmUmu35PbtRVjSKEyMh8slNDeNgdiN0jYNNVa3w8eqfO3M5NlcKB5TPH4/6HP9aaqdk
SPL2tEbSSiLYTHyUSrkjcndHZScQ9324tadbzsEtImSnEzP5OTqsh5j+/8IIuJ9WJELhFwBzBc1h
L3xo4tahJISXeiuJETinesNBer6GXAPms9eAfXxuleqJ+ZQIHCyq13gqsL6+6vgBRw8zN59cGiUw
l8GIO8xv3BuxMzILZQm2Gsxpowv3kleKAg4Zf0cTbuvUqMcjev9YKIAuDFU51kNyUfFEnXrLmX9S
mQYg3HEWSVMpMqfgLDqq4lfs5RZWqosB25b8lhDoSlJ/18Zg2ZVB+Mp+kkRlL9dHevhUfdmVBUM1
o+zfJ8lSbh/NUJOSKv+IeBmTbBoA42Wi7LN55CDGrNweeaHwkbWWYYwNThVViPnb/dJdR4avvrjk
FF+wTStXsAjuWwcK0YHpshmLgRoAhu4sO3fIprpGSviYy1zplIf2tKWbiJJLLs6Q7C0R3tomOc0B
BsrPs4suK2xPuwDHRf+9vH6giiRX5yW4ULXrqtvyXAwzHd19t5Inlh2naCEnRUPNCBY1xYZ8/I4Y
QHFCRXZ9Ngu7nreQ7uN+fzm4F3brDCrI4dy7XWsFUfqLwxFLfK7fa+fE/Xkg61byVdVTv8LsULi0
6MfDxrjgIRlyH03rKoJzzjPbWZ68FEVpOBIKWG2k78R75E6a8TOl6AgOUlfnug1cvNnEdVkos7wl
PjQiSVtzvlstnvxSXe1fp9IL3gtX/Mc3WZomMnR9hxnslGj0SeO0pf2QPhZEjkPQ0L2tLP2NnnrE
AUFMNMOeVmQwxXoOr50WWBDf1ucVoObRrTJiI6UOC0i2SnRlQdKNh1eqCp+8rkoaSggkimk0ivWw
qpFiXGhsbon3qJZeyNcAWpsBZwBgBjNGbTOLI82BZYqMyeH7KACUBEsIN6Gq2t1GDS2eRYJ7Pg5s
b+/Vpod30ibWn8gKbbguXMc8WPp39nUuNIG3Y8Wvemt1INP6ZkmAxdZklC6ZMUPrEMk7xwKlvpet
Ry1iCoTLROqiqiDphNc6FL0np6p+zHAyjRSmjgvJFp/Rn4Gv15F3A7cJ8ux3ru+VnSaRzXvHZpd+
YPFLjLmbfebZDOtseUiepJAs/PS3zxwXxv+Lp40yaw2IDHP/S/yxQhjNMOLymXxtUcpXR7mADZWY
78wwjaClIW86yOwfAjh+oCat1f9+LfEkwtXMt2SysEtEf/NEjpDsQM+W92v0YIFT7pXcidrKj5X1
JItgMSmlQ1aKU2qAQ9j9QR4oDIT18FYuapxgdqy8heRAM3ZBRtKKQwGIQsTxGkxUd7PO2OF+TcNa
s3zsEoOHyxEEuL9TCco5MqdQ7nmc9pjtfMqe2HKV6WM6Z3trMIae1FaJMhMAuyNRhJM95zL1Qp90
q7eAbf6KqztCH3HO9eF6YnFegz6upCtC5GdvdTWTLJHQ4H6w5sNjlRA83IHavlhPYvt3hFkoEr4b
81a23un9FybL4CU6WnbejOkMGWGvh6PcoO7u4XuDNdRU7gChDW4I+fbbYpjbGxB8lWxJIvClu99H
G0hqeAjJei0cFDsxHZjbvVPS3knufJFECe8seRCjTZdaHIxKjtXR6FoObZL+F3t5KXVlR2OXN6tu
930xFigoOv+rK4Lo1Y+Y10i7jtY/8tEFwmGTGSY+oLUA3r0dxESvrQwQiWniXeDIALCQ3Est75eh
NZQSpGjHN0PshSQhH2yGOunqR/9AeH+AYNb+LkAeOLWhGULCYHFFz7AjCtgoEtaltXGD0goA5uaz
19ZYos1x88v7vxNxAYh41OtTX18+KDrNmrm5fqtA9SArEY5vpBH45xUYJAhZbUsqDOMkgatoLI/w
F4l03hAmbcSl4yViXARDbN3p6UzI3VSIvySJPWbGreTCF66wjFjGMKZNUaxJTmf20JygARglntU5
usuS/HQVJcq77xTGOcMAXdZxEv8YsiabBbFlRiIAyTvKElUfaXx+wvJxH0uRs0GH18w24OZV4Ufa
BijcrajrI0GnuCnj6aYfUXhIQ/KikUnKdEb+ZqvMXGkuMwNzmmsUG/v11faqXxwDsA95bU4VGxvb
Pp1LN49J4tzlsdJTdc24KZyMtJGOtu6qCFdSJrIw/Kodzse0kUiKULl7diuKJB6goVpXorLfJdIv
I+E/hxcgBINYSPqK9yCEwR02icOgh9qZm94GyCzdbfZNPUYy7A8Oo84FkASNW0g6jAT8k5sxcmRk
ytXCwtzJrBWvdnKQuaRTc2WkyNkI+449vY38leUGsxOandJlwkZKRc5u2zNIYkkRmO2f+EGeM5l2
Ka0YGzcdPz3aSeN+mSBE1AnHnkmtbq/vvZFa6M/9PPo3s2KHipyD7EgG3wfxV3Eubk6Ayn+zjJJg
nowPmAtOttZQVugVLCL5uZluo/JZded+kFJrOSWhDZ2VHVKZq2CE+M15Nl2b2RtoYWYK69XmQqJ7
/VEKwmSTTg+HnVdI/STJ/XdAGYpUU3gyv+75QxtvaOQluOqIHupK2i3X0Yy3/4RFnrmn6Ub5OfJB
mPM419HFw0b7lJiCDJK/n4Eg/HthsC/lf5M/k1rZxZ/ZsM+exzsCCWBH4QyIbO0NADBWWGvIeiJs
2Cvzpodr3lKOpFDXbL51yDAjlxEBcsRXNWeI1S7w8xHKYx291i+kr+wtqXKiI+XFwJdN/MfJzrF3
uB5a+gX1xmUuJRMwloCWQ+9tuN2oF/GoXB5dXM+0oo0oaheW7s7tKr1x2p3cExU+eJvDBtmqoL1k
3olM3lwb8sD7XjtKoSXLlbwzt4jMXqDd3imfTJij4WXE7ukNS2K/7C/ddVWWlMin3M3MnKFjNGxx
WYVwFk4PUhjv8k2WbC0C+flq+sKSd/KfH9RxtVT+bwaFt0S2WKsXXEdKQwGQDZsOLcVCV8gihNw/
MsUx3sCnsSKyXPzN4Tzfr2yMVFT4uHWkdL8TxlBbQ7hSsqiBqZjXcLX/RLGXCJuKZsCz8PvmdXZN
iFZTZetGoiRQ7g7CgEtlVf3Xyp+6WHVuh18vEb+oZ0LhHFdABdBrno6Gs8g1PaiN0kygUrZmnwmY
6gDbz3NK+8ZHD6ElRJwweqPYmmyFDiwX66v6hr8mClhkGKWcqeLyWTLWirm8oZ7gWT6HAXZHEVFy
m9Sy53nFxbetOizVxrK9zJa0/L4W1De4ZWbjm1REm7DVsUKTdd+tGtp2zbfQ9bvjMsHCPNKfLtxM
noJPgKnV4548ibSbnWtciqaHwwbAQMhhaopc3F0OJS1IXKqCxBfOU039U31QFy41v00U9SZqjYJr
+fnQlG6hOPAMrbVBuuPUK/LMoeP1Oqh92QhnPXicPOOLSugR5ZbkH6tL50nEIAsqF7zpy6v5BBXI
4o1sqSh68+7G8k298wVxnFs10Z7QsGZLCjeSIvl297o5EU40meEWsJDJrfEjWMboEzNziuXrPP3/
RRVmYBRvZkq+jYFGWmfZfYAtTLXFnatslfKylnnf4BiT90hkUUtDc1aNgnnchXfXK32jD2SVIE8I
d7k39MhjB/cMBGrhL8Q2yqLFuujJ4Hi6B6r/UNs5vj+QcDI6/L3OPnHhxQkPwhGfImjC5tkq9Ypv
4QkWjHVV1xkGHi+ZbZftLwAH5CEbT2Z7yQoND2nTewe4krHNATE/oHZnGXtmLZ2mg+LAEZ5shfwU
QrLtlzrRsRy0LFttkdZsBFT0NkEDrqY2j+4vs3JmEtkm2oJerMMvUS/7o4XDd4zuxgyCubedv4vX
XFYqpCXkgrNJ8BSjHuKyo3dSveuiH2eO9mrZbLcS3NKziUH0Mtv0VMNu5pNSGCWM4Xp5/x0Pux/C
xqaAQGwzqnlPZJdo+VwDgPBBjJoLAEL+FSc0ofbBXSxGvTKdnZwfoUV38lJj4M9n5KBEniXu3FMc
4XhGXS8rtsMR99wpKkYdB8PqZYzhBGYWPYyXEC7LhpvffSzN5IgLNw86G0mkPZxMqd0/RxAfnHxs
ccAEJCEzBYPhOpcewpjbZR/dqnTWRsZqp0QDIgQCg9MAsA7zcd8r4EPvuGvOWb4d5vv4PXmNdggR
mylT4zAVMuT3AOhMsGCYy/HUGhpF6vDr5PK+8hd/DEbY/4RERsUtS/iEsRw4450576m10Ft+Jwc2
nyRCodt6FclDTe2OVtLK8ICDGjoNXhlRwkCC2enoSnZ9ONCVI4Wwa35eT7nIwHoUOGQxh+cTLrbk
GsYu/LsoFu6jr7BT7NDus9Js+ImoGtt+VG6YH01V7qdY5C4H7mto7qy58nsRTuBr9gcX+tB+0Hs/
KfbbvItNCicK+/3XU0IJ0e56CqerDrq3zvF4WgAhW13qzDfBFXFYLYHMP6QsOaxOJ0QLZz+xpGGZ
KX/3sV9ftkXZBqB3PETbaKVpnXrnA9Q3DyxbL9vaWk/+oGwqx7lF87cU+noYS28A/rxozqx2qBLl
MNaIDYM5lgbATxDuFOFDMsnilZFO9sqJh0BfDZC9yUqRJY8ezV7zq1rCct+aOVpHDSK4Er78AX1W
E0zagd1ZLRfs7+8qJ/kTPxFOLITttFmitOtyQqHkSzpCAkkZWJVQMgCYm88jXMosKOPtPWKxwEiM
geIIYsqf09DRVNnyM4WAROUJBN5ghg/wD9gQjWzYmThKLgQfigV44wWSMImS3eTql6P6aCVwMo+D
pkzfHbsU66myxtr0M3IKRYNOjyqSqUKPBDne2lhzkdgOEhl0mKzz0fPYdyoUCbiHYqr33biSSmtQ
as9r35t2016KXHkkwqmeB4yyQ0SZvt+1WgIVC+WpHzczb8MnMRcCKRSDDj7l4aoIgGRrVKaJSSSV
odfvsXt4OYSeV52bnVd6PMHV4Tgd3Ato2uVcTjOVdL1KVwLO9uWtfgPhuF6xAuI5rsbnsFTEp5X7
lDlhKhVAwMCcIRRAjXISDT+XD7srI6x+exU2Wi4bdpkjgb6CqOjMN7t/09/pCXHT/UeHkXk/Mxdo
va+3vcOzoH6a3/9IPXq4eJDYD8R3og5GeITxiNSiYpbgUlx9+Vji2yrZV0YqwMKphYXfNaONL1Dj
g7PinhzCNK8j1SB5lK4tGBJ7nArOdWDgM8RMsH7S7DLdGn9Xo5mQfFpDon21QPnh9jl2JHEaR3Oe
LtSGqq/h89DJW3e6SvJzGV3p055G/vvD93pUqfQnnr3tfZLN1osqicR55llFxySQksVhm0VNAha7
Z7ncZ4aqSW9keo/gVLBVYTvv+NwrqAJ6iW/bk6UMWRR6Lt9tEsGmFeh1eByQuUF39GaL4iu6PTpp
nmOxe63p6FDpDfCwa4UPP1LRbCVjZbcnIyhjTySeDUCeofCu3JDzMU2mTYScJwoncHGtUIHcMxNx
JOMLyGSs2GshD+uXwkIVPgsqoDPpvBgwy00cYxFTJVJZXc/QUSjK6/cwQ9iOuwplNL+HZGKZQDHR
7f1lOKCVUlLGNRW/PSLjPrI/GTIwDekEs4ZD0fLUH8PwCV23Fz/2svco7ESijYnlCry+glrDXjYE
k1BCFpTVyVMJsk/nxDhb+/lLCBgwk/AHkpKkta4eY0H38pN1DViREAZVJXBOvFcgw0y0ZKTpyE2X
tUq7bG5cXb0azpkG0TcmBS6F5nH1CpdPusT1T9yTYD/2E6U1jOmZM2bEim4KcZjn+PLj/OUw46F9
NExD5gEylkWyEqKZApnxQyMHBUYs1S+hovbzO3sDViNlekLm/7gJ136D39Fil/qQh9zVqJwV06TM
WEjgVJkvQvKg3dJQESlKhmJpy9ATznrOQAefXs8hMNKY479lro8mB6KWKQdAJsPqigRJJnsS3yOn
LNEH5EdT6xeLcpjMLnbSLETPIP8xDxQMJEuxzXaIfv8pjgtQWnhovrsdTXcw2vakJ8kQ4DGon0Qk
itsR1yCZ5Duhg41mISye9vUhhDqPPzlhYnThd6+4bQtvZDW9PlPAtg7OtTxWDBF8T4YRcmHSHSCB
tiflJrkKVhXuTzx+ig04DAmJJuigivWHe6bR3s9V4WxAqHRDmysT5CCI1trOyQrW2nckM85pCKz+
/BDyuuUgLggB3DGY7s19pCD/T1dBWtebkkYnl6/SRqDBsluq3Q0fD/8+WkTYJF/fSdf/aUcB/BjM
c7HLHQqu0xf8SAIh8v+TrLeyKq7uwpQhAIit2J2cxXrexMw48Wsh2oYKESUVpJu9ETLlWzxNdvXs
XH1f42toV50lgcffOkIpRv73mhiAXgmyfwwOYiKUbtu6Hra1pzzV90GWbPpPNl3DASkZwdCIncYD
Ht6tz017a2uRwk44Z0XCryJQY8gb3t1ueaPd8zsBtPrlw2FQl/vOrZ13nP485OBxYH6IYGLqvtO/
o+f+YtUNylFdFxpUC/Md7UbIPxYjzAJYJ2nCPx+WNXfZWF+KfRRJqDzOxZfQBadfjsCz7FclQZTE
p0jZlP/KKj64rqLh4wRnLjizFMDfD+rIsE40Cm6fwlXni6X4Jd9G/y0nuvO08d7l1a4AP7vhdDHm
OIE7md6XyMDFTYd2c61FI2xYTrQveQfH95J/TYNLcdgKMEhqdBzsO4rHPMsgw5Y3QGLpPIgtD0NX
n2drojrfdBsnERjoZeaAMhbDGmqFHPpw/NegkdoChywLJ7bleUKMWAXCMcV2BYHgnD9gBVfQvOp1
l5sDkerN4NuiJMwrXATVwZtL8cwkvs5DyxdUZy7SKNemc1SpfLv6NWishAL1i8O44M/B7k6hqvxW
ACWnX1o1RrlpQ3wbto3SIoM77qUa3ogtss3wIe8UuBuu8rUiUOsZg5yRr8KWua59XrjKYp02IfsB
o01+9jd0LUDKWtLywIfpbSqRTmK+J+kFA2PIrmv0eCKbukuB1H0lTBFkGwCt6phN+E5CvnvJ/bKu
/+ZOnZVnF+yMPP4ckkrmV/qmwilVCcB4iQ3T6jafTAVdugqKQkzVYtQs5QB01+calAZrod+a+BIT
+ai7NO0XQ5fd20ofLv8TH4+ZAwBNgqsRYHBJ+OSpXJuEbiWS3zZZGW/VDgePensmUDlPGbwpLqKB
Wh/OKOG1PRbR25WbZics6XMRtC10nVgZCtCdnx8Tbufv1nfXcabzfqzqqzCHZXI2oaDDqLizqr5o
hDdNRxYhGUamBxWBzx32xcq/1TDYEyc0e5JMcNfVohpcIoNoSpLjm/nCoOfflv6qJmcv5tT/u4I4
xkRjyUf8BU3gmcVOuWqQaVS454RH3sz69otUPZnXbsm3VrJSg+k+GPS6Gw6INfv0b0URjKRbNleo
2G1nW/gmrSkPQyloG5uJcO2DP5cPMuwDLc+Wr8zonMr/X524NE55rKnhnN43USu3YVkxJ8xQE0nl
Arn/cY9iMmeQc84cQjFE80ITg939RxZJR+thU6XJZQM2CMubiYdEDaTMledCmHrqBts9AmFBEgTB
MPna49TEDiMuNtfaOvTM79Bn1ur9fiYWgQDbS09UanuNu1UDOdyFjfvoszOmcNX2Stw7RDOyBXnz
nKeC6u5ENeRT7/GnNnpN0q5um0/HI1TMTunjG7e/e2QH6ZShetPX/ebWO14xvPEE2COK1iAFbuqT
XOWIkUt9OxNWTmd0yisLD9GTC5OO2JxJnXgfo7nMwlMcsH9iS8ShJIl7r4RQBP1l6RFqxDKz1pd3
g/Y7niJKl6/44SktdZSI47YQxebh/lWR6AHBKKDi/vpSvJmYIYlxKX5MNWpnfrYF/4gyPnWw35rj
QOcB7bAQ8Le5itLXjQcXp+1qgN9/vIfZo1aasViJ3iiXTrjr7dhucV3mhtS9oMvq28l7cB/HPJKv
xawu/mLX98HfbxYKlYZ+9Dn2BIw+fRwu5gaddlpTe9Vj7V8KxLxInkA5fRM4vJ302uw61DxV9/A+
j9IUoJ8zLeZMBtJJD32hgB52M9b8sYAmloJZz6BfILvFR8uwqhTMBWLXwEBUbnXuYjgwaxNJZhVH
FXcwibP1wvlH2vj4gYTxknsKYY2gVnZHH3lDnV16vveYUOrCLOUbgk8IN0UoVOgfPpYr4zco7cxk
inYutuVicmK0mi0WoEDgjML7Te6eH+XAQ3IRm/2OU9NbYUJkIvhVHGDA63P/2E82QgCWjS05NjQM
ACIp0IYXGvs1N0Xrb2B8LnC1zLPjD0RSUUv4GAmJKzTDgoEZu1jJHQLiRkzjatqT09sJhm5Y2Jss
dtEyCWDAXuQlx/5Lr4kaTkvOTNSQq7EjkSnistBSA1i1Qs8wHM6sRH4EhnxL7zkvv/kImRVt7iJa
OPZkW/c0BvFHX1OQmeK4n4TxUiqaSIw3AzUYwsrrff/gyQBdjkr/RE+LPXiUO0fttZRrJBVIE/tb
zO9GX6hbTvcWQEhw667dgvgn/rorbK47IOU02v627y95ubDK8X8VFVE880/KJuR9VO8T1Lwo3L4G
uXwL1iIWF+ZS7veNbnocLLqqzcGmDRZJ/duh2BRiyUIMuK9elEdSY7ui9hP8OZCAetmaqs/2bQvM
ZQysb0OXAbU218oh1ohgNHwbXC7n0A3Ourzg+3BZVQ23Qghd1CC7zs2LW+yjOfq/T/OYuenKc4nt
dl4QFxRFwBJWEU/Le37RWidmI635xdmYLo/lWcFdX6pI8/DHnjF90fYn+HardNIEtlcM8kDXHbTU
68U/oRgCDEz7uePQVvzNVWBQkdgJ3RVXNiBJI0yPyDkJ7uQ30sM/5oRHOhOm4iktRGaVyM4kCBSu
mqbiDnJbYcvt0cmfE2XXjW6+zNnXld9C1DYbgRexDzH55WyysmtFz8KTMGhyGSn+yfJGCayozlC0
j4UsKTDXm8DtR0kwavNqqVxiRrUd8zRiPLXEZIc1Z3KYk/vY4kCPIshfy5XRyAQYue00tyCIYCLd
LMLEhL9TrMCb/xZUwZoglgBHgcQOY58GOKo/bzBJC8cXSjFGC0gqGtCLy3KNi7750g3LNhlA6zY7
2Uz1tXnOLlh7/xriXtC8zjhDN37OibcOuQ9HW+BybgbhgnOCQsdpVujaApeOksLGroOnlBRbra6p
+Ha53TIc3o6rUmIWEYkYjSNCScDT5IIaTpqGAHPwatqGH5DqkVnxyeshnsPdbQ5M3/F1xGZUHoLs
s01qQVW06EKlrQAjTsSPI/8HDuuoQqKPiw9ajH25kPaLfYB2pFp8Yvj+N2SLmNiYS8QTM8vwtse5
nxge11CI+wCZjZFjm6dKh0Q9AV5H5kuNI5mUFGbEac/c9sKGNZcfI/dp7uncvfv8qAnax13XzoEa
/3LEkDQlc6ORd+Foy1K1DwpCEvuaD/hVSpnKwex4/poZsA8Pkxqa73CGW9XcwvL3Ej63iQ+ARLMT
oyUn3KyZEdJQ8izHEzVHlFhpjmWgf668HyowWoZiOLA6RQ1rLV4g1nYVT6P/jy64pLvrISemqzD5
1GOC/eM6LNOE/xnWoqlRx0q3NZ6PgOylnfzGNAn2ylqeDnm8vOxZjY5BpIh+qpGkwCWnqkuLhlFW
l66wFJNCiXq2jlvn8lUiTkPuXJNor8yCXQs2Ed9K38FrxHZSeIg/0SckTu2RuHF+K2gAwfuTHJxP
m9IQx9F23gJ5ol5G1bf/1+LcKQ5Fp8PRYguvtJup5Rkp68Ujgn3cYb6pUwEhCAReXVhTzA1aaqkN
qARbbQIRDA5mEzX9sXMS0HSXk2zT2u37wm8jiFct5eVq/jm5WjjrwoV8dnGaDl62yUxfCBBcjNCf
ZlzT0EyFmr9g1Urrl60qm2r7QOU8BqewND2xXgTYnKTKEy+Y3tFX42/DDFD+ktsYomF3FhI9BZVR
ggsdLNkv/oKNsdajuHlegpIscsKsUT0Haa2BgIJkEtd5mzf/huEXNqjsa+tM0HrGmNlC30SDJ5IG
pIyHuFNhpYOTKNX2MKvsV1/gUXkCu69CkAmfaRoYJ710mIkLC8ybaQXlS9B+AX2DHLQK1TksQKOA
64jtU9nx8woYiTmrJIiVpzPHyokksmptE8XtyRN7NjUek1OtiONFvPkzhtK6P1OYrbAlk+pDA+X/
f+lnQdK6GV87fPo09JfhJqNdBlEcSCBe0lvCQhM+aEmq3/qmUOag44EsNOQyolIIsLgTKwmzyIEN
EMXrOFOnbd5tzF8oTeBIHs61fxaKVDRCi4yXUfH9lwoI7bxsf6s2pSC13fIJ6KR+YuZOsW03AmSC
hrPY+bcMQ48eTgJ7f797+92HylzC3hVH2V87wrBc/VuQA7oa/UjCi7uDKms8qVnNsgDZKDuC/HIj
7opfLsysMupkImp9wKfXa399ltHTHtY/RQcESYb6vG1X2yvh06Vc5ZBoIQpBk2CSDeByoaZNCWLk
gPomHAELWpTpJ6L+H4wnSSXYzDlkTtXArvOwOXsMJFxmpFIDlXxqVUy8oVjosBLF68D9jmvWGxXp
cg6kpX8H1S/0u0/MsMuORuP+JnBH6V7ATrVVvPoPl3Zw5PCVYeqvhfT6Gp2FIbfqd/KAyzdLWZYk
FHfMubHfnzIFnF/o/9PkoxN9JqUx5mw8pqmANqZKurfgKIjvrnRo4POgZ8j1ij75+Hxxkd5ZHT+E
qZampf0+V8lzYv+BANXq6XraWPlR5LmEzaqqzNzElRuOnrHVms1v8VLGbpOqe9ItbtYur087M16i
3+yFO35xGLHpftBahslT9xek77OpflKN6o5bMagq8ZbIxHlSyBR94t8TBl8wYJZQ8r3r+tbCOfwJ
xsqMS7HaGMmB/7rHN2bpLL1MSFpVu2KPd0kBa8G9gfu2JZfyokEvfBZHnWBUjeRarGz/HDLB25G5
1VbkYnASprFkQlzt3HG2BITgBZE+OTrfOrkWq4UmWCZ4VYXmGaprh5vuTK8V0AFB3+lmIWqESCfr
BkoCKV4An89phcCR6BPz799F6T/SjEMNZuEd2AejYSOHNXW6DCYovSppDcMUdjyehNcyJkVrktI1
Ti4InM8TubKb8Ltv0p7GsZk4Kqy/WABZG7hWlaaBxXiQBwKnplX0E7fW8Nks3PHTqVWRuzzU2XmJ
ivR26tEDh42uyZ72C2aXLhNkxbVHaTaEAnEkJyoid6XCNXcuRY6rgohl9L8DLnbX4Ed6FCwXBnUr
Sh65YMMlbIbrrlhi76dm0fmyF5EMhMad5kSMZ317XEfW3fh5Py/+jK/KafegGCHdmclbV2jc1QuR
VGmBMi+GsykLpEydziIBLAS+NuQP002rbqogb+GBkP9qmkfZTb+27CETFEWy8fygdR0/rrK8CMBn
B55yPEq7snKAVxqpLh0Y3LMo/F0eME80c3Y64X4vZd1LxAlJ/6DIcnwHfFSqFfTMKuA2dS8L6zgx
OEjFOAQbUkxmz2VBO87AahR0780I8Gkm5nOncP7y6/Zk3yKLyeSCbyPFGUA1+KXwLCpD8x8DRihL
kqIc0xEJ0awAfvBVG1bP8ACiqmhKwUhWD07Mrt/0699k9ahUeUO8SVhz3p3IvGAAWnwB9Jtg1P6R
FnDOT8iZAtSt0l6RvnYjmwjq2cez/G4L9SrZOKbi7QrtscwKeDc+2rlJnCGPhmhORbThrKdPStN7
NBHpBZHjKJGnpw7Mrhqm176VZafM3CaNo1d4s94O/rctqRG6E3gyIQgzxiMNL16QXk2V/HGAel9e
AIKQTFBt5ImlHsmgr5CXgUs3OBVUJDeS2M8bKPO9USH7Y9Gt66ccnCOIUW10BT2bzdvxkqm6Er9t
wzoWjATuvZCNhocwnBCiDwqBRqoV/waMhfnxfTA6Zxkw+AyVAfXw/yVapZglo2mqaeD8uy0SJ07g
L6fxVo6rL8W9bg1RwLovsZZlHA+Z3n48xg3pVWbss5FPGHz/uFCV//ldqjfY1muQ++rxqFbGxKsn
rUYscQpk2JBa5/1tYbc8fZs0qEji7nEstGDNrwD8ETONkOvIWbeYN96OSUCnN9NZefDUrA9rep1J
b6FDWj0fe/ArYcgnccXZWbUmhvXqHsJ2qEyeRImf7EE2nuiLfBVdmEduamyCnPKShzLjW7fC6XJ+
BWYNPHgSgXjGNhbjk9CFlgXHU2wk5pkdUvmW+KhQ68U+EkIinZyQHAYKm1olMABBShFYRZ6rKVEi
4IeGXy+3Z6jltIIVJBq8ULpE2EL5UFoQgwMxGFcNnvNxkcDPEy4dOMxkGWa15LSkkzR2VibHluV5
55WsQCzoh9kWn8zclIMgbXw3heZVNlhEvQEWGIRE7B9DOgvxRfl8JCXt+0LYs9DPA9+ku2XVo4NO
Bj8bs7lovtK3E7uC0FGsvhXsL/XG0yux75qTv1vPONcktX31jdnidsU13hJ6DO2aEhAgiMWz7SN9
8UwlRXWpv/S6rIbIRlm4XWoA0gbt2yljQ6B+LDhPr/cB8nhAqYR89hma5OoL7EBIHvwKCQrx199O
Vtd+bzJIaCSeVt+12KvgcG44Efs+HRuvRdQC5CBMwV5fMCdJPFybb4R4PPpvty5YgNTa1efa4HiB
VaKSc98v9q3OcPpaiKuOqzEWVy+o1M11aR9lzEbhnf46sz7WrR+yl6QMBPj6BApPg1GmJ4sFnP4v
DE7Ojyp8LL5MAF9v5oSrzyEwN4J0wML5Boq1SN2P81J3cPmgGLPH+cVbBejJbzxMqt46dHbM1v7+
LjKjjtljVcR1lOfdMq+vVLiaQWFn16jcsStIQQW4FGjKw6BJ6W6BC7lTE59LE2oLJzcWqLNnphZL
6k08QBSTdnhbrIAuf6yahNXLdDCGwFRJXgfGFG6EQnEJXex7Rl9m5kQE6Z3F6GeWtLed/gjEyMS3
FJ0ZtptsAIRneuAWt2VfudJHTE8YqGLnmgajdkcu2i4Dsp8mvfus9H/Xiqef/vEkvzhlQJu6qghY
Ogd+z6If3aa6vb/YwX9BFDHEkui/YvM0vKHxgCD7cLtD1jHqXjhPIzIqJlgcpF1bx3aXSwNzyMTG
ut1zhhcCl2u44fUNJF7ClTEB63Fe73j8FNnibeDp/tOubQgzNIDITOyGo54nirC72aDvSFd9pULH
Kr8iuk8q7zsp1HjbsamO2br2cnBT5z4nwjRbzNKaIaKSLiaWRMAqmJwDsEdcsZ4wM5yMk6ORUEd9
NTmC7pzBqh4xmaHsx5EFoYTXIORxuw8kxNF2mhPA2MAogbUX/gUUEIwI8raaO8lxNMWRxB+rXqa9
HstDJV6E+EusxvYBqgiVROgF8WxPYbLxpzhRZu1idHk+u0IFQuHoLyRB7TmfkPTcvFgcO1pAwzXW
sbpTkLSmwgRMdeq/sBbFNqnFWWCr2szsizLYjpJMrOZTTVA/N3G5O//QODaelLA8BlfYsjwxPlyz
hfM2Q2ppPqqPceEOgA9vbtfEp2oBvl4vnpL2bIcjNLkAHcmYn3xN5Dor3OMjEga8Dje5DQjXOFNP
FbWo80FhShCyAJxDrpxuUaNQjjSahEw3n/tJOV2WJ0tDsmYP+emAsHnGnPc+aI5uWePZd7qC1qtL
Fi5LDsNqJbOUpflerExDwD6MTFch+6s+ySoBus07E6KkYaMPkTJJhda/stDeGE5coz8nPmT7+nss
ptjD2q7GsUxBqZgt/+DcFcsnqdjcv7+kIV47cSa+NkFjk93SsjNp20en+7nHM6fE9OOMe9XQczki
DhHy1ifmz7wWJbNpolVtlIC9aNAhgf0pY1+wWQ9x9d9052ZBXql5MewYRp/iVh/jYATuYOcxXbxB
7t0bn7wG2hb/W9G3SIVoaoBSc5WUZ28XUovLh2Qre5oYH+ZBtEG5qNZprF3kRVUgB1RPiAzZnfAs
rfDGVQsGPr4NDHAeoYB6GRR8IWvOxr/yJbOztYpT0wXoXVVE9XgG3VgGkkizNcl8Meoyazll38NF
CN3EUwPjlvL06IjutfPMhheF0A4D8BWvPqep4kZz2WMlJvQdjZVWvL5MNvJwNJKcKTjzlJ2KwD69
J+aKziCpphrfvePCpWrduK+6FkDaJBEsyg7RwRuyP85G1i4KrEfWiEHEUR9GA0NPSIUZtT5dJ6X/
Kf/4wUnFAOmOba0KHYhkAniwrOPh4CiRZYyyWoAMkVNxd7p8R7R4HyD7WYbmReCh6LzygPGrISky
z3BHPa7/qQZncc2ZaNyqrJO0ICoKadYX0mEokR1h9iPVMaT4FbsoPDY1xqzRnU7bfvBJUDIG+4Az
DtgsegGnsmAXimnhFzYxnICqKEuMU4dk2OAmD0JLhrkf+2a0s+6LAc9Lkq+F32cD3IQLCHJFZorK
GdXQnONTuXH0axo1Aa3urtyuxGDbJTfSwUuRagBH9Tnd8UHXY5gkxmyaSOoSFrhLah+nLbYBKYqJ
R+wRynh+4iLqrHyI3CIH0Xz+NlD3fZAZaWDwSzCBFxjuCqLC9gWVDEoFwulSiLv7djwr5netX8qo
63CYyiief8ApX2zAXb/UNpgBj5kDwoqxAqIfNZqrNz4uTK5UQ3I90yc+6JU99t+Tj8Tc+Ychj+uN
ML+ujTD2RI0emSy16f9siVDuJ1ytBCIWkon21aaikiVFWgRucilEnB4Myk3hNpoC/dJOK7uENu4V
0lDLb3YG4z3RrIGoAf4sLh8lwvC2jWQ1R1+9RYmG5ALmnc6MH73/5M1YeXtOqn7hRyuoG1YsKrfF
UuVB+NosM6DInym1Og+Nfbx9Ipij0YskU1CgVKMQGbL4khkTfyoT/aYSvYOVmuba1f29AQh5tbUg
CoeYRN7g+fPvdLbyfTBe/xRo2OrBMqzeWFiYiO4TBFVAztCRxE64Xvd33On31OkZgcCxBM0cmzq6
QdksT75AyF+A1rH6A9EUKHqREUOoCQbAzI1VThNrhc/npBbdpENOIQ+fkysF/Pg2hGE79+2fGxzv
xiqgQHoexJ6sZLp0e1y2BgnYvdbcFMegfJdbh8o8zl4Pax2CN93DWHoxyBeOfuWAMc1uJildZzYJ
jSVJAQ/GpnQIKprwCs17Xvkzm7MKWlIhm3223AM3oDSxPreUYJBPOfsfBwxE9akyi31Fu84uksR9
xfBCFbMHUOvG8EaguVqkL7EgDylAg7JVcodSmfJ+e5NMvG9c5Drhm/xDH3pVUpC1hJZ9loXEuxHh
+eP60aIAok+uflZdByPtJZMaGNiol7/NJcxaF6f130zS0uLluR6MC/3bCwxkA+LJhjOBr49yJf31
osHg85QySHgGqu3uYyMJqDepbgI9L8Rc8WzOEp0q2MIjw6Zx3RIVU0J8APjmaC9wps/DavfPonHb
GpdDyTgBnvvZzyWekHKZ/4PweGCASuWc6b0j6ykkkQGKpjAbHpi5aeBQ4nmIr5/n+ENupJIgcO0V
XY8z7yY/X/u0+/KAsh/fgQ0H/ljqq/rzQsyYIw4ZN9Xc9KiQZz0xu2PiElgQUpxxWQO5+fB2nEuX
xnehHf673jdvBEd92TtHpTZvQUCmjZSlVRFi4zQrlgJSmLS9rTlIjpGgbTSvh0g9eziGi/Jf4bXS
VR47yS0oWqxRmC9gKSt1sdqp02k6Pc+jzK+1WqC0f2sQU+tYH5d3btvbCeaSbVyiC+5CWRD3Ug5K
EENsYw5fV7aXwc8AHOSLqfH83UP1ynGdtm40m2E3R8rwklBuWhlWmNljrviDvs+UyrTCxv9wpGSB
kRXJebiRB6P71n90fe0m+ARwz+WRY962QlAHyJ3sgYU/e6cRgVY/9SUNQcUp1iAfTtP8/JmfpjFk
6MvAWrDi8fKMQTyDdPbFeApfUn68kzrbfQP2eS+RYXtMbI/Hq18UAhn0c2HR2rb2jzJY3ek5ipar
Cb25B9muZWySJNVhy68yFgq7BRV7RpzRo8sJdW4t+arC3MoPzNWZuFCFFo7sfxFpjY+pC7M9p8hU
WMzpVQ+k+e9yzq15lB+BZ9rNG2OWW7rxqpyOZ7ZPqUC+o+pakN50clL3JZZ87p1F4oY9kp8GhjTb
5b9p+7hPKIUdFl3/mvY8AuFcpMM3d/rtNUs7ZQDGNnEYvRM7xXQvorpz9f6y52ggnMhj5akoW1Pa
2dlJW/5OxRBziw+CTR13+Ax9BRTnC9l545k8i/blZNkOzA0hpvLpx5i+XQrmP+bCS+p8YtvFF004
muLdjFDbMNu0favWsaVA2HpKsXreVYKwieczQM/JVPnG9x6w1QCek1nw1AupJgjOJdSLJSMhCjmC
9aJXMfc9rlbs5rbkxcTOFr5DOeYUROrM/QRn97d9s+bPsuFb2pKrEErPU4pgRKCRN1vj7fyYRQqt
vomqFLTzAdyoln2ZFnyRFYJDbLddyJfCr9E/xwWqpJS5xmo3QLebM5ie21pouv7eyTNvxWmarB/P
J+Lz46qP2Ia+zwizKAAZkxUMngnwe6+NmS1+Bx5/uBSnCXuvUkXL0kOc+/jOS4C1LPLHr13/Me3P
7/xFcJFlpRuBGMDfm1FL24uW0wJWsAMHdeO7a7VJiYEXuQ/BO/G28chcJ/6FZWb6McLVHNWKOntc
PbFTnfTukZOVfyD7hJe9FbIfhDQ96VyW1bi4IHVijzZl45jAX2Yq//4qLVd2+8gkZwKhhhNB/7uL
t2Gw7EUEfuTmqmBNCtHhJeYpSZZelW998BuHNPlMe8u6AP7oIFLpBZ4tb28Kq5OOvHf0hdEVVHRP
VZsPwTEsHMVBxA+TJNl9n1WXraxAFMUzi0BFqK1lk1Q4Fu0bCrGP8/4jzKnE8SwXuQn6agMlKXB+
oAsw9h3NbvCJxix4qVuicR/xog90JHAacgtqQUmbBfZGk1K9m7gnOFp8I9a3YfXlzkzpGYOe+5Cj
tGqXxgplKlkXj12hfzn9JYcMiux1i1cr8/DX3Z3NN9PgbjgggzIClZYEoxUoeWP5i7/S7zcCvOpN
BwuaVAmYQj+SpUsWZE8OQHpFv3iTMlF3+u1Z2/3oS15w4CWLOMCL6OZ2JkJWkpL50PPvWUWsibXe
cvXbZX1QLBnmRSB/smbGJcIQ5wSrrmX+mjw+q/7ojgNskLflKN+EkPYgVMvWhupNVlzSF7n7HVxj
tx4NGJZ4bPOKo3bfrQvZHG14viy0uvwpoW6H6h1ygG5vdutZgFGoPYs/G7/yskVpXBfDKz1VqzfJ
tA7wGvAvPFQ96jp7SJr1CFQOah+kGsahPey8NIQ0CMsOKr/lvNyEZ6DFwYzJzASQDzkBMYLnDUpu
ykT2sDIIIvONpeTXKuz0qj5PJXe4zNbjMVqrWq1aLq7JFBTeHkU/jrL9+9hvXm+70vaTk4HUwOXY
DFidvYm6tbD2myjAWNOuZKzHDIg/mldCXlirjfzcilPO9a4DmlGAB614TEiiEddZ6WZyTjJlSZvE
/d5t6tRsu1kbRE4RhLUxNPGH/pc8DMOUKk23fr2TpdVzKwKVnOBEUSOI16I3dtAoRrAPYor95GKK
m3alNgRj++IfDn7m1rucF7pKMZ170HYGUqHsYMUeoUYu/Lrs1BVWCobLk0xxOzOgQF3/SyeC1BuL
EQoqwEWRd6H0TGrBANXzSGhVkOA3I0DTvBdxGvDLoSmFMlUe0L27Qx5Sml94YqHOYo0RVX6KGzb1
YwibYcKC5XMew6b2ZngIexhSv9U0sA4IRqEe649YQSwyUL4RdLGcWqxMYdsKpIg9p1SW3CuVVOuG
/IGIuRL2cDQcgmI2iz4R6ni7HyajxZIuJ7M+Jvg7wa8HU973ewWrDckgA4EGNfSlUczc3R/aT99R
uUM0pwwsTQUQeIJyQBnZIcKER47uOxduANU7ohIjkIt6J/HXOeGpbiNCefOpEwgTvNX6igHo5sfE
htAETXcorzYyg4DBjxkXUeDNmwjj99qOBqhMZ/BsDYzd5bfQwi6m9R+48Sl9oovkxHm96P0475zf
uTGhFpUruytD9QnFsgMklcW/elfVK7aBu4+gZevjSasVSmC1qSIBKQgNqLTVTptLM6MH5QghQQu3
pYZlJhuKjtRT3sfdrNNxUIGYGqN0BsKO1B83Fnu5lpjv8Q/wjFVIzyLb68enAKNJsrH9MhHEdZvY
bERBvQBF4xSErR6w8Ab8XKJm0k9YimdyEgpLpDP+7yde/esRSeHbv5qTHYKopoeG6ILAqu6Gf6oO
KVK2DU2NFcMGcjP7J5OcLs70SUrnQgWmmUqjPrCQcGMn7ycBHh9KO8KNZ8wIhKhIvJoTFRRhCeRj
BzjI0CIYqNwhxT1nK/8/WaTrb5M1FvUaFk/L4tFz6rhpvDIB5ZjHjjKf6sNKXbe1S9vaunVn5+2Q
BxvG3vnOobQkWkHW/RwjkQkSVjmbBLyUvxJOaPHd4BulMvBpIpaHlrWrFNBSDBIcOT3khO1H5qUp
q5Y0tVxS/I57lxCUFv+mnJRO/1SnPIuddU5dlnqF2mqXRt3CYDOM0+EIa5a5nlDEsqqnGylFQv/o
j1MYkf6Alvvoc2/D4wy6VExeddtCi5qyI5Lh7AQCuXIRFVaxpUdPYrAjkYpIOZ7yhbOabtgO3xzr
w5bp60IR9YL9IOzZ/rLs24vixWDAidTo4egkB4n+dLv/uo9rgfCJmgitwD+sNnRsaWO0Hfcj4dfT
7W0QXNEcSUOAYlF37IKo7EQJgtVstOcrw9OUpy/9MBeicjcTb4IUYuw4mWgZjrD1qmw+ULmP2jEN
j04IDtpGPkUzFUH8qkk0k1skzGRb6182XEXgEgaPbs9KFcb35bMvVHSMmCb/H5Wjy/O7SaeRjrHq
hZMvqFXnNU/wxAEcnNjJvWJ96M5SRZSrzrFJhaso5Rlin39Y4kAJLHZTPU9wwb0vNZsiPRkcKr2t
bcaU8eTuIrdZvf0kNZlIEkyG5dwQiuSMpi+0UFz6XX1IM4VhDDPE1BsLjTcMn5D/233viIvqbJAF
HNKAOj5sgygK5keib6tmaPxUrdbSrKsgZpg869k1w8Ietxilw0f0TTsjFz6ueFXpSq8uXjOM2TD5
oCn/dmC5G+9Qc8e4CDqMJTNcTI1Yr+EOICuagvldAvnNd4QX0GUaqH7mn1N821hMK9S77pbdMIIn
5t7bNqNiGdV6xTahUOMJKYCcH7EvtNUvF3g479zXxJHnC/VEB0wv632gdeQfL7HLLphkWY60xfyV
qPgnckg5zKmhPMlqbsYY77ltBNOBf5rJTmebcffKmfzLBR2cMGbOKPNfjFkcft5Rnv6Zge6FlUJ4
FV10f3RXCOKr+gqYx81AtvOqe1AgpEkDNanSohIbik3Q/1K/eFWbrbz9zHi68VayzbsoXuToyg6G
5L0Pg9hs175X3CyI7vkaIYMukx5Uk79xFB/+R3TqVRCSjT5AYipeonv6gNmUKdXU/whtau50DGKK
kChRHu5doMFnM1/CFW02FCxrqe2Hz4mbVoCy+1p3hCG598UdEkHGob/xS6OLqZ9qqReZX+/U9DC/
wdLcj9MP/Ce6c50Yhc1Upwa5uIkN2KeEmSmQCG5eeTJn9O9SGci7uwZYI+nKmVG/MMIV2wh+X+9g
VsIBM9S9FY5OO1lCg68zjtyIFYqvrhWJ4WXhKpJFBaHDQIR+h7/S7aKMMQHdPbuaSAxTDkgsJuaf
+6KDBFGJHZA6iK52AVo2EMknUNNwsMF3Rj6NpIHgp2A2zWxHulEfCMEVJiZjeZz8KiyVVXmoG6Fs
vASziD8qvnjxl3tfv6FViVJZqmi2of8gfscFUp0XNP9zf919vwsTpbih2Y6eIPp2rOvvTZ/p7qXE
eavbkOsKNiowqyFBG7On+JbVx+Pt413Quo5wkYrmKju5kxA6N2DiS4ie4prGH+Cs0JWhVnBe3ybj
dfq7bSLOGcfd5Za2XQh1rJZPavJJZYuBnpHjqKe4+9ouC65kv2Cp8Bfuhle1mgIqaGJUaUKVJ21k
4EyNufbsVr7emDwM80jt3wyReCX6/N0DBDBpaOs5PSuEql6b92xsMwKbqrQHVHxVPWH5tBfpQB4m
meDeNK2/6WQl2caL/7vXRkGZhFRyIU8uHZiRhF6gAxeWCs0yovnjZUuP3TFUkx+9wqJCXncK6yjB
y2vk0nwpAxgKxg/nqsxv+Oh9hOe90y4FdC/1c2/q4YLRdxck+L9DdwmKAr1+Bpz4//zvrw7Qfq6w
Yyu5zVklQhmJuBOHj2oz2wxLNKIQqc+g9VDV/Ytv6ClCW0yr5ezIIy+YgG2seXCcL/YJu0YqN2QJ
04ebZ0WqU0NQpqxa8ITCf5T2VbqBccT5JeaSqsasEtj3lCHRNZ4/IELeuPYTNsV+rur0CucUKrSW
Vuwnu/a7oB9cdP4Lxo6vUJSpty5qjwrp9yUkRUNfNoWHchnPmsxfLIJ9RWUg2gVeQknPuBFs6caM
1GyOaaw750V1/MekQ8F07vRSkAx/2aD457bx67EtDNZuuuam6j3fq/3k9KNKeQ0SJ4mmu6q3JkkW
ZpYcHLoIKyajN6pRJ31/6y7J0w/UArE5yrHJQCnhJgTSNpiqNpAEi4ctYgVjvXuayDNoZ8FibvXP
tmdTjbCXITBW7sS3sgZM1BuCBK/Cqv4WZ8G/RAiE6jQYaqA2ATEt9IZP7Pqz35h73eXluGRXt4P9
pDK0xKpvXwfKzqoIf2r1a6uYZrc34A0ejyJcyqC7cvgM46BkAEjFqhzN93VbRGkpCP1vG76t133c
Ack8JWt+cZp4IHgBHku8lLXj8+CquZsB16TpIlyusUs4IpqUAB/6HkUC2Zr4oPqhHswJkFY3Idex
e88ySQYsKhgwMXAOZg1R9P6e5OPW0wfY1zUStvvDBqIkZLP+JPETt9bvpoKGrF/n+Z3siIqwtXdJ
etpoxpjQM2C6oBTSKugy8UkHretIW2IalfzdqCvTmC/57B4ylDWoDwa8WIkoIvIYc+lZc7xizOI6
W9sfisA3YNxyw78ZpBUr35oW5UDsZiwdJIEo3JJ3ySf2bbxqOvd18GBu/9zAoRsmvO9iSNmq6w4m
pI8cviw7t+g+RokQ4bQTz/MVSwbYu6s+hcJY6uVpQ+kOf6RgSMvdJHHFhS26H1oM63f7WWGUmKst
yJdIITtsm/DGXR4hLxcF003nibNi3Gz3OF2CEUrV1f66widiwKm4QeLleCeTA7Q0ysZwrXqhUMWZ
jetTEXba8d5O3679D5J7xZK4z8igMhKPTU/Db53U5DTSyyZiOEIsksdC/qXxj3oyuDH0N+NRf6Iu
c2pBEhKNbf3INeWKJeNbrGOfFY50HMA5Fgkflung2Wt1ya94wIw0lU0mpYigSBfMNZaBcXskPm/r
xliQohQmbaJIMyoMYy8CwwFxD+3dX1Xd6HjP62PB5uEwSoRBxGOo74S76tWu5m0YiBrUsTKsmCfb
ELE2j/4SCAmp8frzeObjtUrfKSpaqip0+pDQLr+lwqkPKxZeUt4KfJd9QImx4GJEccs1912+tjw7
WmogeTZTeDchGGw5X1AwPuiDqdlBcstXk1vJ0XRxCmzSHc0FSPRrlANXAbBJcT6Epcg0/OGdy996
lYfE7rJ2hdGWySMCMs6w9+CKIUgl6ixSMXu7FLEHtw5LkXpiE1e0mvOC2H0A8E4LO28bVHcEnIZO
jTYS3EY+TWxemqEQtCWsE8CEUy/21bxnBlHH339OImpBzwQ+ol2XDum18bjVNBRBLNIBwmZYAb5b
9QScrwsPqp+AL0aOwrjxG/iChlbeTJLLo5Lix/tGebCB/DsNjx0TIFRk5iU2kjLEBxDTYReBr0n+
O3RhNWpsxrJEHnyHvB/lRvfGkgLOEYrHuDo/35sjp91RLn6pCKoV5zL2/8jkVVtwwg8GPEIpXDT3
fa+baFAhNaxz0VjA+2ntKduhEGazKvp9V9/uKLcvUejG7iw6RF7bzO2W7gv+aCCefRuAGgFxEuUE
VqsX8uqVKnbL5OjXz6pTq85/jP19dVb4J6T4pfLaWtCmvFrwBnb1An1iSHQeNVDqqU++KDhbZQ9m
e7lVIzPUa5uSqI/QxcbV1+jqH+CZDCo390rhOoRwSKoqKluL5U96rsRQjip5iYwcGalSlFoSkJd8
016gshWJrluB4TlS/sHuFFYs76yVVFFLusjagb0E96XBQ6QB5pnkeVP+NqChXVu6XPoIChKY7N2R
s/OezxJ2IL4qgJ9Vewj3JcG8f8lSqdanWM5NH5QXP65e59jYc2RTPwkB5wUSjgDILFwT3+7tWoML
7BeRwUNA5OwafJf0H41Slm/YD1Igkb69wiEhCU/ryzKJiswylShB34zKNWDdYH1gtI0U9ijn7/Ix
+DOtFDULOETXHn9rMTLeqsgXIiaIuz4W40x2KTjMGzGnWqFE/ebTYyuWSUIj6bZZyrbjSRyabNYk
Zjta57Xg70htDrzB2ijaulctfdrXWJ6jcgyofxat9zZvHc/ybCLHkpRhH+qXf3RUEWMXGRKoRVSp
0G8IeDJWynzDD8da9a8Gw1N6Tt1I3xdoanhIr+l3Vwvk++sdQmDEPiu48Kj1V3eDK89SREKyP90T
bu4Zs+JRX/ryK1fozd0oEdHBCiRjJ/ixGL6xe/u9idAqJBibjzW5P8gHLTX8PwQF4+yLUeHWA6aX
3cKsD5i7jGVgl9WnTa3cty/Ak825RV/nC6m2uuWPJNzVM+NJoVY04nX+GkAYHapypRM0tdEOpdsL
l40w0rKGNLREvDfcJuaK8unB9JZ0wkRhm7KdjaONhEgZsvNVIPpSiamblQyZL1TquxWbdEbi4F4+
MbdNwivruoll1NtWelCrd9Q/1obxrZJO7elkzPNEoY0iFDGVB1bEnyi/d8n4D4sfyxt+oC+FPLc0
PSNJOTFRnTrcZgGWiyRwbrK0ggwLYY+AXpiVhFwXR7l7JyMWZX2bVZQw7wEBwSaaZtcPdUma1DrR
2aHqJf2MwrWRG9ZtwUtuaxiybqfJa7BM18bloVsQN7Vk0gWLXb/5xM2J4gdXXM6Mow1ldDuA7rkh
Vm+XktUPaF2CZZaU+/uI5hrppCxi5yHgaJ1t4sCA9ekgJf/rPgOQPZjUYhT2iTTVww6g+jj7HuNo
4PJvLfqnJ1TS9Pjx7wvp2j1VP8K3vcnPMRX97mxk3Xie/wLrwdJcJY7M3BE5F/pK3Xb6698nodxB
WeVtLn8TuosLnC9A3Rbxql6ol+rm2dkZKVMTy4xyAjBWTOuxw7rBeuN+FA4ki67djZXro8NreRDm
G3kV9zlPujYKK7u6/Xatuj1ZQG4h9qsF+nQ25ZKFiDLEq1nnTsE1nmh9mAHd7g4oSHRKMRtqXUWA
L4prUovLGjXdN8o0kEiOm2yJLkbib6zOUmZWOd0Hx/fpZ31vahtpg0yUJcK+gX/oCKBzBzThBieU
YEAAdJ9TKxm3EUDNecfBWe7/3H/+cfIR7Ko2PFQT6TEYUNbTIADjG9ljt6ixGP3rPrdP+nCJLGQ+
KMatwasln9QcNmGmPzIubwGf/6lIIxHr4YVjYNrmYCeYz1G0P54ctaGfbxot1psmwo2+nbS9B4JR
NQPrN0MbhEH6bjUM3cnGWU/MKLoyxxkqCpEQ4lOnUdpPhE26YLhtvZhtrWe2+mXlSzzyTKOadlv3
jvfrrX04DYHNXbtX1tvL7u4dG9jU47hjXBQaMKcbeWH4xKXwx0O759If0lo3jyUatl6SzWOOFWJw
vkt3uy9DfLjZEtD2JlWn0ir75m4vmCs+VS4+3+tngHAaVGog2s3BNrPW4eL3nhIJhwf+gshz8Knd
ad5seYevyh/HT0bY+dYI7ZYT/DuKOTTuzEuqal+HB/XqfXAotUfF8Sm4QJJwZ5rQjEdDJKVZxn5y
ynvRW1JVA3gsya8IcYsN/JcFJCWvYFxcNtVAfVR5IiQngagSpV8npKHfO9MG1aWxLEm3zo2vMUUB
1vofchAhVU7dMOm+EGEIkUsbSX1x7r9R3Be5mXJ5IC1VtbmyxaPA3GPzyC+G+WYTigwpjqnajbmO
i4QHQna76Oc+PcGcfAu6h1a0JcGDUht22ySVHWmdbF3GiFmAGMhyqotdrfbqHLvanYt9WML1T+/Y
crKDVMW/6wjpsMptOaGfZ2IlN/fu0h88ls4NfHMpH5qvBqZJe/Aoi73F1pifffw6UQpECQgOnvBe
L4j5Q8Z2ROV3BWfyjgDN+z6Z5iFkwEj8//U/MONs4zOrHA8OcoDwR72LKw6NKDDq6zbtiNrq7oKh
L1eoJ4j2MvRkcDMb1mCDoI7K8yfiaHOGBtXBIffgkiMi0Qx6O9XRGwFm0KRHYWvC/Z8FAZSL/HPN
Cl7eCcpkXSoOSihEQM3GcwNsrpeO/ywENnX5NTaLkzGpH5odyxWp+Y9/ieUlQNH76dV+FzqM2Bod
gm5I9YxEW7oku1w3ZTwuTCMkqLeNP0Fp/ZgOL7gvcfkRs6uxTEiqEItlvdjRE6UYgeDa+Ew/bpsY
Vic4o48sfs62oT18NAB4Quh7KD96EX2ZOz4zcoDDpLy2cQA97WhIqOEwzlrvHBy5FzOSX8/VAmRk
yuzrtunZaDXin48XZZh0jBEna3J5Avs0TdtIN2rORY11pQRQc7u0rNlaazM9CJkVSWxXdo4eIjc9
I3N2mYzSEzgSEua2tflUl5rb1vbfEaAPOF3xhmeZs+BkqL7H+KPBDNBOXXn5cHbXet+zR5B+c+N2
M//U8/0IDxhm+FLodZ+cpMY9ufR/wXoG84yvcwNtrZqhFcswqndNVlxAcc1PL9DwfIX8uvo/ZDD2
4VXyIoVyaFweWz0PzsTzzhoCW2sAguVg7Fvj4NnMj5LMJxCu80EkSy+3jAmCzzH0uUZF2haxwSgh
40Vcws/yRjo5Kn3IQA/K7AK+sRnVGrJxdDCgR40kxsMnN51/D5EjEpt0FDrzKCJgd+THl2rInFpi
fAD4Af5dVnVoiZYNE25cnrwDaE/8q0SJvCyVSDO+ivncptan5N6ruV77nRkqZENuQNj99BVo/bwB
hwQZe7uHhq0P2vOuS2zg6Yr01d64raAH8HLFzVtoSkwKxrtMLyt9/onOhAX8labIB2Sprk7LBQem
SlplmyCFGSxtbBc4AT/+wtm7IzhsFybKNTiV04fz60h/Xd1OvgpGJ5tIFckb0wF54DUUsTqBM/Az
7oqj54Bgqk5ikEjqiQiBEEHmzH8+JplvTfEiMHi7KpqsXzYL6imtQ8FcV5czDgV4kMSpeZiSroWF
J8CoXJUlsYgxfPTQRgjx2QpTHsRND2Xif6wz8vT8MbBkw2hXl3v1WCA40v6Vm8zlAWgabMBPmWV1
N4UZIummFoWu5dS3CfqGxC0KAsjkg9K7Pv25fWux0snLskK1ztXFeT0o/DHDYVB7GAdpocSGMjzf
4lHG228QyHtf+9nPfVlabopOVso0ru9jx1Co5H5zaMmIpsSlQAlFpO9yKCvb6LCGgKw1W6vmqE3+
PmhA9vctm7sLI7xnj72IO5hMJzDjUUlL4z9mrFzYoj3lePvqPOA8QpGJuiJcZj4V+9YTT3f9gmHI
kMsZoeO54Qe6ntJZ5RtAWO14KNoVtdBjwYBvyLibFr0QSwyTCve33AU5B6840cQN5OjCPVQWAPDW
njrY+Hgq2UKNAQ4vCjHywcdbnrXGgQm2kzqtLbuVTIprcJeTonraiFwlQaB8WCWwMstvcq85xOBI
U78zNR6IoGP2fkJsuZSTa1skrdC7lx6PQmq36CgwNJuJRKI2mEbKwXT6ss7p0MFSCdC1cgF/CaPq
SEAxeWL8SQjvfv2AXyagcI7Nlq/7PEFqWMf2AI3J8l+K7oMV/2/gCbGmE5d5WlrE+td+C5x+eo7w
XaryZOU+RdWxUc7uF2TZ1eGU4qE52bWWyk6A68hnB+dygxZjMJAXUO/Jdj1vhl4P28P0d2XCRjGe
eZjpj5YAZMEQPsRKu2ddiAm+IbCusm74zKkbUCQzI+Rl7WXBnvznxzqFKBoMx7Ch1/pxPr15LHUZ
bKT1J7kiOtncGLWh2I1KpgSxzn3J+RrQry+vAOmBL0vS2hFdaJJ4MneazGKR2ljeLAN1WJp+sD3u
I/jmMx5fgVfMUFC4yM6D/vppQHV0BMC1vlSfjLlFMtjYxxm6VfrUgJjUqyDlji45KfDpAr77OOtT
lmFlBtUrxsbM4TJy+d4h7jzeU1fc4v6J2kOJciezEEHGPlK92eMc8nyRr/22PwR8s7Xex4ae+uQH
7cdauXc4ZI5EmJUGaHT7SlHKIP1b67DM+BjQvOfJJqAW5vvmK+DcMGfj4jvw9fTNaXi6NEBUcMu2
dFLQ1V3vzxdth69CGMMXbKt+gyD6z/qMZYCObc8wdhygm/1hpRpCMmlS/a6hnhEt81FwM7CdeXjq
uBKGOKdRP2LLRjkVM/y1h+vNmAq+yBxsiEcYu4WY9E5iNJHFW1AEtuVOEaQAhtoG7/xOEQl/TTWO
4w51S6DfxwGsKxvDkmFawAWDaeO9S9Vb9p5VUgWpq3Z8upvvbTXy5aIlyZ73qYBxsfdcxpiIUwkF
OEp/6e6cn1JsEO7ct8TPUwz2I/PS/zMcPj4OrMAa9vkx4IF3x3G258s7qhqledQS9My9XSmBirz8
NdN0FaOXfedwd/7JJBR6QcVhuUPRCGsvL8j9JMkuzViC5lsuD9VfCy2XFtEIhFf4qLrCLYJJO6LV
iBlCNvqgy3J/6W7A+SjjtNBVXILongKgRdtZ2YRsHzdiIpL4K7ylQ211Vg/gbqvEXCbNHpXtj+jY
qwTC4o/KMsQRrZseJn1KZ0Zuz8SKdBN2pgDj0LaRPGxx9TOb+6WqqH5f8muFH33WbboZXfsmCdBF
B5LCVeOvbhGfXpENMkpncUifhL7NVrYKwQe6t1FOzSywk1BUq4+XRiFqL7FU8L3BUld35TegCqbB
neHpyuE/Lc4IKMgG3iDP9liO1nfyPDFbdcDYC1VMJFduoCxm2YuHmSt/T20N+QaXiFOpHP/jOapp
lQa5jJiDn+SFcOZrZ3cffvW0LDX1YTyD6L7HRaUR4jFcfG6gkXUicWnylJqEzfcVhreCW2dF1MfD
eurs9sh5MbJROW6Bt0ZSb5F0UGwrXidU2keBNejy4fwEwr18lAt9REjyksPlAJvV2FG4w/l5mzRZ
PyM+ipda4BU5lxfZX4aCYFHJZBP0FslQa4P+nqGdOxKs3kfpbhWufLfe8nLFF34pkW20SMreM3Pa
DH9Xsoh1+DifIzWXaiqpmg3gWHoKvxi4qKGBV0nGh0eNp0gv/OwNsVuUySCOBO3wQOdoViv9lrmA
vqvN/CJOUtmRZoHnkKyGSoDfVj0eZ+adRYbV8cF8O3zWyBzAsqm/bSd/Scy0jSSa9/lHgQDyRFri
gVt6e30cEuTj7FVUXb4UN5O6hUqjZ2QT0UgxuRsdJ+cjhMdSKmVSshYQomdDmQhCeCKARxxcY9VD
PFbSq5EYp3B0O/2gn84RLoAhSIPCGWdqHP7f4ROiK0CEkVkLxwL7VPv9N0h7V4kAtSN4A44ApzDa
RCB4bX9Wft1SuTVgTM/Yt00VUl/G6GNObOWJqCNlNrXL2neRDBFI7boezxJa3Zv6zm/xkpr9BTxU
pVAsc/BHtVGC/0Gn7EYVPj6JEpv7IbSrP/TyyM+xII/pCtn00QtUiebgj7vpBWzx54X9KSdH24J0
2Hydfb6wp+6U31+h4j8UWTAkgEWXwbyJOA/Ciy8vBfzILRiEDKfELi3mjLAize5b/zhRYPnKpuo8
wdzBaeZNcpsHrKqnDRcq2AEHynNupBkqPzO5Bzqdah0ZccZFpDXU1RlJnbzIqEI3aI6aR3gQB1iH
9rC7wxqCh3e1OgOmp+QOYlimb5O6d1pFVXEnqnmkji1B5nppBZcnABJ/6NgCvAsZYca61ADGsg6W
ADNdQbrLJL68rZJ9Eh5t1zuaOQe4YMlsu/QiBZrxzec0kyfkV+nOEGzmloRt/+BvG8R5hX5jZjV4
hswJhmcptj76H3HRrBJz5tm6i7tCz/u8Pco3xLtwvLeC4WFOzFhP9bCeETTt3hQhJeu/aSqDBlOF
qwAZqpY7ed7XDMfpJ53Nq3IHFIMmgKLNM0YDKiZlXVSCrsYoSsw/I/YLnJYWf18o9j0uW+AV007K
+yqu7guNrCLt738LJwnF2K3W0Az6b1HYjTTd01tqiXqT2Hr/FvNE8u4/I3GqcCfnZi2pWhBXqqzP
38vLNAbpaoWYhV0UVqeiQ5I6ide+z2dfs0pAq/XQaRy6bcnQHstlp8S7aOJKHYhMWHNb413uqoS+
gwSC5c9Iah+Of+FJTsBNMH28Oy3wHedHjeStsoUbdN3Y5CwS5S0aVU+zDHxL6vEsYayTXXUVYIuu
hVByUDAjgvnKc+bsBp+nUsPdVjHP2q79/UgLC1M1BLXO18pKa2GMIANJdw02cWEwyDGic86qC3sQ
UbivXvOqYdV6gXLlDYd/CQD1y5KfAFQwovJud0OWhB9oFb/idp4M2L0E6CbkBk38i9Wth/s5g5Nd
pNWRBcdymH5QlBG4RtQfDjnJqget0FMB/OhfhK5Om3m41XuP4qgOl+CXfp09JIiZRHq6OWRg4WHf
YkVN+uQ09JovVMWUS8wxvwbAfoeCfa0UpZs9P36Hgpyp+95CX/ys+Z81o3vVoV9Ik9adsCXgd4r9
I9b+OA3vmf6cTcq6KECDCHfRUoj165mTI0fiJ19cb4xl3A7ECuS0Ay8NXRt89ewk8SS1lhjTW1+Z
3NPiHIUQ7zwSmsc9z1K9ivg+hiLrfSRyJtVsjnFGtpjFYyMbU+1u+FBYHxHieqBSv2DccqftFZxO
r8QMYFK8qHm0Pr7JeAvUXGk7mVP1DDVOJgB6SwQ6pYqrGSlSeeeydS7JyJmxzua+BwVKzWhyLR0r
E070De9e0bYrjyCD/bh+RVETqj3AuJOTHOEZNyklWV+0g2LXfJaYCJnR4bPsd7DKEpIDZn4dSg7g
C9PXnURL6EXuv62Xr6q7LqPUqls0CES6EpadvzfSumE7fOQFjL1YoQDr3OtTl9IEyJEqWse6ZDJ2
EEgxXgLBgFWbDORTUET/SFrfyert5h3iRb0pkR+mXKarVt5aBS+SIOJ3Rt/NDdul45f/mMkOaq09
IEdQTikh50MBipIPQIygmLuv7QBePnD30aIpRcMM/3Vj7AGcLpbNCWYKRZXlTOJ7SbEP8mRFQQCM
5muc1wmee0KErXe2+6bDDjP0GUZTH5mKtdCZv4gvzYNCRPJot4aurZHM6b62J5/5PZr8Mttv6ULR
/SQKceRYVDJ6fKvuO1M5w2K2QzhQaNTGKmZvqjVFKdKPMDkoE6zjk45P2qeeEknwSZpScmPnEO2H
2iNFq8g3TyNHlNKpgDougf/5ql7xmCzyNydfpzN990I8MayHLoc2oFjAs16CEtLGpaOyzKoocran
dw91rm0l9fM8vUb6HetfjZNB8RFPTRd+7Cjmx7JgXEflM+ehBbMOFK6enYqt5+wobB0gwjQh8xDM
WVzJV+OwxsO8lJKwf6uq7W4CKKCR610GXkRB4CF8tHBOVbkWya9q1Zp70gZ5Gx7T/cH80afgCAYb
gCJkMto4AOHPQ6BKFzBFCQaeS1gWxuRYQHcOaZn+oi1ZDGV64d377J7emT7L5yOlNBgcLJo8uNH5
e9n/B+EGMxkvfOr5JIKTh2vS7dbZXQKPgn9n/xTIFnU2JUtpOAqj+K1pZwPZ7gj9uxRj6CsBvSJe
jUwAWllTGh54pkXF6rM2mvAFUrAbSMR7S0pPkonBZXglIbUcYPHgNTx3/m4/9XIEsk2ug1Ry/M29
eHgffBgA80wiQDmw4ycH751Ud99jC/VYQiAJhKcDktIcqbj4ZFzjZw+JFBfhZs/YPt8vSO3FHX/d
ngW1oQLP9VT2cZQcakeLOd/PWwnm/mP2Rwe3rXlh/O0cWmLS95PxUqcrpuwjr4BCvCymVrb7zyQa
NfimfGUxf/kR8vaSubFkv7RLJMu5nrzJMOMSNbx2DLsNofVAdANFnrwlFzrUHO/+8LFWwr0r788d
ZUKrqYoLzZIe6AQotxJU/v15qoEtmRZC/gdFzMyaT/51bITA4SlZn0yogX+FcO1JUfDIR4sDXbSf
fsVKIlLP0Fuoy4GZIB1pUSxvxAvhfsofbgJnidwMzijIx7UdaUT5BbuGko3JDFJzL675n8mFUx5L
mNRBTF9sOiYI7dI06BbNU0yUZgZVJTRxuarD/CgM+8vfUPnQ88yuV6OAnfLv6G3RBwftWXDqNNOj
bQo5fg0cfRSRlO4lEz6rw4VotPP0Ysd3GY77EuM/qT5k188rhBJVcvgVOrZMDrFlXJIaLOcuYj39
EGE+F8Qfy9nYjMZIVrVYhRyrvXIBUzji8mo2abR/OvTQM+K72dJPKzgiYSov4o+BjKuTVyEuheLS
uIhiSmt4EJ8E6dHWWLkmjMwgVqVsx9X0kQIarZWAuyrPWSX8Ak3tm2O641tzh4AxKftoy7HjhF2W
k3zq6Arbl6+rxNV7mAXhgi9Q9zluzY8/TOJVY0a/AstqDCAwOQt0smgblO9D0GKvYuGy+19Z0KTJ
TtA2j7ZTSfTp/6weUgz5CwS6PxBs4JeVF72H6V1N8MhWRwT5r4wPH6q747DOmLQnPflOvPCLUp6N
vaucHdx/CnCh9DsjrWj0BdZAdx0qFtmJFgVlGNLMSA5Y4W95wNPBwe1EQI3BH8JjqyEn1tJwAUpD
jtODc9LiynPWuPJUTPKTn1xXI43tprXytZYmLWc6oc7cbf6YQohkpdgJvZxiktn+OQ049QpPgvnt
+izXArPHjZWCBNH0aOzZRrCOG/iVoDZ7TuDEi+CLv3D96MoYTCTuqCgVlwPhK2Tc9xNGdVWAIlri
qhACW30p8GeJGsjahUTcSyZSNy5UK0bka50cow/s7FxM/rpp+065FfpoXPaUfp9xvwiCCExyoy+f
r9+AbW4RGiJ0/H14lW+X0hag9JBlctcXMLoT1tBL+3Pi3tAu4W/JW7auMCUjGdZssCrh64CrqdfB
wEUJJzHr0v/mdXi1L0iTlEoO0tVbYPE1570pWJjHkSKcVZiOwQWAgwbxzjby/kEYsJzKoHIt9F+u
/bFV3/nF0Col+JX96pYwhed/Xc7ZLTL+D8TG3XKbXjA7zrGdxdW3D93bky4YBn6CnKkcUUcnMW/c
Uxu4nA51VPctLo9i/FjbrP6IhGGloNMqcQdHZf5xODoBEwO8WEXzDGYJffZLPTUsJHjZ5OHnmhef
iY0WkbP8XIHGprynjO06Bo3wbRIEPiRoGruFUDaLgmFA8ct0YO0QNqokQ6526cR+EtE/0tgl789A
f6FgrCTuejqDqtaZvUSmYNL9jnb8wkH0FgM67oGDNt5Hlswuti15t4rxOq4IkcMaj9yu1pYqbkj4
AFd1+fj6/VwguNuBo7RogCUXtxFJKr187ukNOllucAEFZAzPiUWMSkfoq55mVoAw6vtM/8deScT4
XjuhkFlKale4EAMZH867rkOvoERZG+0bynZ32/GG56kxwXjtI51QPx8hlMPj6BqXk0gWUwAquCqs
+s/v2We3LkQ8iLSnKManXRKKk/0iepIgi4tri+qplts0ee3xmufKxbARbf6epEDizuVLPfKw3YC8
g7dfMchMn0WQPYfz+vLYUJl4+caHJlg/wBN+JFD/zFoTaETVGlz556MR1BUpycqThgkeWpgsmitf
7yC4/LDnNQKgAKT+ShhmdJ1DeLTsLGCKwWqyBRnwyZfnhArdkWZrY9g50sq8tBmBw8iCLMolVukS
sBZV9nwdQaZix7qSC8VMhIXplBiaTvtU1lLw1hco8LnAs/8V/I/kHb93wDQtybw8wIkAni9JZzTt
CgCU8VJkyrB2lssp71/3AOkJvUuRWBenJ+pptDA4gpPA322Cn+LppOSxkA+KHpa1rVCTTqUyCCDz
yE9EDDNLqtFYzz6kxXl8gpa4BB2tg1yUVxF/sEp/Zf+w4Q3X4utHd1PP7SK5eXPpiw8CzNbNEbSq
H92ZjInXir1JAgN/cyVqcdiAn8PFKU8SiEpObXJHWuDECeNhxneBlmI2SX4av1VpfGCc/uP2bQ35
XLeS7LhwYXZr/EkvitVY/RHCPM8JB8+dS5zkP0Vbd6qpQqrfDitNkQbhE51i/UQKF8SndL5Dhv9Q
VtSxRpoz2Yy0z/QIq07Adj3mHsZ+Ngk7KhNEXGO0L6r/jP/mhZ6F51jlc5nhd8x6Iq8MUh16Hz7R
WgGU0TaiavftivKH2KtEB5Im34zGDC4rxvsno9c2rV5V5xKzeYxbPUHXNfqNsGsdUVEW9JYxgM1j
/ULgWWwsdlp0KkOlWugs9e65aOM51NXRnYLgAMzgnmEanY1mE/EIam4OL5HDOTC/oex7SrXOfj+s
dB5zJDGOwQ8pqYWB5dFB8UJlwPnQKRErs73M9Y+bK9dVrzJB7WHpYXd9et8mMnZXkzKpiRZTiOTa
bKq73yj2RrC5oZl11LA0Tr+X+MIvIX+wQbECYm3O1tYwf2SgEpacX9LTRVsj4ISByZ3ECYRGtA4X
l7IJYGRg7TinqSJK1gh+bzpEgEnlJDZH4bqUKHOIyBgKBI7uVEGYxoz1rjgoFgQBnmLc4eNmcUGG
B6HFUMZ88+e4ujHh3Qz0tldj6+Qwa54RIkk/4b3RNQhvgJB1MozNk5six8Jc99/0t8worQIU1s5x
ZJ0iwKLD1phnmu/T7ctPnKrjRzXpqi+yVkmPKcJlAUFJpVLSXVsh+k+BjNvFmwUnQbHz/UAp8JFK
StRRefdbU9Js7R7OwRPsoY2gCfsmqN9S1B8E4FBpkV56tB4CUqpYv44Kv/8sj4f2KKrwjTXBEydk
Lmy/RB0pswEi5a9uC0tbZNTLdyhr2+kKxJXOvA3xL/2htRKC4xXJdZ214993y9MVexreTmHysYoR
69J/jKWygHLEMP7DDJu4rt1NG+nRvJr6gYFow8OVU/9gks1YKQrEvNisqDarJWXJptP3Zn+PZu+f
m8zEjYBSf58+AQe7Ce6vdYGvfo4NiMuKeatGQU+vnj6QF/nvg9IPr2c4NJEnPbYAjcfiv7jwZuLM
K7D7StQBSD2CV+oYn5lu1C/x4XU5px8qWzICVfsj8lqmOGMNaRThEt+zrsURIYTsqFhAkePg7Nzk
3iDWwa5mOtyhFTkD7WtWPafhU1bYxZVJD55j/OwmWTTTYrWPoF3f2Tnl5xub3UQyXv/miQfH9eKp
V/Amv8iGBdU4b3PP1tLn7oIXZkj4rT/nO1aMbCk/FbL/+ZbQF4jTy1eEpupy4Pi5acIXV4aUbAXt
VVZN7d32YNU60s7pJQukqK44bX3QXVEm9rAgJDyiRZz6IlSva3dxcJxQQs9lKjyK9Y9Z7bF/8lFX
W7D73+lwwS4Wb2LM3kCSUNq5fY/RjQx00WezB9REpzEy2QFw7G2Muw40U8o4W0r/cVhZujSeYub5
25nLE+XXUbBGicuJS+H1WkoG9gTjKdb+IxHOaT7PnSuMhPSRwlL/rnCMQAYNnxOdZ4bCxDwySZqw
0Px0+X1MYzKUMi3s04xi7dPCuHdMLnSMUAp69+12XycJRSpfDuagaibcIDdXQmIUCQTjR0EglOB4
zOsuLrRf8VuO0XfVHR7hElJ4LuunW5O/t7XXYfdXxARcqEVXeqXiVIi7NX3mNJneP+pM8P/EmoXG
yXHkCRsLwcEcpgzuYuje5cjDkWMs5kAnvzgJDLTgIaU9idtsw2NI3fWV9+ihBV1BrfIB+RyyMjty
ycERNB7t5FYBUEKFYvJ6NF3V8VZtyDxGMYsJStLiK04vjzTI73XgznDnuvjcFdY/A371BY4Pnv1z
x+LAeF3mp8tTVNfmRmeKtJVdakQCeM3Dhb8RWmsXcP8gnUUm8Gg9BIpAq5J9PP0Kt6BRmRE0Vk76
CcPacqbtYXGw7BH6fTnDrGEoG7xRcD+/psfRi9fT70My3wUsXueoePlYeXqoc2MlSpRlFoV5lQKY
aGgbulFVm2//IweQTnlkEd0G0lMvgcR36uogUPPW+uL2dpHv33/YrtI5WScsL6t6s/h8zXIsaLL6
Y/tM7ZRXGokvKSBSP9GqDwhrb1c9r+1dyXuyh4tK2BizMPFtQ0XKrypfSrS1sTjEAgPE2pN7MRJU
WH8s/OVmJy91aEvQWIY6VH3q0Wd4JHSoTWZPba3zzbx+CN1fOauoPqGxpKG05+wQvXCeeSrUsQmw
Rg0cXq2rtFcFLvVYNE6p+85XsQsedAhsXq0gsPn72GvlLNcNvv1KHAm2LGJ2E7NEpHuiWQO2LrNr
L2uYVkQt4+qgE56b0eeqBxpSTIU0CRdIrbwpRrSP+atv6/hCGFEZwEX2S+t0M7ycYBerP/k5mR51
F0WdhhF5pW57/IHHqm9jgpaDmg8XGJwGRQgbG+aLpP14HNg0qhRjOEOQD+UDHJlwToYaFm8GyXzw
pMvuPTo4rLSOmPCHBqPSrK4WjvHhEvKGE/R3nliK1BheLCcPlyGtlP33b+Dasf47nayvmxPoOMHe
WbMwluSTxHVVJPc5XUHc6crEIIW5ia+m1Lp4GC/OGkOGGBi4EFapiBYtsrEhOoBRI9UF0GXYe07J
P+LRGbn2Z5XBp9kr5utJ8+CUWXmK6SG20rcJwZL8v3lgtAqktxxrww1HbjDivjX6llOt3hmBVp7I
5kmLGWdMSc8mBb+wUn3juINpy3QuY/7kKY2br4mAsGeD5NfGeu7ZC/r+0MISVHC4VBqw/L6uiF2Z
sZuPs06dgJ+gqFQeVivD45OwrcHoK3Mgr8oOLNS+dYst85pmjhu3lQ11XE+zZcgthf+zZzSI2CoM
Kn49Dn4MbPBlsRz6lMNLuKMi/gu956L7RnWQ5PoAUy/VASehTSbgkdE/wBn5lUVIZD90p1DY0Evi
pOSWZMCjymjuEISxsNFQBIseTWmiuJBUGMfiQ9NKzeC95J32CC6D4BvoPq5SF66SFt96lWif4jLA
gFh/tr1lC2H6B0/svA9fu+pIr/dzNniZz5vVwJRuz2NGyYOra7epdNhORBAHmdQtuixj4ByNuN9c
d/FNhIcguV8jJeD7pRAjvUZZlQ724KJXb75jRz9LQoV94BWxbmzeElhHYe9qQan2P4/EA6ed2chW
dA9BkCC+8W8xqe5ZKI3pnUrWYKpXr0L5RSZnQ9nwRLaxnCrckW6pImPcE6KAFzjp6ChAgcqPBg89
RGOoWr4f2+NDCVWyb2RPSBzotPHep5dVDq2b2Y6sGC5lznc6yqF48qYO+Z2FtBHWPohCZFda2q2Y
JSxG+L75CxkIN5IcrPs4mQF1am8TMfRaUh+WoS5URv3DUexsuAqeHWMeQ9FPRzOXkhRQVvIg/oDc
RFScuP0RykU0eN6YQaN79Xc77zT86W/3fCe4b6aZljbV1C4YuN3tazD+EFiJoMT2oowRdSLdaD4B
aTf1KEs1pv45P/FFpHqEUH+NV/ziw5ZIY3/beuQB5SHx6M/dvpdK7/4q6Ir3ThOgtpOL9MHZ/zS1
dMEancZKYE+UodhuG4CX7fUTlAmFTxenPEcUOcAjBWIXvdEKOT6I5Wr3etgpGFz+q93WnVZXwStF
vi29sSAm0R2yxEDEb9gt/qde5Hs0Px8tVLmXM4cpx9+9iwEDQTGtZrp0L9NgMGzeJolI9z1FRyMR
N78wX/cVtdMLXLZLXvpSqQ/eASp89rKF4y7hPjduptfkUit8cWYq8wuP3XS7AlsF14z8hR+9ZKBb
eVbungCw9EwatFfUm+sbkxDR+l6uw3pAQCrJCeUx6I879bta47I4ba62NKgQ2NfldceGsf0CcJZs
ovmruhGAcVPUh0soLc3fPY+VWNF42fViR2myRJzPGevaDtGccmOcxSAgkoCSOSG40iOJa32mILFa
JQ/cnEIEvgJbdejEhxMHRzbuFAaOY9NJo82+Z41SVD9kt0LTMSlGU2u9Pr20b1FRrjtDtuobpVpH
2xdQ4c5X8xtH9HjmFvs8hW1wWDZy5s7Wf/vG2CwfBL+tPc5/cHgSOVIuuxTBV1+2DvnGt6cl/gh1
/if/De1anaGe+5M71PKD9t3eMbwYNLmBlyOTftT8WyyK2HgZjprAluc29xfdtUbEJqcPFDDYS7D2
cyJaZYojZf+O7wwkOccrNyU45MCn9S8fbEUrRffY+3kQ3Kkyf+MdMdz7R8AEwDemwK7GL9oFXQLN
r6nDagQNBJA0i8mxhilVk4lS23bb3h7bit87GZE5+Fb+iNQGLqqqme7Uyg34F3BA7N4xTzfy9ON5
PSIFXBOFUne4zX4kL/QNK5odawuPmwFTrjzfU/7POjKXEzkZ9j8tuP8zR1OHp5TouwF0Qc8qdtYw
xpyKP4bYnNk9rAZTgKcYKjvARA1dAuK4OtQ8ZJmGEEwxI5cP5x/dijo6lxQS+tTXHBGVi+eSfLka
u/0eg1jVY+q7GrDRHobCaU2Y0qVWHXgRekWSvyRA+RVuwnwX7Ryk1g1S3wWnlm9atGLgEJrSnM22
MQds5up7DfFwFjfy4Fi1ta193msYP/phnSxketh3dL96GQ5IOOuzBPMhzSqy1nZdGarDF0cynDbW
S4J9vge+p9U/RLMocf3D9DNs/eAjDNpgyMxXbt8cvCjIl+A+60COoUNwYiYrATTMeYmU7anCY4o+
3Pg/sipi5lO5okUv2WOTute4ViIGK75LFQ9WaZ4TJcmJPMbE42gUPge9q7dDrm3scmKB2UCmQX2R
iCu6B0pZ1MsL3opBoC07jInQR9n42LgF9dI8SYaZME0tdTR5DebQ29vo+WPFYyzICkGGJOmb7MaE
izbwOZSy6ZJ2NiJy+d7QahZgHcoIP501Y7zFxDrCYEfwKPWydNoujNiKZi2ZM1FLQ6iaHUm61MtB
ZioqQh1dnbGMbxmtV6t+7LoThQ1M2uN6/csW/yIgreNe1GsmAT85dlyd07keP4plRAp+ui2BvhkS
kI8JeVSl4bJ9TpvLDYRWY6/Z6GgTHtSYnjgzRx7owEvfKdbe08Evzn9bD0IF8FbWcWgm3CiiPX4M
YE04PXZwPK3e21qS+9tu2ETFofZMjq8x6taO5NJ/DCLSIqgSqFhtPnV0nA9GmgSz/G2384VM8U6m
P+KeWq2ZY3ihRUUq0FOE7uhI8vF3JtJIM+t6SdwpouwtEJ9NTmxA6S2bpTk5zTeQ5S8SBOPLuDBa
30d5n784bQyqXP2aqnkB67A7BYJTuMjwP8Qe3JFsrcCx1OOXDkn6e1Mf3jkUxdSXXHwWV6LImVc4
Q8Sl57tgGMXTVnLvymnoa+Vs7BOb4Kn8G3+YvlKyfGw/1DLqQPLP+gPPxDr32j7wsTLi9qVGpXte
StbmGkN+fEfvM+FpuLSUNYAA7ZfqLXKX+iyMgsWTJ4Xj/FxirY3DrxPQ1Zgzh+OZBQ47SweomyZQ
R3nlUUPali8F1vLpFj2YskSz5nn6KF2BZt7d9hb03LORV+sVJyiA7Bq6M7YmTcoHPJ7wAe0NH3GH
u8e8A4wbk4yzaUHMMnCjC33y7eQ6JyAy382l8+FOzohI/OK834I2JPcYFHGZ7IqsH5aixcWwK1sF
VkSIK0FeNWa3MHge2I78nlDoehzH4Tx83uwwL689xAGhFl2oL6exXVQcEQR9CN9uVhrTtmPzq0rt
wVi55VyZSGn6gXWr1X8GKGfPuQtHl3Gw9ReDM9Y4DxoOnP0k2dkybNuhJZ490I6wKcSh9gLlYk13
r2z/9C+GMRfWrtekDNulvxM4iSzKNbp0RCrgH8joEbtXaB4SiygMRkSEpVXtx8SEtCy7j+jv7tzv
Yb1iqUkfxDDqePgoPvCfZbs3IBOdcOGW30H8Bi4vi/zyFniMejHGiVr6HYN9C/zlLW2Q0DgMTnvG
yQg5kSgydxIVMTJJOphCddlYChHyOTDfWGX8XOgrE03YBVY7vFUjaxZLX9QgBVE+6r1lIEfLze3b
ktngHesiK2hyOdse0Tz7GTdBKoVRCm7eL/CaLIvCb67F73EQkfjpPtcaO+XVnsq7fyfg+ClM8Djh
LGurbK5JwsFD0MNkp9J6xpAiWn81DrwO9uESVGg9vtHMk618c6acx6acc0/9iodeDxL9rV6TIIOX
/N8NP/ZLb2xz5cFssQCZiumSaj/FbXG4eDIZKlfZjnEzCpFkCa5IXiYZWvMQDRglnyoymVGhLdI4
6M1QHmvzPiVNWMGZOM6zCX6Bfaqxfrr72u0FkSfOf+FyXUiqRvPTyuTxvYRtYCCY5vhtakWk00Ou
qMNA78E6y3ncba9ko/fNErfW1Bc7WNzXmrRMUS8w7j7/vPsyOPx8c6+ukxLnuUFXODx/rME3jO5w
ihpJqAzZSrJemO8ZpHoQVcJQobeuZ0R6tgYW6W+dpyShXEw0nMSdFP2gYrC5wx939xboSg98WVRs
ory6U1ijnRv+6672PJMcw539TvgvWf0NPDCtNq65VW+jkX/ZQmCV0SV4Q3gFhXRXcocM9VjoB+ud
BlSKS0qaFRTIMuVqTOwqZhpp2tvXxcxoZf9vbVjKc+m8eZZYO4EDn5LHZ6bI5driYYAJfI9tdvpl
rCVIzwPlVSMTTUUFoiuCpmhXfHIEMJgBZzhCLFomo4uyKcFAfsj3Uz51pnc3aQpGuX0PRzx75XhW
45K0n8oDT+yT8QzKQgQRfudbYDgP9LLh0jGnzQ5zCyZ1bLHBjUBGSwYq9QtMA5/9zFF6F4dXKJZi
/sS9Ysu/WShHfG1d+KFFHmWXgOz5zv8ltRt/ZJ67lOGMiDm9O02JGZ5JRczhojP2pJa3zEisbuFe
LVXo4zPmX5d7tHuYUiG4zBSJiQhW+cZAvGd2KSPwtX/QrZ+5hghzS5vzYLRmcp/Cf6uFE6V1ZRqS
Syjllss1JkOJlmODK9IYLMTnqe1+YaigqjVN6heKtYGLg5fD8o5aJWzghGaehmQoD6yiaWB0jJZd
u+KmrblpaH1uyb+a2fh9G3FYsNN8IV3QFClxjyVwyAak5plc8GM/6EUgGnJ32py/ZmIr5P9uwQye
EUg4tCumeIyXjAlbuc/TMQtlS/6C9VLRezAQTlnoYK/q+pA8fuDq4kzcpRCkvCSMS96/M9jymE18
G1lfdxwu2UDAXlWNNDtvxi8mk5lRSFNSwchfuOVCUavA/c+A13a6QLo82o+/BWrdpe2JVX6QYBNC
LiaIrP9S2ykLAJQNlGvjK/fiHIbtwLNz9chzH5kvjHhdeRNzZo6LmJ8VwEhtq9ytXgH1FnrD4v2L
nvuqt8mbs5KC5pufpU/oaN6hML8OXETXDQvM4rElidFnRBiro1070slsUYFzTSA9l7y1bHs79+cN
4QCVJbWryAXJv+yi40Gyo9aov16wm0i5GBW17Qgg139iqq86hclbMAN5VZe/uwXk0a4lp91Wn4KP
OI5sDWk0/HCtwEEYN+/BYQOHLLL0xstxj2pOmxBwqXXJAKent2Nm6LbADvRufcZtWwJZUOIlsIMM
R+EsC8Da/+cEemEPsKvkqRM+aZBiatvOQXyuqtCJi1j8CChQNOihEXNIy+sBYpq8/9deTiK0aicW
X1jrrVFeZxrY5gkdHAAogHVJKkbie2d3YD2tubuttw6CgUQ7AQHAJub860M4rqOB65iQZPlsZW1l
Hd7NOJn7Rmsn6Wh2FXS8JawqLMPdv1uitq/7sw12KqutJyU6+tML3jo8Atgur0kUxtViM0e7++Ej
SzdtMH+/CKku4l7gpERpV5Nw7K6npHPLRQEeiqyls6zRwAvkpG9aibDwDhMxuJXqdROpg5SHGjZ+
tJ20PK1o5WDLlzi9g2eZVu/qfCfy7TapMMZQF1tUFO1PXq+dIFoo0i3T10zVKqLgG/OADL9WZ6Mw
zW/aMu+TlSPVki3XJj9doqVLuhsFKvu8ZaKyFt6ycsiZ8/7Owz+MkvifyxEbgUjUwW5Sz2nuVI7C
7kaNFKfZ9Ia5CaMqzrRNiEijYAUnf7Hc3S3CyLUt/DCavQKww4iY0AfQ+hChY01gnw6Ucu2PMQzf
sj31sW+JRTPDpHIUbiNntffkHcuA1PT6J6k3LY8X5hcHoScmYzGGvIyivdG34qbIv02lWOqg1ROX
IfEwAIWSFYfVHFKSlD0+iyEsTkI2M490HJeOs5m5Qm33fVChMYRJVFMzvMkxQCofPwevH6wZZCZ2
yNSIUZ5YnRSIKnuwuLiJq+Lkr3NjBABl4v1DDXGNmg5eLiD8EOJ3rVV4QaYfFlfNNIjNIFcVPmC7
iMX87jYfHnH9lUOY4Ogm9e3SqJwm3N8jAqaAHzsgIqJLzKFnSVakTLNJ/cIihtVIhIqRBfusL4G8
PyZEe6JyG50VWuvWsTD0S0gWis6qixAqiNAn91Fw1014RbPmFA3SrrCsnpN3QsyBJ/kMwLouoVds
Tax6H9srSNM835Mt6ir72d5G2AhwaB8+up/Bs4vhO9MoVbasWo+iS/9FAKnp2GyqgrY7S+mVGq41
/bvWGaKqBC7elxkqayxODoqCD1L0EoNRtrYFHyIXChS1Yj1ZLa4GjRJStKiPvJR7XhkiutWZhD66
3Ng8NzApDs5GOXivO4YLNyUxqVkGL6MCQ7RjAA/khMpBPm579kpmezDc49AzbPt6c03M6ukBW1P6
E4gkRtIGZDIIqNPG4t8a+j7cdWqg/qeHgtbnhuLDBXIfin0G6qiCAVe3lnOV6qTvJ1T88wHzb35c
/RntxRhT35RbNqLB6/klLl1b0zUr26SNvlHG98Blt9j7QwqBH+UE8/MFSFDQE1jcWkdh7gnPeMa7
eolO7/5aylYOr4Ji5xtYPmaSduhWmok/6kVXZnjPrDmDNI5tV7GdFNr5hkMOPoIYa1zhIekAPikP
Dc9jkHdt9DI+k5VaPXf9VlHqZ64pwkEKEPf4Kw3/feKR+Xb+MamazZJbANwJ5+iWIElPE+yw+QgL
i7BBOLELH36fDs/bgLxxasvo0mHshKVPJ4jDFfO/GdY5RkHHmDCz2Oz5eHY6VLiNP8QL15tL1cHn
4Vq5ziowWakCoQQ4q/45czs5KixVCb0oJ/wrhO48ZXdnSODMj4g8B/izbVbbn1x0IbMPYVD/3gAb
QzJwztkW0U5zlp6JSghep2PZubc8nqZEmZaTd9om8T9foIojV13749NDjKLuJuoC3SxIXHxBgDxv
vkkPNukhfxecZzBM/8KLcPdEb97yf+M7ZfvZlMBKUlwhO6/lo3s6ob1ZxN9xiGazuQfL3ryt8LF+
EucRAKIjGXOZnb45yyYEP/vmzMY9GYo6ZHBMPvH6b29XIkkOJW3kquxOrHjEodo0XJB23+XKEmOy
zj50TVHYXPagn3s5OWacVz4aTf9b3BptbKtfrIv149+RHYTdeP78cgbPc7L0lhymAvT40NSmfq+P
CwfzVsfQIRE9L2xmbDFC81EmlpDi+eeD1J7LRhAYKlGrkUJ4F+PSlf6k8dovLkvh6rKbL50fX8Ou
k83DZOnfGUu1SJyEodELN0Ol9GXxe3PEtDh/tu2KQIeqKPc39Yb9RFV7GzuWuRBJm6nbeG2PTViM
yEmZ0yLgEwLhA4nPNzHQQkfloUOBuzRwHF2SLoVCcHUw473PEY4yzdPnmEvtIHVenBJHWf4V29OU
xkKySzPBqKTU83JD9VEJwMwQ7n89x+3NaYaoHSIjgv4/IJVmQaddNrgSlWF8ZygjzpzAGNhrua33
IOAUOEL3mhLYjsxG7Y44KKFmYlMXOx5gNVXoZc2ftua5AofvvN0PqxE+1q9uxFEDx/pqtIb9Nl8a
3YM3Nq/vd4gchP+Dpt09iibMzLdHPHZuhAT2eW4Vu6gfcBuAfZfFnPQZFUgIjENr03KRcBNGPNaj
JcI2kyCPhxZhruvdjKH950z87ttBHOg6dPxlpuLg6QV0Ex9rZyTDSb6ykB+VVL/PGposuE4Tinm8
IEh4/gwBYBpL6USsYiq6SYbE8OAPp2ZiCCFZ1O333+gOShHgW/3028+i/9etsIgdYKEcaaLYee0L
sdNBMohN9sptZA58Wqf+ehAsaLTVH8Xj9vv/xzT83yREkxZatLwHmNUikz/QSi5QRcw14uf2MZ/J
5bKXSntmlyGv4QuHxL7orRVFgALRaoSsUGoCAmc0Cs1u9TmkbxpKS8aMkp35pbLEEqdBC4Zh18Fo
2OsbjJZovKPSGihrZ+gUJctkyrA8qddk27zkp0UeqI/cDHOymWhydJ0qxwfBVJ2HJ4nsAKtwqn9n
qATLKKTLYXWaRZbgb14EZvIRTzTEmXppHgcgaCxNMZZQdvshjir7gggFkBw0t6wiAtFHDa0Mevy7
BA0K+Xzlz8QQjWNimBJwDaVWQF53BxuI73W/NvnwiQKYTLxIKk+XUatzNYSceuly1GAZT8HHfSDt
G9wjYpHE7QRp1uDxxebAE/DWQBqmc4RnimAqrj+HTu9K0kb9D5t0DIuo4GD129uprm+/JxRZz7uQ
75yWr7DuX4Js0O07op98pP+n02av5ZmYTPqekTHcrng01Bc+FOEUw4VsNmdQuiyKIdP05tpZV/ji
ndM/tr+xB7QRY/AONcY1kFmM0vqKL+mkvzBKzW1wMKz+4y48xscbshHK/+Y0HGBi2mmw+EGPFUDE
KaDmejptTX6fHwWkPcoV3cZlqq+zm+0RJYLrh2O0Ub9OGL77rb6hFqkRL1OSd8QalDPHE8+8hkDm
kaSuqwQ3tIw5t7trPPzuDngG4hNY4YB0F2qidRfHCoe3Cflo3Tm/ekc5/wOdToZtHbz2SsK6mX/k
SDRkr97ZKPx1FJEolDM5c7whZjOwKBR0uSF6CGpcJCyhRUb1gLJPaYfi5DBYMLBHgmut9pq6WkvN
zslLmnib5V+zF1eowVGFM2ntY79KyqZ4ZRdL/4mVkwDL1YyX0PWnRH1zVL4L7NNhUs82S3hAeNwW
d1Fu48HRZxSH86hBJaJ/MuTPipcuwnRteeG73l8DO6NcXW5+k/hvsmjG2BXoVwlqETRiuYS5V0/L
/G3NLoJAtS6SBJiEWyKeY33uYfqTbkOhsQSlv0uUJgkOCN9TyATR5xVXqzIifMQT+Wq5QvClgyWL
UXujcS/0BmVOnn5ju24Bqbg0Yk7KLvDH1ItIqyHZwfClNWDGCyjSF4xaaP5qtdqCrwlyTrTs6qCN
YW3AEdUqgastAb9xl/k1dMbAZjqJ43dT/vgbwAg+7uAcFBfS6sBkzAQjUx33IBIFtMp3WcoPW7bd
ipjgY+M1UMBFoLk0ZvkuiX58YQOuawE2A6retouyJiCNK1qcbCsjowNE1xF9SbUgdZXO0StrPejY
qtmqYA6P7wl8FUDuXpmHkuWMJzMrCV/CNdfUSE3y6mj9iYuoEHCqeBx0ZgTGqTY7860kzO64zhdO
FoOC6G7zalsxNnhq+0jrefzoukCYyIm3sPcijNWz2W6fJOk6KgTadV82XEusGOtrIVvDJdhCrkgf
xYJw9KtQ7sVMX+TFP5FjHUwisifTiX0RGRS54ruEwSyYM26fAgqlYPIMeors7ETHypS/K8qN898x
DMP/cpXCXHiBl9ScMgPqJiqaxI+ntUN1VICuLkAaRVjwrFZGbb3BqvQYljhPNheSmRdwjxSw9DWe
xX0NkJFOrRYRvXXNs639s6cRPNpyAsBvGghXa4c9c3cd4dyPLLbFlsRACmmqDiMyERSiKM36eCvc
8hK06ISNEOmJjJfBoULvn79jbiRg3Alm0EOswerOdYDigbmUGfei5st9lXCsbdelZKLv0vZovj3w
eUXahjav8Pebuj24bAfMU8WSe8lwXfdZm4OjKFZPSxjzr7WbpzeL4nOg1RY1rIYSQlriVMdVEGVG
4EEaQu17L6UU2NsrDb6aVTE1uLamAMMXmTiSa3CcRFfQZ0JKGVeSU1xlURE6IdWfoEZgiPd8wuYs
qn9eLrIFNta48wXN4FWDm0cs4wgLl0c/NoUiB8tE/Q4wdfZwJcdoRe1BYinsgn0kfUY57Kstx9eI
xQVMOwbj3W/gXkXsWUCS22cSwR5+uPxVyY/RAthFjnd9h/EkTQNrj6FwExf4UXl9oWxxeLv1kAGL
I9PLUs6pLGyp58HMEPebK40PUE+vINv5sXgQ/+q8MYP88KWK2mhG74SjWmZHKIyRLSITMYll7WX8
P05zqaaRQvGIxRkJVcTTc1bw3+sx8uHcsofboxXiLWVuR2Rhb/dPF44YbvoRlXGLMOG05lR7dhnw
L0R8tK5ZnkGZsIo77wvMTliuKoWfE4IaZd2ixTy60xr2uUHpTBr8o1wHhOALnqc/NUimqjvp3W8L
Qcsn8B2ntqyS0bawBU2g+ymIkbmuY2yCU9hdto6OEnZc7klZkkA175E9JGNBs5glmIFbGqhnPR0k
wMI1/5EO8d6RX0EL/0ccuK8nB3wx5jsKoKifhmMxQve1A7P2vemdE6hxVoCpnFULkpcD2g8swjyg
VF2I8iR7hZhfvbowIVjCXjveq7hk+exSKhZAaoLt+f9IPOW7DYfkfIA3ZeTvw5AxJ7/ZxL77VGQG
cdVxX91EwZr69WP2VVy1FLw3R3t5Tsx07q4Yn7XqI7NitWzamzxBeGvSlvQPdk7TMsYqZRaRlNB4
G3OqJEn4ncXPeVDTHtfUvnSVRzGJ2n1YmTzHjvfjfjpHF7QtmYWylUjm6iVUt1IXg/K/aqsLG2ds
QwMcXRxhcY3nN0WJGYJITKKmunc7x2V7stX5bYPQoN05wsEiR6nfKOU7eygwBZsnSJsU8l+sZWd1
zwi1NBETtxyIMPGhUq5C9dfB0lFtrrRlOUWfS/C2wF/wRhkABWZ9GfKLvJJluFmNFr+DAiUMEWOC
RiAqT3YzqgdMJhTVLJhOBhIF7/v0DXgw/FXHVocxKgbALoidRJxF/1Ckt5AGDxGz1H80tzdiX5oF
g0MB31iqCOWWuUdy6litdaOZTOYzT61GIoQ8LW97IQjQW5zfk+FhKbfJ/50nipIfWoq5ZqwH+OjQ
vUe6433yyyG57YyEhXYWF+KBG7nwnonJCmpW1xiqzOTjW+M8PZ2hCI966Jkdej/yaiHtGINu+jHq
lfEjIwjwhuz+0uhyFrBgrVmDqskWYjxnFsyk2HZI2yoc10RW01pxu3qH6ie2jG5XjXQ5l+y+owLM
SP9slEJvsXrbTvwTAYCAIYho/1RolCtPb7IIG+XwUIZcb4pW1USvBJUvLz1GVWt+PDzg2whWnJS/
CKbZ8khwk4nB9Q831ntWt8wzyDtLssIGYHSgNl4+JkO3BFjF0hHOn5Fe/jt33jTcPKbZctSWCo3/
tF9OLiiZIC8gsB1q+gbd47ke8/GFvBwWe2RxsDms43/S/0HV2dxadxg0/x5IVokrfGBU2OdHg8fi
fqvxK1kO64MKTGqU1LzFPqmQ2TJro+LwdHDH4om8vSiLPgnni0wsdaSiefm222sI2j5acclWt7La
ZXUC2dTEnYiKcOS2cp41syv+d+ahJu7q0SrBPh32WqcZB+/9Lo1n7LX8x3iKjO7H7eeSnpJlfkmJ
AMFA3czfh2e1g5UevQ7k1y/TbdvaZNeQXufkvAaw3zl3yX2l43w04sEdzYXTR5KG8zNq3pw2X226
2Vqfu9yLk1wKlvMcv4eqYYUEiLt2EeQugcS3JKDqnxmbId9ec+n1JaDghE0OieVf8qU8zl/cjaG6
48R4L03c1ylfTntcyUcR3lsHwEsRS1LWXFJZAGPmZNbR/nnXf0B1G5ILdEGJrzNta5dqie4rrBcD
iuSOMl0w9EK4LEdKz+Uowl1CyUAiK+HAIXLnU6jCqTneSWCeEwJptngsVrphk0rcjFiEb7INdsnC
2pUsPAXI5HTfbY9BygSxsuX4kM4WRrf/esJySJUojgteBdSul8dGGyJIJrSbOdeFfUjuv2wjeaIK
zd5JeYOr1jcEUbNdHX5sV+TqFwU9Q25vlwKPofJFk0KtYL7BRY0yiZnqdodTj6AcI0BfxynRUf4C
3S1mzvWy+cCoe3mIHl1V9wGDf1jxy80YXsYoavjMg3EIld3ODcHF7ElcAOnhyXHuWk0Vg2zeqvIl
Ftf22z1xonTS7O33wXE+zz8NMySBg46ZX2qvPZ+Kw+t7pE46GYGwF3WuDdeq/pdTGC8BEp/bMwHs
cV4/hQG3fOVSfc+aVEi0R1PKtxQms5vAWuRT+m3uN/kbhM7Q9S3EJ93l8N4TNW7hPQKI34so2NZ7
HqPSF/rUMWZx7xvNXSAb5sujGSGgeQRcmmb8pSPmynA5AsEhRhw0hJvE5yaj0f6Qu/tEnD1+jHVa
XKUcoSTfjR6vsUycBAriVG8ypwVF3dJ9gAquToDTalYzIZcaJSqe6ekGkdmkvXR2dWwYZtYA97ki
sV9Jg0M4OEE3KKd1fODoqQe2J57XQKHQwugxOsY5jo50iAlY6GM0fQilw8RBbtmp2+jVQ1QSUF8k
zt6ctxtZHzVfGaFpCkYxcgEheZZe/tsjcNEPVqDv0436tZ3HfSsoGykemj2IrmTcE+ZpPq1UKzpt
koAnbevpl3nOXLekQ63w+FoacGdDyQNm282MWsD6CG5JxMXrxaZtGdzGXarpzwbP9b+p1EQXEoXj
tZrmtu7+w8X0cynLnZvIwEkFmgcLZMtUEiKejAFniEfPf5wRP6KjsP3otD3B1gKU3oA0actSzrEL
gciUi0v1FZ0T5RiuHPyryYwG8pXIqbds3JoNEWcOsgc6rZ1nGWkpzK8YS9rgBTH7yGYUr1sr+cJR
9bmDtHyHGENgBO8vSC9GKAdTszW1bgOKg7I8K8lrHraxyUbdRFm10jb9fY7DP0fWbVkvG5IJ9+uw
9ajk2JwpKYLZ+PwzlCXN4uiJnPUQD6VR5u1Dqpp2WOmfabQMccHstyq21vfBV62U6/rCVYKIv+VI
j4e5EHmMS4LQFtZ2gq6/QJEkChE2cQMKqQ3nQ8exriS0hU4BPl3sGaN1BAC2wvoLsoXiYKu/mBWz
44IwivSTl1WwQ3gbx49GmHL93qJ9PBVwYuiCv9nc6x22QjKLLyOH3kvMDK23KgcfxhxaKGt1HkgT
2+RQKF1bHHd/AoeJIN/VaEypOiSplNh3wzNbNSBydmZFiPAFJuzndj/0y3TkcYDIniPAvb9bqkrI
NHjXl6+pfB1EfGC0Padc9Ro2AGrizC4KphEv+WKv/V+NxgGgPAyj+K9WcoE3eDyj/Mp7TY9w7axo
TTtiYRNVL0NGkvplSEOiBj2v8gwvmW/wMrjuiWZZtma4h/vbhnNKDj42qKdsigBrtRYezOt0dmdw
2PnoTtPES0h37pkLYVUxvJkcv5TtoG/Rc46RkZsJWnKiEvJOXgIXz9qDGje4A/XK2Osjc8ROnWEM
RblPLqxi+IBrTqsXCD1hfcwv6lGIAv9GO+PdvJqjQhMpqvVHfZJCiHoz2BOLUUIVOIy5FeFlhKLu
UPzlNgmCHB9AjkE9TTTkG/fabXE7epCTQSWEPCSLL0SNn3ka9vAEd3ArQFrAeJhR5L8kariEQ7vR
m5CPQ4l711ovcSb93/0dYWWor+MUvJMzZ0P0w9pW4QZSMOa/AmnLkJfKmpo/v9iVA+mivFGk6cjH
Y+vqi5I/UuY/wCGvB7x39UxtDD406oPE/2wjckmzQgg0zcYthHaS9BZ83DnHqpX1VhwVDADdrTXV
KKFc4Yihd0UR7m5rnDPeqqYch4rQF5TOb12CQf27VTnSHj2I8Nu5YJ3/9gv/Noy0TBFf7h7mFR8D
Fk5hKHexmQvTy+aJ7x45RnM42e3Lz2RR9Q3/tYN9DWBkgCuMsrEG1zFvrwk10Ny57/M6C/u+y640
u1OyR9h0eF1CIFZFvdRiMux63tuS1vDzzrjkKfhauNuVehU8+Ccw7OumO+idSa8IS4yd6dp6citI
1QKkuj5bB49AXsHIZ6C+kzjCJEaeu/w3zmD76SGcE3dQr6BESOirYFjoi1R2vk0siv+hYAnMhvYY
/Fr17R3VChgcAFwT8GT5lPeF85k5EwxpIV9IE2LEjBt0J56KcTYk5etxzs5Iv0/81gx8OgkSnoU6
ZmiZ5caXCaMYnWtYxrnJxFM0izqe6/3L3DY5zKiviZIljGNZu/hXDwGrugYBd56iWLv5Q5yDa8tx
KQnHl5cKXzQtVAVJPZebi2uIoyRjfcsbayXJSEsYea+QzlPordf2Cutzu43AOMtmRbEkyE0hDSVX
9jWXZ63detMMRIBvCs5/p6XW+g+nd4GLTS4e6rJEWgNuqqsJypExYNLWxLiggmHQ7yrIBF+7n6nE
A1OSsSzdLCLF3utfKwET8W2gpEvRCGCtrYbKxO8u1YFPR9z8pkCynAc24+jYXNvLBrhyHGe8zJU1
VmcO/0GzjLc542XtvkwuhxHcgOz9Lf7CIFAiCMVMKXmCIE9DJZ4fHtGaks8e2KAv8Gm1ZqSDYWec
YI9kNhstzHdAMbs9EWppCX9Y5Mhhv8TCLrb0KrcVW4M4+8P+YMIy5eYrRhNwsSSC9irGLCOcOai3
/Wo0/JDtQuF5arVbyLSYLOMQZp2G1qgwe+C8oEhcNtNaM0fNbdsn/ThDxvIlhdqjmTtfughT61lL
QV99uTrHj++3Dt/OIyZO1fWXKMbzV7QFZ+YuLWJ3O7ye0q0gwFScsoIbsGV+R72ZymHzoeNagmGb
/xlVGEE5abfjCdEgTKuJZJveNaczg4b0SSJRYHTtjYsieljKBVl0UxsXOnMgDVOwLmgB97vv2qz9
jy8sVpgGxeGA/Wiq4jWe5V9BwBlMtPkO1EmVektumBcOYFcGXAuCCi7tydDYC2WvqqC0YiTx3ub9
vjhG/x79mz6pN8YuMTBsMYPJFKYtfV6tuFJZZ+L3fEcuJh+DMXNW17/Y0b36bDwCrWbDCCKmXtHJ
BhkteBymmOLLQ2TkqCq9ZMxpNKsvYe2A3GoSIdnCwNfZFxzy8Q2HYLxLHrOXZUP9zqsTQYg71qak
TPiTFtv7CEKu9JUzXYspkx1EShiGYzqZCCNl6o37sgs4s3/bqhjaxpEKrbOTkWW/S4p508aMCtS6
eMglolU7vQvLvpjvaM79PK+GoR7Iov4ihjzl44waeUBKhaVTU5+EvW+rnsCBm+ZPPz4m+FeFhFAM
zf3fEac7mSLjHS1AM5+ZRZBCFpCP5Ay6O/WuPydbx/+TDGqmEw+6cQ17aQyYOrvAazw/1Auk59Y3
DwoxJiuJMkEx+Arh4BXLDHqO48zfBRkMoCYqGFE8Ct7txWKCv+egZT3RgWpR/kzsfspYX9zgqtT0
WfjRRJHJiX/HYoR2Bw5Sl5Uq2RtbUD9MFwdNVaoxF7v2fiGlsicMetq3uVTmEHFmC6KmVum98TlS
ZrK1m79U4//4mqG6YfSLuqBn/rCgUaIm6m94I6kFDu0ByNot3zZhx9l09RvEgag6R3aH8rnJGlnS
249fehST5Ql4PKZWMfA6QRDvtoHDMPHK0fXstA+gpx13/DxhgOhgyRKoObvsxq5edQkzknm2QA96
4Z/EFoy6eHTtZdQ0VkkGYiK2R3UDkOhwUoa78t8Za0L7LAfVO2PdX9YnxHYOEPaGqqsK6KYkj6xi
+8MNLXr48V4Fzb6s0X1MMs0xqfmzeSD8COsN+gJqcQxiI473uXALVWwu4vTMuHb1AaeA0CaTyC+L
ogsZgymysOWIwkUZA8kKTHwa4++1WE4dhubx0oFMjM7avrd1p8CB2kGOsfBzzqs7rwEYZY9PB0hD
YpLwjzZCD7JciSB6Jyy3wo/tTznyLSnt1jwLCxEGAqLmjuKAQVi9p+0Ogn2EDdQ2EYqi+x+urDOw
cT1tkpQ2nMCgEKb4zjP3aozVYn5BdOmJauXr4Ss+SDCbTX7U7xu4b4JJvEhsYZNzxn9UbjPAzbtd
b8w/hIduiq6H68sCOoodljGZaECeUWgkDh8soQfC1fU3L6uxBOSQ92EPmPQ70iKyfsdpZePMzkyO
xPzzvURobTLgO1L4NoJGJ/T70bCBnD59TX8VoPMlQrPmvSdak2t/YotWzdl0bR2C0vNsIkcVDobC
gwKkMEWtqPrBK2VHX5bvy5MW4xQpC471HxcwZIcOxzeVryIhJYe9VUPM+60SMqOzwkEwsBoQlrQS
IOVy7rxLjSy255tiPQhxOqlxlmhEYfgAbQDL+sDrrEe/5gTjz+OpXnWkzyMq7J9t6qykB9iWG9+w
A4uae8gyAvSN50Qhx2G4yFRvGFx6fLQCQsw4yWV6HR8TUYvIU4Da6Q6OQFAmMbOiJ+2MaSppRLh7
rroUVGK/duC8GdyBdvfR3miIfzJn+wsaSq7IKlCwc1AOv6jq1REegLaSp/0LGhtB0wMVFJ26hGtt
1ZQJ0r5XD37DAPO2U2EgohrfPlyxsoOybS7RxDvV6PMZnaHjBnuEHUgK3jrgzGWBn5w7DSbdsiid
ZmJMypvSb4x08LFHqOPU5n7v6lbMAr7eBr1Ta7AovP94+SiGGRh2rWiQiNO1dVOuHjzHOxUrzXqX
Umidzg/Q9BFIgrpPmm27YVmq3kcbq4lZoU9AX10ONJV138pcHLC+RCZFwxKXkLabpyBv53zYuSWr
PwbuHcU4Wcjqe8Qtf+631MasWDb24AU8xfw4YQQkuAMb2FxUctYcg1NcBUyA8y1ru0v0shcGwmX0
clLVaxSn0CQTW+2p105kA2mZbtDCsCOYZ0SkSEdfQdLKJQy4+gXsp8H0jWc3EfN5qcmDtPhEc3LB
pyH5Hkw5Gv9Qa9prVhfrItkU72l2tmup9fTIkRlaNFM2KLFAZIfMUgv/4vzXQvOp3AaDoXy9mcGt
fBF27c27yYd8q28uiWRmZNdPOKiz9HLzFLK5g33IvkIBIQGq8Tr8aDYWw5vedfhbAWbPM7G49d/E
rElXfcCEO6bsyxJqmg8XKKmnPIVksexrwvxrM/eVK9kMz3g1JLV2Y8ki+h3vBr/UyAe68bevyEbW
Y8VZW4oQdyr+X8c9VI4KfjmVq6ZqR0nvphGNEe7oNOMVZh21yo9dilY2xi8JARmu4PyiwRNxoBPO
p8senPHCJukNARL0QbFleIVFefmx473/0kY6aLSEuAIaeQpQy2kB7C8KTQGsSNsqgxut9TE/9TWX
c3yi+Jj4WbbOkRvcNo7DpG2PLj8jvi5r5/A64ReF1lcizHlA/Q0NDhKMq0r+OGS4PyFMkfCVx3Jg
qyOlcSZb/P+N2JWeCrXr0URG+wBSMN99xurMt7aCkorgDQLZvJXHwa9NiPsdrZx43M9iN67xXuSZ
hauZEUHWvnG4Y7onwedldqD6OiARdAlPOkgoBiYkYRUm9N3uWIX3DlfsABTYhy1Fo27gGcGXMGSR
w08KGhr99bqG99Aa7xCUErOnSP7v3LuW+F8HcCJ+k0HzBarbkNR9E6ofjhy7G05G1k49woOapIrO
r1ZobzuCD5HIsygO/5PUsMBxXLejWojNfOicbaNyxM6GUXC5LAGnR33wT6HXU0jiptxCw4BWilgm
10aD27wtsgmQtSFkvdnR3LT4l1qex7FjjX2CmKC3mZZJvVUaq6wZR61oUIeauZrjmD3JmmYIJ5VE
r/YORpOJwRtpnCVh8QnnNk54ofnxAugXze4bmeGCGmYghZh0H1ZpIfC9GKcWbngUIQ9NyzBXeFGx
rhe/j8eBtEEl6fUfAXwF2W/Qtksxs8/TICC+XSXLlcqOIlK74rMq6ibPfg9VcAj6fzZkoEBYE4Wj
mDgKEyKtzjnD653MdNDSls2B7PGolu5w6bdp7rS8HzISriyhfzp+1tIoH78dRN9e4dy1Ssds8dG4
0l48vwbEeK6F4QunvTpO4ps8w5EKgK3Yy/NVU3bm1+nR2B4+BaaqV4ojfqDjE7pWur1b1ocP3PjV
XLDCJjbJjUuV73hack73bB90jQDM3yek3yGXGCMidIvdAb5GNTgHUcE1cTBxsB/iy2RsfCg1hYwB
K8Pr99BHYln+66Nzi7r3yID9Oh7hUj8+ZE3mBf+yPfsRFrZJ5NRAY2c2IlduiA+rSR3b6GsFP/UU
FHBwC1jYsoCRl9Jf3ukWGXSPRlhadJ6euMgfyEzUuAE7IS/aQtDwaOpJBtvRaQvG1azExoEZOJgf
2jP2JGJvsQANi3ZrNtshTfX9O2+T2g6qR19Dr9HQIiMXYKW6Ee0F/XUUeHCjl3lIoH3fuhSeZWsw
0D1OPihLEVHPwsVnEL41fTtOGSA+54VOmcFW5e6WHLKg0w0kX5q5aQiEPtYiy0eDOF9MsLZFWW2w
PTGd3CdL3AwcUXZTEW//+WGxyddVyBeWtBgaM+jjL7UVKQj29Bbnw1dy1SmJ/wELWe6UInu4Pbpv
9s6uLHSPkzbVZKfPex+Jt+ckDO50JXCJIrde1YDOeHr+0Y/OEkXqAqVZnDtDj9AcNuJElTlpsZf+
jPxLbGMMvZSduzwmnYmmEIk3Mvv8Acx092VZhmyS++qZrBkAFwUfT6C8a92CMAEMvuTHGMjY+V7j
+LLm/EQ6Nv6cMj9MPFXGKkcCAdbpqecfnl2OAS3LR7GM08wI/NCo3e12Lcay/I/9bB/8UQLlFp5t
Y3tU2sNVzjFzay1yJoOzC18hneNuLRXnwIYtcn3r/TTMUHwO0uuZuy02BtqbVDmi+P1eVAwkvHgT
yhsz5o97q7ahwoHU1emoEWgWSZ3neWQYmD2u29zTB0EtUJPGy9e19Kk90AbfGYmC30X7Z4N3rdU/
PCT8i31utMDVQay+tLvahbNsQWpoumcfI0eDRf2zhZx0lqcFwwbH/Fny3M8pdlD7PBIaVSU2sB3N
NVUc/ZOLdFitdyNeEju35mD3NHAPSo4Ytx26GU2q2WiIqV/xVJU7E320S+u1cgHzbuAKQ4gP4xIe
fxGosh8NP2ys0brp0hKEYlRODWRrSSz9A3yqxogB/P1+MDADW9mXVNenM9tHkrxPK+/Nr2qP2Mwb
HHIkzcqL6g7RQU2p/zhmRLI2t/ZvfHRSA9MHuRdEF3RSy0d+R7vb5lIqizWjJ+SSOiQTWyVAF1pJ
26CGcf+kHd5WOf+4gY9rnBvUJ9WzfXfpg0vnE+DUxfMZaUqdHjeUE6/B3jdkvp/VWD63j8ZN8Fm6
6Ie8E/cT2TqKOMOWem3Wxe5UmNUlCKmboB6b657kYYZzVaKrnoGTjEU9NkL0nnazvAjh/7bJKtmX
xrPvGIrjg6Mc8mFeCuT8gxp60+BpCepo70gKIA6gjmrMQwFX9tJ/xtFfEECwEYBu8mHPHQeh8AAj
RjS8DWr5s4iEAwiAUlAXt8znCAkaph3+Yazfbvkcl19BpN0x0L6XUy5ZzaVSI9HH5AXqWebjiHQM
ZONvgv/s/30lxq3g/H65dc6XHuJlM/c4n5TlemATtiG4GXk6Zauum3I18MNOOVUQXvivhbdondSt
YT13J+EeCpgI00CXBxiyALr6/2Sle6d1bthSSMlG1TxOO9JPnIdkl6No+V+CnV5hFA2a1JfpoLT6
892G9IuOI+qci6hwsPavc9JTc9UoB41zuubW6NG0LYoNhcTD/CZ/a9QzjNh6yG9Krlbq3q8Y1YHD
Q7HLH7CjU3wVtmk+wZoXfro/5iKRT9D6xtY34yzw4Ezy9pKMlj3VnQjN5VzOYHIXhLac4osYpUQ+
mtyB2goNi3zuxMoYwla7+iGWbXYQRpKiGFB7ucYqIjZqGD1UOVOf/dQfX4wsXE2vaMFtni6OYhOw
0ozY7XaXpuuMDKtKFks5IT8QLve5zWhfcST6abxwvoHCCSJsdUWcZRrwmtM+lo6rJ+hrZ43HHTHm
w+ZPH7VlCIq9JpY4hSNj/+Mk3cW0FuueTPL7HSRZe4fUFTnHXnWbwrhC1kSQ1YMpV754v7uLFPqx
p9Su9Pzfo4ObTkFEq9bu+Stlf20KQlhRCwIyQkHeJn89DeGJbUoGnLxrBq8EDh1B/xigy/wt5Ygl
5X7VZYRYX4FAgR6wYt1bGCc4a7slYFoP4pF/Cu7es+XsL8qDo4xF773mJFRdSK0LcaMNfocQoAdq
6qAZ5ddTRPDFSN1PhKHGynbDASb5vWjv/t7PbEWD7cV236gcwhuxsp7xj7t9kjPFH+4STIzMNl1Q
TVzR9XeEoncpW7H0/fqgtSnRFh0HL9iAH29x9QoPtBw1+2b9p6T7xfOvK4D/4nHITutSdlIwcFb7
bWmsqvkXhTasr4AB8nXgb8ZcZUF02LmeeRfgLhcIwtX/8zwMn1NSMadJrjExeZPR35NCyrykRYRq
8KuLy9/mOHSPDKhnrWvlqBwUY0SrlwPs6Imud626spnFYV/xQ+hP79+6D6vtZMHeoewgPpnjLZgC
xUowolevJ2QLW9bhI5SxOjD0BvkXpUyplVVK3uoxWlcQ/IWK+D1adcMTWuX7MzCi0717qrEuAqop
BpTHVnlI1b1jXLKKPPWWDYAQAdJNkzwWY6OP1wnL0gAvVBCSE4R11Af0VdTz7GGoYlyzHGyVQboz
QIB1fS6USNjka3Rwd5kt5/zuxlAd3MgYLSs2CwQW5ToWzJc4xxbDq0mxsUtcVd9UkBjJAFm9KB5+
/RD9H79GLSEIvJM1rLYv1uxJbSfbSwnuwSs+49pj1tcwR7+NG3mGaXk3EeL0lxJOeyQjIrpDBROx
3X53wMvbm49jnJpCWBcCn51DI1Gmo3+drIamQSqBaBb2gQ/Oxr9B+QUb19FWHQxysOyil/Ttdfwn
3REOmyARs1swK70mfLV2nfs7DGaxfeJEjnkGkv/6FZ0xFupiX9XiINKNRK8Xo+w+0xCdyBx1e+yQ
Klo/ryx69/t+1KDXuKzBfNIaTQ0FBDnmadhBxd9KQvIyBeg0Vf8tbYn4MJ+9LiywKorcQy3CZ9i3
npceNPqnTYBIZkilpfT6n+VN13b47yGvesfvCsGEX41Yk3XM26LXCdqH3JqiSkBTKpg7oqo9OlkX
oCGdDk8QMhsDnJHdd+qRM0HUhIhb/DxqzNuPovP0Ayq8u8B3GR/7Y8L2OoRTYPrJSbKMQsgmvkvO
vH6GoQrfygDSJEXTM09Qs+8E6/PFdinJWaZErnnzwPttpCFha21yueGeqU2oO90fiRBis0OR4bH3
gVFXm+zbsTDpijXY5N4y7omKEsWT+CXw/updeg5W1a0YkGi+/qCu/H4dNZ6e44O3CXfXg3YcKTDc
xKYTr3yeNH0LL5Dr4rWZPYuzABd89WLcZmFdBTIL+J8tr7SsrH2TbYrRuw8fQuvH4S7ottNAEhUo
oJFN/bSa9XZgBy7Q/3Q6bVFTFcR1YaP7o7A+5onZ3vJua4GeOwrLGJRjP0tdCwK0AY+ZmvXhB6iI
HHOcRygeKzU8cL8P5HE+9TWg2C6BC868Yaa9qACOACgOu6ZzgI5VWHg6LWjlaeTgUQj2rgxdXbnd
MQ5Kx3+0WjwZYQlINUKTmmFhK2o6OOZnX8ne3CDaCA1TqXw6AFyTZjq71cCp1tpVNCvXCSyQv3ZO
FQcbid1AZQGcuIVBj643xQFQ84FZh5vRH+E9jrZJUgTRr4DcmmwdsdEoaE4U0NCN+dnIQrglgftn
Jng2ZQ+YOy/ji551O8U/t51fLyNyNIFWBlvzzgRONzSUpNy6QRKVtUg4FeYamZYmTvUNRC/NzZgp
lQZS+IOm4ILG+Lj8DvVVbBnEeDF2YAQA0zedgRylmXb1KeX56DMxNsPoTfY6i4OhA+PxFjtotUeP
9oaQBuAURzzKOYVz1ZuUvuEdg5apQPVTT0CDm2bEN413VPMH21zVE24JSV8VuGe+vQBYCzW1lBOu
5O65tqlTlbtmulwtzVQXeXGZkw0obVYPKXUDBjxPSoVce/OgWXGym4MLxiSxSjMrU1Nh6NDCiyL3
sBT4b8cnXMSED7xdv4wKX1o3/aC1Aj45sb8EtrWp6PrjIsJx6raW7ugJSGjti7ltRPlLW4iiP1Lf
8Co3kczeUfpp2zjGOwRWPMVbnkNLTJqaxCx7+clFnn918wFT3CwLcxVjdpBfdyxtOMTy6qeOAW8q
dEJbtKQwEdhMMR6y5t9jPC1B9593+OK2cdr/rsLaia0vXR9iMXMof/iSahiRSLRBebWRNmAsSgk5
xVKoHhyyTqD9XYDi0ffi+XrrnejTklLdR4QfevsAyBp+B5TQ/29sAFKbxvx8d5C1i/4MsuSf8Oth
4s8V0dv0WwjLHYXm9SDbiWo19K+OyVo2qKv7GksDbp8fI59p2toeW6oruNgnpKRsS4yc8rV/lrkI
QM/fI4uTJb0i4h/s13BbVd50TMelCyP7WGPJEf8G6OsESWiI+sBR8u3IxZvT80YxVFZJLoP7aCYc
W2kSuNeNOgZrYMmUmdjldb21HA2iazj28j82w4Fm+eT2fk4nKCiQ/ci0/nLmxjJSMPfsogJbVXnq
Yh5vDrn1mO+wakQ/NUfBMz7INu2msHm23bz/1w6uLDAGO0Ch1sUG/GB5bmDS7NschEWgoSrDdGil
xvoP7ebd8pGkyFDeuq0Zrhc2G9YOtRF+kr/+mt24G07N82c9cnJOjPBZCkjzg/NLTqghuN3yYjnR
I8DzSjX+9tif/821ART8HWUlgDsdGR53OYOp0g4D9DnotL8P2T2/tLuVB/Sm1RCHLbm5mIdvy43O
5mNVEtheL3Vu9phrS7NxNPrjClvx+sBAcn9oOBnjUfUcCHPJTSxpwRQEFpOpQMofId5QdrA3YGmy
/RzBC6zUdE1ob5ZFltOAlhYG09wJPuxIZ9ia3KfSPqw3/uLZv0+EsDPBm84swOKoOG1e4S0Q3+Z+
bJCu1pRvVN4YrJdKaoxsGcM0J7+7zoJdLa+sxpA78gen8ubMxNDIo+vvxUyrDfV7Qdlnhoim9tou
BjA5fk87cmXjeW8044f5QEax8gMuqVuxrB+IDFJwSOvlqDnKVPNoe7BQUDT5oOUHfd7e+qrELRyP
GGui2CoHwUjIMk4b60ZBcC5xiBkHj70ozljChWYO1dWbd44k42uhUMO0sbVlQe3Vk8TYjGIvmkhD
dkeS04H5mZbMYSkVChGGDjrTdc/siMBBPROJmtNsCLc0UCO1LZY1iHkJWoi6azM4bFVrSLrAFi6m
AV4wfuaXMs5RHDhNC9w+/b+vOV2CdXr/EROMH4VhG3+eRklkhenoZfE5qbWnxmpYY6fEFSWejZxk
REz7cN7hwj6r7xp5AsGvc0Y8d4GOzqhFi/zpSgyT9QwkGH2AQ+gqAoESWSMIumPjnQi0jYdaymwE
IZM+rl0hvhHS8vndtjB+t4PgUNfQOGb+AMKlqGa8teXFaSP+MVwJyltlNW97vsTHaKvC/pJY1dFu
4eMfGasLsVfYkGVGfTYpS2Cc/fd+g94kKxbqM4sPyacY44qWljjIG5bDdiAq+YKcHAHTEXomSq6K
Xkn101nwmS/WU2g13neU6WOy1FGDg6se3s3DAzNG5KjQzrFvER8uf+6Tx+bvWX//ddSvrkA0jrDM
wePZxhLFsD9qtjQiblmE3XyHO7z2Ky7rx7+clBTzpKVbVHuRAJpdlC8IMhqvMbmtcrerRT+CoSCg
8HSQTqmomM6DB2jRBWnAhGc9cdLuMKT3VKRw5hrRFJbm67Ssxe+IiIHbPLr1F6mZzrUkzkUp1vo3
9ONJShC7YxaSLBqJdeiEQKQj6LJZHQ5R2Td+jaWp9pXCvfasSxgrh76R0XtU5JmGmbmVu/uOkDpg
1oigHICbGgKDuK5wLW3EOxa2i3A8yvrfNv2g+j32kw9htCxBZp36YAK1aXL6eNE4XwbxtcNl9b0K
YnBlaLmeF63aNFcstMY2cwkPCaY0RvHM5+Y3pEYMp9vq3WVoRl9XwsdG8uf69Jxy+DfzmOQfMvvp
D/y/nWkUxNvpYplO6dCv9FRQoiUZUeGX3X0u/2av2ha2x1tPb2UuOSqZYLFX9eSNdJKc85NF/9M3
C2H3i3BzCIFKkx63CpcdM/GX5gTGVy/6fqGns4Z+g7gHSle8iYxFVWKiDMvSnoG1jnAT9js5uroy
GQlRN3Q3NO6i/ATzu4EgDUKlEfiTXPZQc2vnLxX6JQi4gvOwTm+DAP6W6cqo5EkibX993J3wmfEq
m5YtVdU+gVoDfw27ERczkd/hbkZEiFGfyYOyt6x9fCzDPblbFnCASis72qMElt8LyXt7U95WFyku
YSXVr3N5Yd87LBUh7czlQNkcvL57Gnn6dxqLE8kIq29Bb63NXezAnR2zP9+astitQftdQ7swDJz7
1ASkKgex+cUxvtscVKI1UgTcvfoxpSOtnNu/ABVQ4gTwXsn0+KxmwEdIXMrbzO2u76oIhH1Lv8hs
tR9pNlkA8Z4C51/Z5+TiVeXVvE85HedaxJuTBie+wGF33QRZYYh12D6tIrsTpIPlzLVB2PZvNcVA
X6drv8CBTO7q6uKi7grt+xQ8LJ/5P/fDloCTv7vX/Hi7zOaJBh3/KoaribSKlCcPJKzYUZVJ/iZU
C4GIEFILhDyBQ6q3oO3CGnun/ckacbzS1h9tzJFqg5xlaowdqOPjo0lISb1nKL1CqL7PUV2KNqdZ
zsCPHhgKdD93uMFH/MDmTj5M9N9+UwRd+rjLeIQ/GcSFon0B/ZQs3T4/NosibPUGLh+yHHJ5EWTX
dqD6kVPJsKygvjlxPFRWVnbg8KG4noM87uthxVXsYVj+SS0KxMv7qdJkSuPGIe8mW9DxCCbxZIPe
znZNKneGV8rGZ5s2xorImxMk28RlnhVe7KNNRErsYVe2kiSxObBsNEsHIJvl/XjjdogIgX89q2i0
WAXmoFQ/XPJdX3DiHYAaKHBrBtyv4GNX5nFNxUbmO2W83sylMXIU4kEiuBE8k7VCWOwoA12rt+7A
Fpkl0XTUvR7moier3q40DIa4D5q7EF8Sv4pdbceO6sUk3oH9/a9wq/PlJaPKTqEwq5Vdodd4qhn6
c23kjghC9fgXHmetNjJaWQbPlU7QmIIyQz9HCY0+63FBmrJdqzqvA1weJeTmW3zbVbYwwcTq6EBK
nBUz945xlOdfWAUKxJ5EFTTin7kO0+jHgf+W+sN8Lai1bIu4NTLqtECr1sNWpzDEnk/RD+YHW4Dj
vzIaCeb8I950aE7bCRxzOHOMcCTNMqfQFSI857tyVXYMJ76TcoFIlJ36DUGEPh9vrzR8FRAnelXk
ZgowyxEZpo8B0iQn4N342rC4nox+BYQ0oAZ1FeV5k/fMYCF1jiGDS+MdtWPB8tQCGiTFrSiI1E74
swi2qo8NQ9m6xDqBWSnMndB2eiAbpKqoe0vjUUv//jO7VAl7jfiynE5KruKdSh0mWd5kiwwTgicm
hsIxQa/N/iEWiy8kTdLUXlwt+04DbPjQQgZHL7pLVMQQPYPix8zlEKhLmGNJ7U1/WHh9/6cQ5+Q5
hkd/940sWJkNv2kMRbUaFS32ec6+UnNirDCMsi1QP2uKfp4Kr8xSUTXJM2L14cPR/DDxa2aZkOn5
mSjZzdMgdDdE5bamuyGRGKzpI4ot/FYvF0BP8fNwNBM9Az9GvdXBdcgaArUKKNgLwXojugduDpiJ
yIxp0GwzrwQBHU0c4HGY+GUoR1RicuG+dlbB84hILXe1ZsYdLqLJ4wswXxGcQxeo2wqLSCzmZchV
8X7aCE/5rEjdFyb8orFd6jXRQTokbpBr8sQKcsXWqLYcmJUchC7OVkN6zVZAs+WMF19JCD9FHNO1
IJIh71T046Qi7S8Dh+eIAyORNC+kf/RI49LwVKG7K2N5jW4SSVg8oTL1HrVAm9V9zSKu6S5yHqSo
s/HvGbLGa57NOzZ3oTE4WTnwtSSDhTVH7f5kczOGImeEIu0Ux/Eqr4RSjiWFiYUSaLfwkF6cvppr
QrVkZl6xyWcsq+34A1VtGoq9ERXI5XLF3487PUxtpLDmYyFFgQ34kRP2xYBUoTSwOUh/Tso/GMFO
tjOs5b3YYcaL0jEcV/styBtpm5v36/Fltg7ygEze5K7OUlXhQunL2HPHknwub3M/Wo1btQJAdAJU
46HATPo5nIY7mXl8HWrCxKpnCLV3jKCokfTiyazXFgm2KXIRsZfeFlihSmGb+9BheZrbZT9b1WZO
95K9+vHdLDBgt5mMPL+t/wb8oy3vITnuNn6oFofPPQmElWgkOx9V8fus/VofXDWNOTtIhwP0YXpA
mLFoLSf/Jqead8EaQGKA5par5o9TsnPp+nzxk1UlDXcPfoAPb1HR++oBYcu52stcwjFnA10N+eIU
47kchfxCNLjp8K16TdLPRM/ZNx15FgFx+YDsMW5JPluQjYpB54vs2DJK5NwQv3q50awaJDpo5ZOQ
4Y3+onF7A/C8jUeEG76yRfeQhUG3rOCpj3wOn/9HeQ581rlMjcsPJctLL3xf8sxFhIhy/K0DTW6U
mljAQKBWaPCwcVQeN5wtlVX2+uz8VF7lZhxM4vzjIwsfbvo61Erk7jqedk9Dlyxn/lBMx0u3vpWm
r00B25kNeT7sUngWIVEcrugTUT/plhSsl1jE6z/0qpNVihmR48A9GaWZ81CBb8RgTJcvZ/YMDwwf
X3wkiddm3oeNr7JpyTJs9IuaWlkGIB1sJCG4kTyHEgg6Ty4fK7zn9JGhmC2EN2j0fad8+dX0zotG
XGQHrJ9Il9RYni6F+363WW0OmXyhnQg3EvnZcZdUqFw5EY0eaYhjjc+k4YrGYQNHbXyfzXd+QHUj
aizqd9QlXKdv0K90VIS1kYR3sbdeaFSGqKqFdLPRBbRhG6+CGQkqvBnjL9pSvKaN83auEfr/8xeF
qAkd8Wr1qhFksAxqXbN7o9Bz3FdnoBT5NbOeD7Z0VsZz1bhFPHk+L9krot88M3lhE7etOdWYLOhu
s5aAJ1z3DRyPab9qi4fwp/CuM4fX+nix2yem4gkCj+eFDy4SLBcYbTKWN5smWQ3h1sYQf27abbQu
XKRjb7jRjPBlYMP6UsoRDjTar5JN+n1Oxcw22LBH1yCwyIK2oYacCHfgCxgtQisCWWrDFa74iNBu
7/K5k6wBnEyP9ZCokS4RaR+cRT+xpPqbVImjD/AVU+ZjKxZSzbYwr8nr2FEdcf2vAZz32px9xF9B
b0QMwo3l5srISc2lPAHWFjSpRILVPxaNLtWXFIpEUPFC0ZfkU5zLw5TESOjB9+sopB35OLz9CMHR
fP012FmVgZetVmf4QXWhUvLs5JEni+CS+1wPutEq7Zo06vEWcp31vP8d4CGZP0CAYSV6+NKT4TAY
gvL2lQ+gYlJkO/5UjLXlEDhhTzxBTDlilXp9sD1hOsDSzsX+QRkU3pruUr5rjq6kToH+WbKnD2pO
0Mu3zrdDQXZKHRbp0/8rViNi4FkOr76agfGhCsFBboKnuWSnq8OTFDFeBlGRpcRbTaOseu2OvdkZ
V+XnVElniLd4ARvc6Lr8Pcoa1tzV25+7lfYZX49yPHQWgMV0B+Dj1AlEr8Tt8KkVUfSw03SU46ha
xP4QzvBByY0dtVXJqj0kGOVvTnTU8ciJsOFgbQOtNV3HQL60QzG/23odJT93bxTaCh71+NX8e24l
0MfmtiPTnYlAlEunsvQSyMn/VYIa5dqwTM/EOzX9Jao3tmtYvMSoP1ssi57ro1dCyL6IEj4tT8D7
4qCpd2yepI+ecu59bnH8qjVWCfq/bIrEFv9AIwjRV5rMferA1I2m6Jerpc43cIo1bOofPC6xLzSW
/XRXpEewYeKT1s1rPShPMJKKfRXQhTxxG9txb6BbSnwedTSALK7rQ7l6QiSuTBdDpsAvRQiRKmWL
dmaIBIUnsAzJrOsFJuRbHuWvImi/T4029nRNkP+G5pli36LX7aeBl3flOOy02ZLPlCPExe8lZk5x
93Dx55BsjWY1GwOxzTMnOatfPzvna8KMvlHKJfqEKGQXimjT4EgFaUZPnfMVd6jGnhb05Y37iTmG
suhCJOYohXii3Oml64xPvp+9P63L/MCtpViAIBNOo7HiHW+S6JPX743swveCgvikouW0ei5Lo9O5
XH0GHGXa5WOE5BrGjEpd0USQgp/U8sga78HS1cWD/WEhVE2R8Uso2ksOlxuyk6yNaau58UhWFusB
DpHih/Q14oMdWcvh+g4e4Dyak0z6VrsHABIawLxFVgRMNwGt8RT3ayoY2nsKN7EesbEdWgUGGrtf
4ELQFP8/cLFqJQhealFuYOBxurLyDfUe4+dFKIdL+CHy89G3nS4D7jsp1DMCb97rk9rDv4Ai1Xlz
wlBAamDLunmA7Fmn+8ukkhfWlvhz6WQLdFHvi6KT6cYDlVeOe8D7+5aLi2xRiecYRfa9LSMFfo9+
HAzWNzVCEvhm25vDNxqXacXA9OZu7FOFARGj7O2ROVLQ8Tdt529QtJ1G7mjwinG4moCAVPainH4r
nd+T2RLx/A8JpwGR0RECMh26tP9ChIj2UMCtZCZVEl3DEZA5PVMe+wfB2G5pVwwMC3WfyJXwOXt5
vP76yvKBCz8iyXzOstZRu2hfTP/tI81FSBGCkNWlKG8ASCljYM4ul3pDobjxusMWbp8amQHkSrTy
0ol5e6q1ufdGtoQxJOR5WwWhrS6J1+MabRVvK/qYZUO6o5J43dueIf0qZBB8pBMYzPvuEswqh8Eo
wy4fT+lnVSK5pr80gmIckpfHZE+WR89PcTQUtTI/+OHU+PczwYB3EJcV3NixxvWQWHXr9HEiK+rC
SZHU55UTCS4WTZ1H5WsxC2k1kk3OPoEbyLZ6ANAJxldESlXsHq0sKHRBAOZ6Kwb0VWKtt84YQ8OT
gxSdnm/J6uy09qoYrMKumI/rBF5XDA8WkE7FyE6YlAdPBpSPiaeUTruDeHWbOtZqG60b3Ees9rNF
+gazp5AdWRgRv2x2+q1lZ1gIw83947hLKxPP9e+lAc1PGnwE7S93lKYdbY6XGZTg0i7u776oyAoy
7ZVrPGmfT3kt33jR8MTYFDaFdwXzyhSG5a9Yl1tDzgxhKveIHfCt9voy1VG9U117RA0bYaxCgiOU
VNgn4tuOB4r/5PGZB/F/4HwMD563t5uEbZMZRroQoPmUvRjg1pQDMRZXfDzhslVoa9PCBAoMODpo
LKFQ6dAKuMy0/qOTqklSEFpb6hx/NHp3ZOAw1Vkw4suhBJDEgH7dR5vuEZX4E2hrMK8oj3FTEkUt
HTiYqzm2bg9/6fajdzS1s1TAwS2/6QZIQKwQc1ssH9NLxqBSQEfiQI9nVecBHweYNxpOVoarNYck
eRUrvcdsLbBzhxkzI/KZR6vexSgm4O6E+pkl3jibbpn4/mHAJ0M3KfOIWLGBGWMwcaOnTT1+eMXI
4fVoi1t3YjxgpHCyo6v7iDugcIOamRR058fNEMtDH31ejCV/+RdeyV4TX2wGjmsHK5knSM9EfJjr
FYjkejWXHONv2XyKdPue9/n6nN7GvhdjAcksjHqzKmnJRIVqmXBeYBgX+wzSHF+LerS42eauNaZv
uvX3xP1+Lxe6kIZ8ojLttyGt+ETNUdZBq81/i5Is3JLny8XY9gjNFNpyv32GBEXReIlp+M7kJpMe
9B++FcuKaj6RTuKOqEb1GLvVuA4S3f9/P8IxarUMdMpDiuO3bUzsINYhW+xGhIX+FsHLwkWXUmvL
4Qa/coAPiBkQFUpr0evZlw59OmXpImeU3KcC8rXd6/FrOpgOn+EVOty9cdeZ94ZeNYMP/A7uVKnn
NHEsU6WcUKdwwhD6DaV3eW+9aidejLJdGhyAJ1EKH8/lZ+HPgsDc1WhZwoUuPjxUZCpOAIoBiBqu
WWX6/ty06pCZaIxKWJyoVuPK/cF1Jn6orlMga0IiAp+KKGK9yaY+1rxg+UEiZSo3Qm4HXHWBOGcz
THB0eN4ag1lpX8qDib013bAQQ14PHbCsRLSPyZVvXhvqRhcP/gKd/LrYX1okBZdKZ8EmcWDJCAss
JiF4QvpXuU2Uwv4dtxV53SuUtiytazm05q33+4fTG0RjEBoutmiBfBoMyKZy6YpG6j+nLDzAhVQu
jo76unfHi+VObjaj8NgtBNzxgywbYoPpevfEX5sQ38NJzShTcBa60prtc3rtF9PEmyaPHT7rR6lh
jRg4We3tTqAYVpMqueWaZTQMvClsDgDKA/12nGh1/QNvuhZMEhLIpyUIpcnCw1vVpWg/AzdTAWUd
0QCzQqxfc1gK5ouVR67pp113aVD2adNV5hv+sxi8+zuuErvNJRKyMdAZ8cORFfJ+/xNQJcvLtOnt
TkPoh7gWZiPMDWKEPwc9ukxdL9BPdGvW9QEDqA095wWFxF11fH3iAiOZysT/Ue19o12FAIhWN9+E
BdrOYOc10rSi735Z76fvtsI5aZOSJdqmZQhIrfRt35i+R74xW55ONScU+72t2ZDI6N1ckdgv+fF7
9INB+DdoDubBUQde6D2zlaljzNMKtY7yjFbVnGEB39VUEMs3fuQRY0IRptoNfoyoGJ5MD3WZXBDa
eHwrr7W6Sj9m96Xv6GO8d0f+RBPktrkIV+1RjR0IgEroP9Y2IvTEO7cwm2Yg6wbwxLams9wHeXoW
BDvo1NyCddlYVrn/Ovhtg941sESCJA4XIRuZwBymEhta0dCVwtVWSpJxa+m7v1Ks+Ilp4X/6+R5k
T+p+daXSWv+OTHk4duDVoRJaK6B4qpsaStZ8fj4wBPi/FhdtxLpJf/TvyOvd6xEKZZPd6JjUYTCH
LG3fEq4RTNx2sDei3girGOitPm18PgC/qhm9cXLYaIf+ZFuAYkbx5dVqs1aeqXskg4aZfyh+G0ed
gZbtpyAse8foV+ntT3UnnAS02c7YKRNDN2QVlZ5hR/EOgG0tVThtgIiY0XV1xsDHu+NaKnk9U2DH
6rkb3iRbsjovcwLF4U4tUNKjDNZOGWIimsu1prU5VwTPbf2I071fc54E0BbAcVExoJmXLBf3QmLF
yCXA5zuOb9+ZCjFz0KTojI3BGNDs2MtaEnYvIqLnLasSY8QG3kRuNFfp6TsecK8DNZcC/pkP2PWG
IYBJ6g3W6IEg38Ghh3+RdztZUx9p0z3JQQqZ1Ykx9xZwgFLFA9i2URCz0g+Xil1JAR72DGuVICKi
orCbCwPDO8oR3X1piYeVCxQjkvt4DCwmu4Ag53X2Jpkd5DneitWqlOPNDef/o/V3QpANwq2ipqdu
pTKsG/wC94O1hrhxbMhMizFhWxO/+KE4ywCEC5hPn/O9HZaXIoEGfP1qL2WXM9+dLHXLW4yWZpAu
PywsUDBv3VfCfGuiEy5/gBpsqCizB7bDtot7xBFMuq9SnQy+xeATebwqFG9eA+vMh9G8fU+xwXks
j8DM/IbQLwgJdIXEDUSQ4BFhC28mXUX3fJOdzvrfV1fJSxAeXe2KbYfCUXAoGerAH/wpYls+4J2m
hUUqdMybI4Y6TPk0NtatwIwo88qhnNoNOIeX0n/Ui88WJ35FRdgVbfdzV3crLGEvgvHSt+OVWsMB
FgjBGTdaqq6PBv5vV0z3Kg2xt6ixSak19/QMCsuQnbZ3/r8wdUQdhnwlrtmJrptYW3Lkf5pw5BOE
shLHQZgr1M+kAlbNPub3M7jHwR3EbBnAuXoBMr+gaOij2mXC3UIlLAWMwvGgj+0svo75spRvfTpE
hAM1Wa1RWaDRJawANe4Wh6fTo3UcxmLvDIHQj1QXZOn1RgefkUTpF/uM5Zv/8ojnMIpZz/7Cwx73
hujqLIiAjcWO5t4vYd0vwhhde7u+HW2eA+NFH70HFSt7lB+0Ofd83rysuazecGdEm2hrI80dJZai
eIaZpKh26nJhgd0EmDP2YMOz9uqfekNwptGkwoY7ieYifvqmElolXjaQUkz5xCEgGHst20PA24PI
hBk1I1AGGey26ta5av7H9P0RUGRMIKESi0R9L8Psas8WUs4hZIdO96n2knlMk8CWOR5zk30wyk45
uYmtHCp2Xuu3/c3KmDlaLUfBpuqfuDBvsok643BR1gwsqJc139rAxydCe4cRjnXmERpwvK+OZvAG
uubZTJhRbf/7LHLJlfmfwKLsMzVYb84BUg8o+ExASbJsz9BDTfRjBaNlP9C5Vxc5B88x+D8BQ1yg
GQUAPF2e6+PGYk1vJDhqlzqA5XePbSgXyYpIk77OugcCqMrvCs2cwFazNw4iNSmxo2mu2Qi/AkYW
chCtt/Dl014Y+vGVFe6/x9hGy5g7shW9kZZeqXo3soH6I7oSI4kIhQVQqxKtfvXVpJdk+bjeNAf2
+nMNIZIiPXLaFeMsfPMNK90PH0TASjxbG1YUuAjOqvQTjtHzzTf7H2My7H34s5ITEkABb2c+ey2S
Zz2OShqlJcTNe3u0ifQD8CM0044MWh/oGITvH0cTMgeiuCYRbF0keSf1e41tKLxZ9aADLQ4nf73H
R3H14GuTgjD+f3r4hTgcqc6la+dfSnWTJkMCfZ+CHepu+ylkxv8dYWSsiWAIRl6EK9/GyMjwywzW
vHMBZq+8S/hLGmIQY+wieEC6078NWPYqa/nSuTaV/VWwpxRl8qzp07gdq2/B+/SDEYKjrwxiVfNc
OrwN3XZPRTHN1Fxl1WgTAmNyRwt7a4Y2ALjfJMTx7IxakVEx47aHOtxr0j6SYpY4Mfuea9LJTHAZ
JyZuKrWepvjKhf65Ucc8MWonmVTdwAHHVN1oIoHceq9RKCUztpP0gr93Q3mpuOdUcQUalL1wRyN8
4Hg4VQj3PQZqLf6sGHtUWGERxpxmAj4Cr3+lZN8h0V+dPcZSt1ST0FkPhlPRmvNR+e4Bvdt1G0tl
eS9lUj0Xr1jBhlzhgp/p5Apmvuhf5RSCUpEj4z69nT3hRW0MmxaozrV67LY0GNc0XZvmnSxZFLRs
pcZzgQR+2Bwm+RIWpgDpShW0BIOlno+Z2dMVckcnRRnVueFv3ja0wjMisdDE5tlr3DZgzAgqw2uH
f0oCpSNGolt8MwfSytUdhl8CdAEB3f0Ni19vhnB+sdwone0ec+Ph7OdRTj9zmO8tKD4/h9L1n/lX
2205gJ1BJLOTRN76Y5CfQkKXivP+Xfwv4DeeCyvNkE2maedWEKPxcEZ/km80dUASK5Tn5wOU0Co8
4rodfYE4B/UeiNetG5oR5JGsN/B3nyd+ecD5Fd9yy3d8ilgVmxObsxiRMYrbB2jarWxrgKZoTp9z
ftbtMv6eRtW6FWUzYNI/o+09IIaBqTZ6+Iu0t3C94Vs3DE/vGUV1UpWEiAHi5gaAjl2zcbJ6etJU
nBKbKKPC30nkiRTz3WJlvi/b+pDjY+r/Xsc1KFS+1mvrHKrvCBzvXm3VktK5Y++9czygBapKt4f2
8hxsVsbUV3+EwgCpUvme/LuuU6X63Oao9ikWsMPhqHaDG0w3/EbpgEFtteR1WFwojW/oFKpG7fLF
9KnHsojDZewdvwfpGr9LisVQcord5mVDiRpTZBETMCSdROQGCLuaSkl2HRht1CRhfuBOGTQYGqqm
KE1mbCl+3PINJ4gjEWA2oWHPjZ/PZkFgHb2+7UrJiF4lDkV+Hv9niyohrMK6OPVSvOPAQtWZNLaT
EEjxlwlYNo2bGg/9dXl62yL3lYdCfhRGgf3GqdPQac5dDB95afpBslrQ+qyfVFcUGz0G4aTzB/p3
zEAMsdR/vDhijJBH2daoiO3N/7nVrnQOiPp1i8k7GgOXT7urfllBzNnFuH5V0y2AL7+gS8KBu0aw
DYi1jjO5zrbUUphccqDDGx9clP7m+v7a82LUU08tkkBEIoOZciDQa4AbtCEtjCOCxDNOSuIJOy3k
ufS65ZX4zeFs+y/9O54noZikeY/U6IBXCP4Aie6dhPuiRZz2OvLQ7o8RZYligAm8Q95dsc9xzSO9
mjEhyFCBbgJDwt7VNCoAlONBPbVLqjFj56sOS+BaMGe0Vr0cPvpHaIoUb1V7Uar/ko5yLg2uENpy
r4pqeJvDyEUHOvx3VKFXd0UOpGGvUxzH3eObxM0R2nVRP2BvKije6OF/wuKuArAAM8zCLRdVgkWk
xDHyO+YxJWPcaq4SQdVvoTXhZeybbxqPWh9mWH3YIwYJrKCgtLVlL+XebuckCK8u2bt7smGC3e94
jk80pBqK+GEMHdgavbgsVzlkwYdtb/ywqH6lttVXxJ4gXqBIhoeU3TPpevPP+UFa6sAPfJoT9CdC
loRt8q5+aaMk9papDmqQ3bRve9BdZA44QfUxjv1TrgwbuGoK06zRsDUdd0dp1VUe2lBwvwy1TGsC
02XM4dtmMkEP4p+9BN4J2TiNhQ0C4rYg4krjh2PNDse3koANSrdXsc30iLYX0iBBP5lXkpRhjd2j
77PpPdPVgTnuleRgdKTRmPX7cCDwjvNOk8HVsAVLq9mWxBjjnUtDCkI2JNI49/my+WyCQNsCZ6VG
RkV0cB0P2zeiUZQjNvwdXLaoxm1DPdSIWN4odcoxm5+1Aa0W+aVPC/At6fxmwVe7w6c0ZIAB31lC
ax3BKJGHpDHrGArX3l5Z7YYGuWTbATreN8bbNMjMzbSzeABN5JdL+uaBprZ91o06+A4lUyCzFWoc
T7ftr0jmLHa0upZXHJOZxAO10qIuvl81+GDRJgHe8oJ2urGSo3D0ctEUnpwWJIOrVbck+NoONUSE
kcdYzXamOWMZCoKvLeI+PdxAAXZVAvSX9rQmk9FyoCQEOLzki7q7UyfOgQ8MfFVDlUiihoABXE4R
BRftHg6yEKDGYlnJPhqHttNmnSZgtK3lWflgmHilft8IGoAlS+NCqo8ccu+hp6P0Ps7+8pnsevdT
703oYRmX/AanpGIeiyOHznjAu14Mt8HQQrxbzmTBSoQDpN4G6HUo6W1a4x7o9lsBxOhvav1prMrs
i/KG6AmgY5bO44vhQxEiq5JFdOqtyjEIGMlQSQEIUoiVfv3NQ5Lgn6oj9zjHh1/+rm1MkeB248nJ
dXGU4czRQ1mAtlQG1g6b2ulNbj27ODtWWlgc+axtfqDYFsRo4wdSMASQBOifXhf9nSKVWTcCu1fm
stWsesdsR1TGBK4PcPqg117wpajyxYL19W6e5ivOEJ39iEtbv9AE1TRSAl+vWx62E+3u8Nb4gsHR
FVT21U+y8l5VCQhIIlNf8uuOhvbaeQg/uRfcIZIgkgGZ7AKpWB2qK2QNVT+gzo56L+Kuf5YJmGJG
7zpGduDEO1omQxsY+KwELw4DKdzFBnzmclAQ2jW4d5VXpdMNpOB6uEwJ7RDq9X9xKejMHLiOij1X
D6hI863wKOaNqsBm6Gk2m9WqJLdJy7x58U2CNuDXEKos4T4Nhb3BS45FrFYcrn01xz0ousBZtvmv
SCFatUiy4zUFDT6ju9u+LGCBg9Y35ggOn7+wsgJTujLn/nBOhXcUm6bl2l3MijZg8W5NEcGzV7ak
jhB+U/x+L1pISvrwbnsOphBLN3LhK/j0hMbbOVDtokvwX3NNHGungOoWEWVTikZWTFq4+7gt48G7
cOSEF2wgfgN6FMVk5fUbqWq3nYRxIdlIa2hB0eJ08mB99N1gz+dKvUnh4s4AuXlp933kxpdyR8fN
7fMz8W+LadvOPHwHrx+nA28l27tB+K1ZilukPZhfbbB68hTiFHe3IyKDG8QHvK+F54vqgL5C7s3F
D+ZfYJiYgayftrAU1ruZQuhkXM8a4PAyBJ4b3p1+ts+KQrOF7/vb5CI2BQwR7ir7zPJnGTOuPJ45
3w1sFvV+qWNRpkjaBIfJ/bKj39t/O3wpDpbcsR/QSO7LJLEsEeVIGeLK+hzmB7MrLX/EJ4+Qmn2G
Sj5m9rHmyCXm4TSkq+WvBPK14tfI0fNOnMgW6hIq5V4ECA6yc46jpvICpNxUXOXRwvCkSwf5LHjZ
H9gkz1+bvJOTdCcXDPra0YCwWN1EUvxlYfuOyPIJcKcJ4PveYLF9NKGFXk7NM6xXvGIBtLpp35fs
m/diQkadi2GhvWbyQExrvmUgeo3XtKAclXTWexw0j2NzPzL0O7e1lCXnpEBrEI6CV38O6ha85x+l
Px5q8qV9aq/8lTPShgEQljPiDQphF9+hLtPSAQyw9HjuDW0xshHuS6XTVWHreXd9/GUodQIyoUtV
qK3VFf2l/ntgjza9+vipXuxY+wA5M+IaTvosAfTDWKjnwwi3XhO+RoeWuTGgJS04fPxN5yhWUmWo
4CVNCvM9NrbBd18bzjg4W9CbxI0vyHJ4iIDZkjBs04q7q1GVrV/FXmNslIW37+clhs5u4sLaXxR/
FRH9EBMAa9WtfAdU3FVtbsEGTXf+Q5kg0lfzV6MNRTOS9ZGW0PFS37iA8EO/WtVvur1DW9kTl/hi
y4g91WSht0NVLId1OrX9e7ZVU6TEiqVqbsxlD5Ce14dR0LpXoSM6jEL0qtnB3V7DkmHHgYyQMUN0
N+xtkRb0n2g1v72ORYDT1btvtXcZ1ttzhN/d5Mm2k5EX/RbYHyOVW2GIPpBq28q3lrG/VUqLfhmY
pEbEeAwzD7zSkQ9W22lW9jYSbUUkYP3/nreU7hhQRdRCMVTEZRZjtQ8eUPm6FIHtlgy0ozyUcGoE
fsXOPu2eGiBqNEhFJg2yaO5hdf9VAWECafP1gbeSXcy1UDo47p7V5x8B9EEjgd2BHP7dQGbWnnso
WxtC9lAZCRrlSGRvRsvFWEnbpXKExSXWa9R87+7K+f1XsMxHq+/juL0bzFG2asvNnN0QHoO355zS
SCtYy534AU0wn4qgTsz8TaP2KGe24//EanCCN06XQajY0IyTji6k1Q3WWKLk1GVw4xpfuY893/dl
4ycHNB72vzW070S197aF2Grp966wMz3ickiwoCzWkWaLCyMcWBH0QKRrHNK3TN++ElHSm9z0PBqW
xkPaff84XsVEPxYHdoK3q7KwRMj/nYMICdbTogNwXKvY6pGMdY2qCeChdiWzK1gZxHKLAK4Ff331
NayE3LZv/+tCkZG9HoKWp+qbh8UqJ186ts05Gen/AJZSeaL9leEfK0QlQG4Vo+HhojbKCjsVBYtH
he7cXu2sHZq7bAmN/a9SgBRXhANcSQ8wkQX0iz+8hUgdnxvs0L/Q4bgTgCD89sDxnnzssh1aKElL
C6bYkT9GXWKvFi0eE9awLN64qWnaMTKHCMEV6eEc6CvXcRiF+qIt5RbODAZ3VnecmRvXaf4kG18h
GmnjbXA8j3tDdWZ3ZY5ixv0tareXlZyVVBCEWQRIo9iU3wnunbH+FEtV91YRtpIS/p0cA2lTwOIw
rni4jqDZT8fMPlSrEBYTifhYkZG378WUg1CSGGg5qGce2xcJtQpPjGpPMubuqK4DGQJVamsPgWGr
UQd9tqxQ3k91NO9WnnfB9eXAxkp7ydtA6rRWyOxbBxCquymvRVJVwEDjZ3/VEkaC+FOXKqf6kfVi
Zczcsg7bTob9q86JO/r8NkNSIHlUTwLGYVfsBcV/1Aj0jEAaeSM+XFfhxgHB3rasS7qAwCROozpY
U8NyxEgnGydU0+abGC2MDy1cvrpwx5AVwYXmXQ4c22omkppiRvo/SBs3oVNvT736OnuxMa8pDqLl
Jk6iHl+FbnYv2eoqPTQ2BiMybdQ0iS//S/uFJdcCCDSc6/tSMZe8S0GKCLP8jsv+U6JpMmJYyynV
4nI8RicTbF78MhTlfTQw44A2Py8hFoCdCf1pJQkuVBONVvEJ6JdEE2+pJ/g9+i4vkzBIVaiQ0leH
dMvfZeOlX4hYTjNEJAPAz5KDTcJFGGe/ix6w3dDmzFQt34vG+24ommqnBG3yzHvw1dEgf+h7duZX
s1Uxtrmx/MHd7ftLtm5gN6yS4Lgqdecj1I6JMM71fm33mlYA/nQh5iUpZkno5j2cjS1IJt2tJfxL
wZF0WwjVvK5+WHjv7W3s1wkAusAgdXu/wYiSIm6R2e6Mn4YIPzSztOHlru7vjE3Knahvgtljgs/1
zPG45qBfSuq4y2hvQrI/TzCt1v8pccn/xj0+Nmk5j9IuTBAjerjScuG81C/bRl+jdHmfKQgWaVKc
RisIQOij21Pj1d1ZApoNWv9vISsVwdQjsTwIhP3+FKIS8likfjNDk/Z4ChjkBEcmcVoVNN0Vv0S4
mC24iMFKQ2RjKC+l9raRfAZYuSqcszYgv/XD2RkAQ5Lb7reuU2nWgYqWEq72BbMgrHJzltKt2np9
RcnEO7VkPxNqN4MX6q68KUUhiKHOs2cLc3oMVrpp0xOva74O5v2bsc3DErkoJ8BrHybBWMlRqRRr
51uNGV+pypCoL7raPRGqrXt7dllOmTsMMdoO1A0QFgLMWE6X+8BGqZtQTT4DFz8zHowCBVUziNTD
TY0OdVU4cLRPG43apTBQ4l0Hkiua5p3GnjCcfc6hHl/0GQ7jMPIKdMiAGcL4F8x0TAsnIB9/uG9W
F6QxDs6LmUlBrSfNSaY+7+OjsoeFDaIGjz9JtwzecBJRdvtAPCUdZG0EeQ5uDI3AwEtYgIkBAN1w
UMjDIyyTeYQWvFdz+WSuI9UnZaHudlbygvztcbrJdedo6rPdstjZuRm3U5fgg/aYK9J8/JNNL3m9
J+1qDzy1iCLXJhoAztAlG3xX1ejflV5xRAzoasVot/KDtRtoNb5hfjhR/GEeRR4VHLUpRYaFj/fb
jyNWHrvYgFGJFzh043DhmKuCbzcFunF7PtrMUZPtVm/nf9aPTwdNGmPx5x5pdcppk0HHeiaE0GP4
0ukppLUn+eHujnLZYPTUtXKaOENLlZ9MamUhx7K/kvwGzkAyDEFHcQJkvMo+Svx/Tu67EzMNnEQ2
E5ZmTYMMFss5OX53tLtKKhNe0p2CZaZ5zHoYAuuKiXmg2F6FJc94cK3QAUduDM3paDyCYHG1yPUJ
NDT8rDI2XXbGYQLc9W1ng3i16mz7mWvS/ZAMgipk/1nM+Hg75J/78135+yJg1wpnmgksNIEvefHj
nXriak4GFFCQdH7nCIEVi3na3ukSEuqon8pIHnhrUtcSgdKW8pwnQUgeLO4zJobJ7mlRT2q9pJgx
fSB8rxmEtQE7H3sx6C+onVD2d6+TcAXYhe9NpbNth44r3AV+u4gl5qC+ex28OAV6Gfn6aEWmluTg
j7NYGKop0G+qgwPbfXFpM1wRV0ALExXWkyTd8JG+HGRJj3CUMAJ4aFszkdeikG4S7mGeyjhIRmVa
sTJjhjC5fMQxQLfmKxUmJEIt8/LZEB2IS+QkKTEiBPzN3NBqC6DmehyPhZMGav17o37ejBmO/v2P
AgVJ3X/olDQ0pkHoxn2CvYrmytHJn51ctVJgHK6uLEV+khJHWBeQnznzyeEmyLMOQDFYVvwMImbE
rfkCORvJVXdFyyZUMzEmQDzk7Jp2Ha/AVbd5Fts6qJy/UgS7noN4RRVG5ylttIIIo8pJjIlyak6n
V8MPCWvjLjcQS41qh6184Y0fazLK3ubedmc+c5s8ckEBc+kQ0oG1L675zE9+7KpTrfpfM6CykI2K
9cJ6UwM232nmWj184ZH3JVkNYkpaVUGB09GqfYmuReT6BnCuOiVHWc6RRFbnSNmXFVtVCF7JSwdG
kKJxmcgPzSJCP74E65d2ThFRa4mdy5RBohs5N7ak+eq3l1Ll6rE5v/SV9QFEI3LrKT7nhmm6HezK
4vdUHOhdhLqiYCuJB+NE2yGFoowaOdVVrjFwIdl2LOny14B0hnlcBq1W4Zv/nIj1ER6OXk5DM2YN
PR7pNHb6dTOATUcJNfeI93YuRCgwG04uSXWGjs96uKTnNQ0n/PnTpgD/Z5IyCxiFJkkuWQkL8xWK
D04hP0x4F4HI7yzNpY5XfJFYvCRAvSPJM27X5jdqGY0CVO26D71V+EnFaBEgWYjYQ56v8npMSpWh
32fdKbNE/JDfiiOPrD2JWPCcFP4I0f/DcxVFVZT98u+G7h1eX8E1YJ30aiqgMCKKADVbAV0kDUUg
0O9Xgo8ywAKgceQ/K4Bbl0SkQ0ljWVBjfa8Wf9bEDgbfnc9WTVeiMUWsoZEx57p+gyyytYWx2dBA
PTilY23RaC43AooDV5cUy1uL9Px4TwQf8+jbxOxGMdSXUiO5xOX3tAbIrlOwni1LLwjWpY9nEggV
wwxHvGkWG3NgWKCuWQUS+AEMIuUAIq5xxr5rkiacOJX9sMRQW2QonvS+TTRqq4/LfFgeeI62fSKv
YmwKE625ziwwck8fWMahN927zASIF5FW9TcQtoEFmZ5yx1o9JkY9a5Y5h3nuiKHqp1OEApP/BEEt
bJ56R4jtKGaZPP1clFpQ6nDSukwOQb7UMmvyykT34FfTSI2B144WKuas5t0FTg6N9Jq7odGxd+n9
5JMiYLv3PVE+4hydo4dokyYgAF/mgjHSH9wz6ZCHnzbRqz3hCqXpmrBrqK9IvAx0nl1s1bELjtE0
zrkpq9QA+jrcPud7P5udpLeENdhp2bicOVj3zZ6FAdrMHEqxDAB31uRnqyaMuVvQGLLMsReO0fIu
Wt5KsUk5XlWblkPpZVodPPH0ehfEoBMHKu71J7t9BC4872oauAH7yWyESojxB3pb0Jaktelpzlz/
Nh4G5K9q/KzcnwXHyV98JM00IzbawNAOQOiolfCQfHV+mOFWeihm1aHkKAg31577oKLr1+AeC4do
hXlfrJA+tUYi/0cv961gocGR0JdgJ4PAEHAhIz+VAZhcadw7SKdnZD6qbdwpKYI2zuklDW5EfggC
rPkxBwZKR5jA9u32yo1Eg9lTAYqY7GoZrbjCq5gICye8VfMTUnw2wDQQAD7hRkIKZ5HLfSXvJq/O
KsfLDXa1LNiZob4IcjxwXUGOZSRV4LbGIAgdk5LIAxkvYlGZrsru6RKtPLRC+OjVeqkTSIhzlV7w
CIcyZFINjd4IupIsVWltfEW2dGadcy7x94sRcdxQ8QvOXU81vDAm+rTKAunl+YpMQZ3cHQoKWVqc
mT7MdAsy6+71xDoPqnjN5x2bMQEELGOWVzEJ12knDZrMj0do67V+OR7mP6qm9ciYHfcMl65lrCBY
ZwLAqtu8oq4PopIH1T8JfLwydPlzEmgZjcRUZawNHpQ9lySZuxy6B/YwZKOnjwvHOT3XqGxSyut7
K8jCKDdR473sFuuCmyIsFx85GV24xxwd707TPjg51ZYg0pEIUmcvBq9iD1QFuN/6FOTvIv44z9fy
MlW6VV5b1iV2YF8CMu++2OoA4GXpvfrs7TqqMoD9DX3Th5al22Lt1etkM95geItlD2fipUgM9715
LOsoW0vO8nt1qh3DrF8RGcbO8nCmvwBt+S4RvDjTDKWDVu5eaE/tXwGt7BQETT5XG2A7quxrziUr
CBfLt6eH0aYsur52HAAEve6cqG45dCvZtOeazxboRi6+QE0g1lB2UepahuZfmLC3fe9s9xseJnSr
jKactNQhxFkq5w2qOdB9SmDRWjP9M/WbzPLX2CF01PbUimE0y/qEAVZjWcZctPI2qbmWUxH86MD1
zhtLH1V/0z/M3rRkLbMKU6jM6fKqGHgF/jIjD1HVxg6ZDSWK7algRudGjNg0b6kLLEG31aTvOKPB
F5MU5GAOmDGsQQArKGTy8lvr3F3pTpP57QPOn/N12qFwpr1KhlTHaUkT7FylO3WX3BDx7MuRdS/F
2mBDL59+RMyI1zkTuMMhbS7uPC5YVIAm9cXzs4WBGh7CuCUHmzf9Quee+T+tkUf7n/dWIUst/fkk
oUx0/7xKc9hR+2LRWzbjE7jKvzR7k5MaDmPyHd8ekaHMXmFbbIaclbNsq/np+deHCdTh2QewRF/5
SP81h7ZXpMvLvA59FkR0lGMO2SXXwcDTGLYNa1FDq5UrfrKwbsMIpS0TZ3LNRGPgMxE9z6z8iXRY
eJygDxOYQzHnA3//mqnYMsRtlKxme+FrxW6R83ZyVHIY/2o7ZXqxJ4D8HZ2Bs2JcssgTHfV3tU1J
INY3otNbkII3trAQmvsNQOMexnws80bQJS7kFXWB4QcxGkqemd12q07bCdtxtAK59/n6wklpo3fg
6XOig+doVKausl8f028WaDqp5BFzDy7TrEFAlepxAWcWqRNHV8vJ8rUCRua64AtAokuYXcgmZg84
Uo+VW9kUFj4JmopojlQYd+kufDCVyN/2xFgsJQDry9p4mLuxCr1B7c0yMqFru8e7FkUMaVz1cAhm
yGh+MtY5eG8Q9b42di8C6aLvk74iiXXVi0BvzHU+9qnJcJ3hZtnNH+KB8h/B97mhh17yu3X3NWKp
91jX9tS851eNR05OopF5tV4E71cB8BTtT+qYUyNKiMkKgkWR7cH+B1qnlBDUASgna2NB5bX65j9E
WsQ9BEvpdzoEhiinSz6U3++sbrqKtzkOuXIOqi0h/WcesP0FcYvHQ+LOBtw0CHuxF6xje7wj1QUT
6vksMLkZFKi8cPASyurWQbs6fwQ8SQ6KrYG5HS3QBbR1QnVpJi6xvZlrSmxis8kpCMM1DgQtx5zQ
wv5venSIUj2rZZ2RfkSCCIEir4owdSqPsAbV+PKViXHQZYGBMZDCDFYEx1WSVVY+whsqJIL+RThK
mo2XrQr+cjFcyKMY39vkNAfBp5h24zzCESH/2KOjBcaQwC/O2FZi1cwTFRb4rBD6GL/J7de7fqKn
eTHmgvDPaNeE8iduPc9c6+wHB2IMqKMPIo946Ka+/NAi/qaEnshIUTQXq0S+DGsVL1g4ThKlnWqZ
bOOD6UjH8UtHE1SVqmf77LRnSPtEmXFZ2POyo0vLnbNacJCI1Jmy31UH8cxhNaJSMg+WjkO/NuG2
Lx6e8mudmVe9o2kx3PmmY7hDolVXJmfmVTcNF16xTdhGL6LgFC74lZREWHFhKjwWlg1wMmzMI8mz
FIr4sQHoe69HvGSNUjzSMlh0O0M0dHuDvhpbs1CiZpqalq0u0MiCddGHpa6iiLD5boGlqGfmR8Tn
oadiins9KG/hBk2/BozVdOCUzk3U03RBWP6HT2Bw1FDNgaChS+nEnB4/7XxSna1R96ObcZ2AjCws
DV5xPaLK6b3ermul8dVlfjTQlqQpqoSkXG6GvGd05+CHgXyezvrs4yT/ZQAc+V0sfyCTvoAeFXVx
Ixws/W+BoOdlez8D+tpDxfUdCbJAEfZf8oDvvs/ilweITzvCNGEU/9VE6L/XhdJrO9hG2gI6gZMR
RbZzlpNTxe8eFK/1BgcIjNAgkqT/LRYH0HeaLIk8vvpGSmI3DNtm0OhYPpMqkWQjFG9SxhHfduVS
3luXOGofvbTmg4tIx3kBAt+dHAR/njFcfwM9Zyrv3lF4YdYyE0QjahaX+Qdu8tdgo3O1zwpdLqTQ
w1sChKWo3WBRAA75/vAL4W2dL5gokJ2waAFWLCgEjzSrb9Rbrv1MeNHVf1EsPUZpiFd859OC/nAY
LPTy894g6oR9qOpbZvpeZpWIwkCmaqixTvrvcmd1mBAxNOCuqTF9DzTli1PrZbqACiYcMJhwzQ5c
yeHrFiUCZ6IOiWfkrfaU1/fN08WYYcNI/qlT7lFc0+RxUIVENw24NgsL80nGuwuDKBOQZ8zatT+A
NpML230UxG/Mw1r8prH6EvFowtSXIG8Hr0Hk+JccfPiv0gNkAetfqFVBr/ziJ64U76QS7cM0SD0a
ttLO5HQJtevA3jl/dSR87SZMmRvW/2lEXPTBVhcdVsE7NhaeAqj3qKKHjaLnDx9rWIIkWlvIRc7U
XPYV384BJHM8YqPyHnknjXf8OiCh244MtCZWW2w5RFSyrHDcyV2TtUfyc/+cIcTrU3m6EAhSJDFK
2Ccvs10RwlOvFHWOqe1BbEpy6Sq2PnwI1Tl1qVBzaZx3hJQAEUIrD5UhOffv5DCM/gM5p4FuDu/M
w+2FvMZUJZzpSE7pakvjUA1qXkvVKrJuUeF9nnnQX4Khq63j2coHvA/eQcQ/bAEO7xSDwnBxVqkV
spvJ02h6fzO+guL1/cBk02m2aT+32Krufr7KRy6mMRpxjK/HExgNSDLveHSHWT7C6yShHeqPkp17
etpjzC9za49rR1XN/leELFG580xzGlD7tUDHc2PggvCcBNM9l4bAepcNC5jopTVqtGmsZVUk6lVY
/80tZHIKguQbuCCXKV2vnTp8So4cHWtPxrZMglm/DMl+1l0PQbvJDlr575+N04jVLCtsSAEnpWrR
n/qNH5fqkIrirm3K/LZcUJPceIDLIClJxoWbzu7QJcaW6VDGftqB29vupe/zZ2P41bDW5Pq3Mw1q
5uZdhsouSGjxBcip3X6N7kqwcgTcTpPH8kHsee4UccJ7vP06RODoDEhhED+tkeQ/ecz20u9zq9G+
66jvHG+s+eLiLurngp03M5DiidWpiNQkkd70CXx7NqdCSx1jUovr5eTSKd/ck0XKaIwPJrR5KFTZ
cQLI2GOo0y3RyW1EL/gXhyrpeqT8KYlRy/YKVy3qmZMfDbcdaFilNLxSY7xHGXv5TxGSeMvTINZ0
2eECpwFi6Li/pa6/p9S7YqjMQgpsCOCJTp8EdM0u6PE5JnMnyarEbIZYfDMjxjCkgvBjFjs3EaCM
FgF1E6AMcXAaNtMEqbOhEkv4Wvf1RmLgyFPCtuVjzqtU5hV4Mmj7TIp2f6OQw3spUv3QJ7Vd7M4T
2LW49xk6gg5yHytH8g06XRfPQzJxp2nCK81cLS58Lv6nkmThIswR4E5CT/Zk++RMBtZfhPh5CaU/
vO87JkVUi2LI9dFPoezO1noAkYtKnCFAMVmvCewDoQSd5VRXrLul46zvobVjGCGMPAXhpO28gHac
1vHC6k/67asH7G/S9HQbZ8KwXG3M9TvhQUKWJ7/oOvCB91m5RY9+4xlpVBI8NU0HKybEY2Gpxiid
6inhCayGE9Co8NWG7YPRaplvxobJVJEF2pG3UlnFbVE6cXEqZ2WXhxHSs7k2CCiH0h2kh4U/wZ2i
xPUX+UbZ5g+xSko7hMsLj0Y2e91UI6V0gZUjwXX9YksfT1i8hj36g2l+uGCP+h0GyhZpcrYADzTV
T5xLSiiEHxe7Qc4c+5IiB5ntOyNItx2onoTtRilOJBaJ08pHXH9mawaGYsZkA8v1mq/9KxueHOq/
fDE35WDAHOz2mSScT9hekhBlb+0Hy9YWUtvH2y2A8xSx5gbnDnpTzaNXUg5Anbk2pch4TGWWyab5
SCUDaANayF1Te3jqKKu6xiuv2A1JQ1lyHxkSrJUCONkALT5LxnmVvE8a+9eOW0edHAHYFbMcXD1K
2m6YxA4W3dZq6OqcF0huWj/qd/kgbhQS5zWhfp+eMU+BRrd+7iWfVJrVxJ2JlZ3AG9/fdQOWm/F/
n/SAJokdA3e7TOupPCYAGZXWj3ogL3T/KW/kq2Hmi9RhgWqnv0xu64uhY4/pX02BB7g0YdDufpa3
2zEZdi0iz/uZxTTq6wA5Hh66iXl7vw54nGr0WJCxJ5L0llW5fOWUeXdV5xgFR4LxzhlG1TaFveIJ
4zoeoar+2h8w8LGbOkLnP5dlNCa9/ILXfPYomMD3u5eLLUWYKgofJg3orUmBHSvfo+P3DaEfNiwl
aMlkpjAw8djGbT8UcscC2bxKcxN4O1oiJk3LSCzAAGU4RjVktLutLUasd5bjR1leXMoIqZKZZnNK
Uu1xB/wtcxfnqHNzWYmlIqo0i3lwOnPhysAcH4FrlW6ZyyX/r5rwWwR4bQtByaZHwIXz/hgtZqjg
eOxAdiyKNknOugcHXAVf8kXtPF0wtSNI+Uu4uizU5oKI40bxwi37OkYH0bO1fAB04JWji5Aps1yY
JDAvYF2FeMyA5hSBTAIU2o8LETwcEAxmVbr65ttEu9ecFTTqOuQlUROG5blDGy8G77lDUGQJOODQ
vAWUvXy7DLyTXQVD7WKbWNi8TihskTzME3hVN/tnLh+53LgiiBgBJvC0DYQzU5FW76N3qEnb15Im
Z1KkU7TXRqHcdr8P+EwM9uPOlcdoE8AkPNkDC6DralNSw2fuN4y+7UgABFdlwXtC/rNGorYK06ke
JLVXG4hzDZBA8Pbre9Fs7ZbYJiJPHZsywmgb/zHeFyWH7NCQN15b/Y1sAm1gVwl51PD0gmH6Oyiq
NAIkUakynmsiXzzzYYGLq8jGarL9ElKVMdNPhDKYRWKncAGizkPVYMDkge42VX2ydwIbos+kUt1I
qM7GMZqgpdJN1WhN870zG1aClD2axlLWAR/KqHmAmAApM/DPDr/FF3Yxnb6DqHHmMZCFsiJPLJy9
0k2sRCkHUAuaEgrGPPdnCpu7gGfK8NrkLMThQnCBqqVsHi8FmHLi/s6nQiFSc8hdEleQCTJzW2VC
hRWEQ32Kz6MSxNJR9RXGAeKGA9auL76UNHBLxAvne/jITBxUVtsds0et2ZHKPiLB5bQLfNYx+OM8
mDxQcuh7VKsEr0gZlEgneiyNJPLPnLul2OARl1k8FlgRcfKhAEpZfL+yvfGi49d0hvneWfudFZqX
KPugToTcUPYveib9rBTm9cEGXRbXbnP54rknnpjo5ZZIb33RTA0F9mG5s9ZhMb8220WQ97t8f1Rp
DbUyiLqBwY3wThCYFLsTPjE4g5sDZRR6hm2oMoqrYkQzzBMQSiHLqzpfZoO8BE0qav0wrcwXqKsp
CQKv0vgz0UGxCdMMBc5Q4gncEHDimocSIsYZJBW1c6tavtkpfs535WsoV4lb29GEdmf621sc4dDn
mHRIoKEnQB05Ebqn+x+6IuUz48I38Fzo4naEQ8uBRv2kGhNtJFvNLWhsTD/Gu6Vf3TivpS9MtxAy
kqh4ffWWrKX+2JHvrXjpnGqUUDRdHR+iPyD8cyHFMMLAcvGYbbBR7JNOl8PTLHQhC1N9ISOc5IOf
b4pjS52cr6B0zRDQfZf/YhBixXnEhdOF4FfY0FgcSz9vZ5UD4InXvMwJ03KofofaLOk7R7LfJnWJ
9gY20A8vc0kbU/ZGfH7/U8T5FihzDUckyaOHj39HsPguFTXgGmIgy5DhbDI3kJhjm5XwTPv1ZcgZ
ZqRItx4CtLt7wmq3pRNZ5Ngy1wyzXDv8/fUbX2GmVtGL4gqmTxQS04lEFn+cQgkiLhdP/IJTJBMT
6iximU9kkRxlvP/qRtHMlCqGZ/hq+L41P8OoN6FnhGHrudCQw7qxSUrvnzFiZw6NlMVrxk3zcxXr
dPsM6UekEJIQqdd4fXfEr5d8qr6bf65hvyWXet8lf4DoRjk4LVgB4TTZxSaNR2nHgbxquBvmJHe4
t4jH+kFaXLQtDEPXHLxh9uMHuOOwuxPuekrctMwrJQFS929sD3buaDfO88BNIhNF3yC3NvnO5AfW
PWMuTUiOuY4qSOw2D07clqa/cd+yc1mw83v20UGOZTZM64qW16IdL6WXQ+MeQuCNpD2ntPsn7x6m
wIgiXPklxwSYh6FH/Qx7FM1+hr1JE3rDdL9+WeFw2B87OZj5Uu29jgWTlqcoDDZWyDfACIZymceJ
l7rom/5vIGoC3WQvHpEyc0h4V1iZtalMYlqQg/rdSkK3N2K758eP+7qJbqDZiLtgN0VfqkfXkm++
Ae2lHf8y+9QMz60MFTvVDvRafEgtSc3WB29qr1HJs6xpqCq+fMW6g6+5Bkl89kPBc0UTw5GqkSAz
BqcDVWRWS/lfE5bqBmKxxH4PaeKd+5MNkfYvJOpY9ZU74GE10zKiPA1/wcWk4sSktgAiCXvEOItH
PIP5yZBbC8+/btfSBdVEVzlIWQYFusnA0LU5RAIHP9GNDesv8d/A54O7Lj12Bc/pWKPK6gxuvFBi
cs6qcjiCH2bSSxUQvC5PRdqw9khsncHdUmHwYDSb8TVj/aK5/GAqc/uSl+EhR1WdgiMxMBTH6kEx
t97f4+ibAtJkZQjwx9LhC1snxHMBiSztVF9D8dTxXVaJyPLnwzqGmx+9U6XVBjtisfLtavTnKRF4
0HfB2xJY8brDHnV77Yb3i3kmBCoXKIIQTEoJVoj8DftSGWtudiGsNTDI9n6Uo8feC2kizVJPxV0H
zfXAZJSY07HfEs41n/MP0U5ovzQk1/JeWBR0nVSCynu+D5EIYM3lsPZ+6pbV2g8IsDHh0Ri8UjM+
noysCngdaoDqjPP3pbmlhcdqlMLjo/PQg2EeOU7MJiUvx93pNY67/T7V4+3eE6WS8EoxMbRhXwcq
AtmWPfrYwJkLj76XnVxL45dog8nGBv5g3uyjVsUQdJn0a1woVqoe91NAPh65wMDN04v3RXQKTB3f
73G2kC5OWV1xyW9WBga9RBGP4fds6iVJJ4VDp+eETlO/1RUTNTHT0fi3SJyizRp44qWpl5fjLec6
EbRDrRB2Fic2xArxlkf3hkM7YUSJ5EK81B1GQ/qYWCLWtVTZI1WYDrgtwIG3CdA/ekGYKRgyM/2u
RYd943RYoGpzKRsbzdl7tUdy/Q6UqHPp3UF7YXps02VAoa/1BmokllvyoA/vVk3xTsQVTjoS2GO+
6O8fi49CvhQJCrVradM/SIoQiq8dcT6Cf9n/1UcExceXOPZlrfLfxl1Ktafe4UMc7ZzMgfCrAEm+
E/e1pKkGFYHQ51CwzXOOZ8MPOpMxsbCCY2vGkN3UIKS2aeXYvzZJPbGGBqE0SqPLJqYbvyKvKvN7
r/oTQCjYtlX7YBDVs3WgBYamnibr1bKgAWSjdI9uBpXW08vFCFxEPNDcoXw0Iom65wNqyH886G5i
o7Ldo7ZY76AndDpFQJYJdxb0VH+4pSryPYQGlZkvFTkkrXT79i/lYwcweeJoplJTGUny/qVc+WPl
e6159tQs9sfWy7SaJqulkFjWCrHXkRxM50z22funKkRi2HBjbPV5JjIiKw96NWYKXTIdlckvMdcy
yjizHwDU7CNCPg4jCZ6pp/75cJ68myf1oxNLGMjGku5Gz1AXkee1iHdqC2MS8YYSeekcW8Svu03K
h5m23lFhpdfWoaDuI+Ik01+36F11nyw5t+T9hb7uPmL1PCm7z6a+Os1fDUz2JdICYTw+e9hm3N1E
DKn6sFwxQ4UZgW8UyhGw0GneEHQ1XxyR/iTBoFxH7jOohJIItm4F8NfSuCU+8ogjAJVyZxYHPzLG
mRIm8SOSeNobjDfRMJgNJgK/MWSZnhmUR2TYLPFu/Y+6DhwNgSTMhOl6HvvZkpvethPssfrOjoCT
WIfUaSSQaMOpnrJMf+0yo3mrP7lgu8rE+3GqJwk5f5Ig8CuBBkFNqJayQX/0Olt8R63PDajj5AmX
4jK3uGsdAZDDCGRO6jbj6brKzWrxf11ncV6LT0lOn0KY76qgdVlo7qTCiewhmQNBq79nDfj0f+lE
DREsSh0NpfuCQf4pw4TDpDA5m6o9e49ncCuK/hyDNqDM9qRmjZJooI9oLkGRPUdWHsqaiwYOMTD1
k8hOgU9py0MoYcip+Tc3AzN9piuKWeYgJ7IdFCfiIrXaxSTy/HGxFfK8WbGvesZMsnasw9Ptuild
4bBoDPMjd1tQVYaqm4iPGXTrle2Sa3mR4MY5T94XT+Xv1A9Z/RXldwqDodyHBcDmQ4cl52Ensp67
Acnl8OR6UFpM/fVCEz7Dvcto6xjpVtUjQ0MtN5jN1Scoaxpd6I5raWX7sB6hW022fWM4eJFXDt0N
rDN8DovJienWMKEhJtvd+ClMZhk1HTOev+v8ect0hBVHXFfBFKSaitnxN/33Qydd3zlXoGXGQG7v
770w1t/lzbqgckHsb2bdgnNjuy26RnhkSBWdXYX5Z+YbHzs3+QkSQqF4ohVoU3xd2INRqlw4XdaZ
Ae8J/CRPLFKJoMDdNpTTswYz8dz+nxELasDvEOTnJ9kO1GAc3zoxWl8DvUIqbQ7lIBowcUkqwnVP
rjiaZoGNM2FzDhy+O0Gn0QO/gM6kVwM/7Pp/2uGY39zbE2da4JwAPwYsdayq2IFyizL8ML1Ja9Ji
BBAbY13lu8okZbI64TOZI6LRun/x/uwZ9Gc1JA8u2JvPfjMdOGEsHRNPbFFZYr5+2nZ4eBnUMzAW
35rEwJCYZB9sdTRpoMNyW7MCLiN+OLxWnSQlzurMKnPk/B5jxunD03J1wtpR/yIBu7eUl30/GDhY
++LZYonIjAhsmyFcC3EWrKtyi4bA0E9FQNZSBhPAxd94Lpxm++25Lpszo0t+sbLg+tiQ3CIKJaeA
RhfvcQ3+XAo2ePtb6spMc7xh1R7Ia7rzbpgJ6XnkxOpRLv5cp8QH86EZXfMpsVqLIrCy+KIxemry
3kBbzCv5swfA9MgigKVw0c2hEYGMy1HMHXP6V69xevMB0ah5GGQU0Qw9OGAFYmilZxxAI6X5HhqB
i16iOKevVRzf+35MrHoc9DVuAn9hL9thu5zBKQ0XEwIHFWA0+H6ohHnRWh6hqi/uVFiuvdMWD4jZ
rsVMHPpENkn7cnx/3aNFWkQQIUvIqUnxYCgRzyxN9BhQSPLch+0rVH+nCGNjj/YP5qs/EKdVZuOh
zaIAULbAG+VRjELYz7go1TF5HuFpX/lUjstF6AXdPQvvdoSa6dnxvf6B67NJopteQuW1r3+ura+e
V7M9bpOa8ErgRwkSVgxYjGOf3GqaiTWIe+c6ZnZAtz/Rd7vrkdfL8sqpK8NNxvQ5uIbI+BmRU9Tj
tD1N6DMdxVuh+yKISk98spf7oGWL8Vk8nG16s16AJmrLeqL00pKOwSPcfz3ZWSsdtWzQHIWW74AX
YdHvVHuuljeA2DQl22ldLt5PJtgSisbgBkjIub9dfv7IPQU+Y+SQgU7ceBxN27yBbs3tt2S8vyGF
JVw9adS7Ghd1rkMD1AbMmx4Q12osNVqzzDANIGZ1ORMKy7GQga0oMnmWyP1T+bJm+HaNCaeMnhN2
lEmetnM7eZDsc1/S+Kn0Wh+PlJTLhVjt8BI0LpkQdLAhD6RvYqdOJa3fIVu7bgcnbOCTfELLZTIH
nYK0Ixo/OLFo5k4zia0vtFJQM9cX2A4AMpe3c6JnOHhawaPKyqXE6u30wTTeSLdOUp8D1PIV8Cf8
r53dNTTi8N+e/NMTzqeFHO8/Ythth8hGFd3v6+SbMzcmtUscslOw+DvY7Sjmde0lliqF3tDUPaQo
TuZtIEWppeSZwx/yLbu0hsUtZUhsFNr6ka2KwGZXI+M2SwGhNuIculAKGJGDmiPhpsryGNfKe0Sk
jNKi1pFDaF7vv62CGiOeJ62wDBtaslKAuVjdmvKPV+v1/hzk0+1mQTWzAqiqr8RmQ0qSDJLARfqC
uDeRF6w1IR2lShUNhPhT3bPBjdgXsL+OsQJE8Yh57k8oa5hFbvAjEv7XVhnCHON6OYhYM8NziyFi
I4zmE/mRrtC0pqrviIWCv7jhoUvO5qElY64BV7EdVNNOt1BNgi2O3+OPE4ZtKv/YSNn/fO33zC6e
fsaXy1SfuaIqP5DN8aDvfsDEFWA7o7KYCB1ZtNFyjp2gp4DC9BgdSHx6SahlfB08tro5Zp9ZvdFX
h+Vu9LCsHpmYZCL0x5YzLX1JrBrJPIWgQ6kLsItlgqC2Hln0l5dq8cPbaGzZ8vmI3CehkBzVpRvC
4YlcUA+Z19hPm/hdX9VdC6v3Fg6QRYwAMc/yRzFd1kwwZ6Ul1ERSTAYlYeL8D0RY7fiveOafpxqW
NzNEeqcaaqlC672kkxaS1gPFGYblrzuCymqA5VEFnInsrNRIxYAt7FjfkfhTW1NkoZuve8n2H3WR
J8MeqOKzXD6/bzXmnXvrZRVNBmeuIzc9p/cKzrWZ2HIuZsSghWT0V+IdiaQAMFFqo0G5cORdYcmu
CwDzBm5/5ES3ILKL4T6EA1ZHV8qrXcySTzsgIZ5axnmBKQ5MGaQT0T4QqhSyZJP0aPULRMG+HHoM
ETp+hPGH/yiOfuZK7+X8AIdJPm82FFSyAjUcr4HgLJ7iK0X8vqcAPloHr2yhUAjvXR1nw3frUepa
S0TFKUCSDThn2aqEiQdmpEb76aGBs0DZSTatPzZH5fKqj2C72QjRl2ZiNwAdHWYirLbLeEXjxATK
55EYcixpyz7rAYZEw1O/b2DLArNDMJMErZfY2ZxSGXRntrb4Sz1oM/uytSOOZn2HquUhSmdHSgOw
r49Ed6DhONPIVo/cuG7B1zKWrc27lInYyskR3QqYG+IvQSgEeXsnc+086B0DpFXwxxmJK4Bu1zLR
JmXNGp9hLARYRMr6j3LZtptLWqY1N0VgEE+Br+B4LfrFbMx82s/4+5xpcDc6ERDBg7HZOREv0Ste
diqrhbP59gpQ8vOlP8mvCJma+2JYVQ71THfmccw8UnFbZ5c1hei8rlFIlV+rEf086dw9VIiwMadi
LevWGWqMdbJTDGFsp47AeW3GHU19k5THPsvMjZZYauHxmvw8Jw06BNjjwHFCr1CpYmYE3Yrb7Fzz
aR4kl2dXJUTfdM5E1qWvx9PegktmYShj8c4Dm2NR+ivVFvTHhstqxfoPGhj2MraLFOXIpqR9CCmk
4+iqLBFehSqqvtLI8xvz3MHkaELEN0L1BDxrM4ySElVZfV/3cRhuwaOVNRdaJY6OqUlTnFGjFf75
JZKuTyx5OjDK7/yQkecTvlKk9JnPximIL1JCjCzT5S1C6HP3J/p/4I7gYY4h2i4ITkxio9K997Xm
Rk5S3tT0ksA5/7w0gbyQXV4Vnxn+rDPmLqlFtVuDUMuCYRCV6TO8tNK1pfBA+MH9EXcvFSXGvVVM
nepbbDeyNzlxJYwJsm8b3O73JUDqfOK1pl3UqVNKHbnFrBeVCjw3/9L+NqxutxTEZEzuA9akSMej
uRm+Hnq/oJ0tMOgeSgtUJsqglYBPkuavXRd4/Rm70QmNo4ubiTe2EUcwvTfe38LVMEQwfTdPmix9
lyHScbDaOU7uhBdiQfW5RmNfq/xxt0jDfDcZGY9ZkOQ0DoW+2jlDTps2EhXl8lSjaIdm2AuOZurq
rLhxZSmtZPg3pL7OUpod9tohuQgF+K9WgJg2L8cIHn73EH4BEVVCbfbhl7VkH5oyfIk8StIx8i9N
OlUA8zTqz8WGHaaAnIMkdVI7GIprGiNIhSgeQNuvWyzMXZC9r9245o+QXyDXRGsq8qJTzGQJlawD
gvaabDRsTpISoE6oh/C/UsnSmDbo0aUenqkOI+Y/ahA7w8U+/CXstSN0LqdE2D++mRzOzcwJmBPr
hI/nK+BBPClNn1sHjp/2HBn+DrkWBxVXYj4qlVSXxqpHc+0yKoAiymHPQRzuSoMLy4XeL5XRaHtg
FLnzt6MMnbuwVb1HIDBs36NNCSliaEyTg0646gL9mJoG5HkYX8MJtqkWOZWZoHr+NFpABPKiWlBc
hhUN6Vt9FE3xDoJuhmEN73/qyOkaxSjYW/i3GXCLlDcIgpzrfy6g1wX198d8cpXkBD6xBT9uRBF7
y/D0L+JsSJYv6DOFS8+SZ5ROeu8NJJl+15lNTSoLTpKf5k/WcNDSbYTaUm7cZO2l1+RHDgqwJQTb
B0ojYvlH+hktALc/5I15xLsb3blDWghMFXQCJGpQfDrp//QoBgnW0m8JoOak1hOwXCe1DWNE+bN9
eSY72MgvsWUe/06c/s6GklC6xlyhTVpv9Oy6vUMbrg/7hfl4DsWJYWoei7r64sNOPi2y5E85DJq/
2W3HSQTq3xLQT1KNaeMNBps8DUYRQ3M5kfkejuDxj8bXtiPtA69Nsgi2ySKSpXaYZ2goDn79dGTf
JNqXC8KKKduWmCDqRPvcRAz9XGF1wF7fOYfAr8M9HDLFy2VJZNQVaF+7mxHQFprqAUCKOiW2pYwd
YzplCptWoVkN+x95bavICrLaUoVfo1bzV9hCubrcNRGrYAt2k2XJcDaJVaCKHcPh4cD9YzlpaLof
eQGs0QVRw+6zI4BOkmkvLxVcN62wuJtSt5m2oVLIm3mudAG0vCYUbMz7rgZ/aAX0uMqKFqTgLnig
JlI9zWleE+GQiD7M20cdtFrG/EK0UwjnwNo/9R1tPU8L1K33pHckEiJmIxORkKpy2/YnpHefYMjl
TeFm0eJMNc+NGkNGK3I2beHcuEoubDa07RQR4xi6qp9DtQhL+uK19Y2UHcIBgKhaYNv2qk/fYSlB
1OnouFHCdVLKIfAWMti/jeTGhZ/rncdDJpC+S7naBvxIIjMCv93AogodMnsqp6/ZH/Y19xbZTcwK
s3C6Zbr1enItb8RHFo1aoH7jnlsWmQRm2NlpU7LRSZedeUuPJ1Wko4GhxgJwhrzcpS82VVm9IMVM
2xHlpEVDqunrxbOJX6WrmZO6K87OrOwZpRhiTzl5JWAlB13SqY3tA9aEJJoJAFt7DQNPgrWy6vEY
TdM+a7JO8vir/0mpbLixItzHyyuE2pu6/jVWf3JQNS7rVcnDclCH7BlipULLe9f826iILf8rTwi5
5kaNvtmXDjJgsntCuVADceY2EkiI8nT7ozAAalgKlA8aNDkvqPN+xCmMRhtlrVR41DvoLKc2+79Y
cZ0sWkatTSEZ0reDv5uQmAmSDHWYeeQorLd2wH2gsUPV4gMrMzMOaEvFo1EX2pdmQHPT6GNbQBZ7
20UkFIlDNZ1wFCfRPjp8+nnAe5SokbqEyrC68olvU8VlJFd1IzbJ/dfbngDO+Tp98ZElBDZ8ZzLE
O4Lkh+IqVDY2+Ta4dhJpdeGdkBtFm+/tzekNsTAtBXzdFnRSfslXnavRpc6Q9y/NZUd9q63ZNDXU
Zz+NrTtF1ZqR5HERUYksG1vzFrwb2zit+/+OaMr+CKhZFUdXrVJZPm7bwxzbofDj1Vt5o1WVKm7o
55Mi5/h/tgZfcae7cIygGPqXOsbUUIVBJJitC3iQFuzHfCu+axr89z3OwlqzPVTBkEpuE9PQMtPg
dM/q7qcS3JTiSk+lHxHh1GhsBojwDljWoHx9uM6S8QYn4xCjOQBnu0d2wbkiR0Gi5Z5sZwvv0w4c
Y/O+ImNiaeVXRhFUaQqvtaogX3w2j1iCDFXYgfwbTkRowmIte0DLGNekb4qC/55ObIaCVw4VoH0W
ZCf3ZJ+frBr7gqdcHfIQp4kq7RpiIo9t5L+CebYb2498dg7KHBP+aDd7lgfV/JvuT6BhaGbPpu2C
nQhtwbsm4amumOiLz4wTVmgDZjbFakA8v+qLOL2peyX2ZkPDlqzwKrGO2J3x7mEB9j+0vnwzn60N
1zfVz5s7iOLnfkwfFGi5PXMnU+tYegU5IbMob7eeJSVhZjV7bFLyr8PJFXRikhka79JK0l7oTAXM
6eCVTi/7X+p2AXKSlL7I7Yl5O7Wav/USA2eczWh19iipLxgzPKlBck1hqzgTD+1SLA6hBF51QXtd
KeUEfFbQ7uwPImZdkwDO6ueyRY9E4EFrY3Iz1KOyloQ8v0Biw+05MByt3KeEzWJNkH+DZ3/77Whx
z07mKZeWHQwYg82isR2DhwyQ1BNNOF334uSvmTTvfXjs5bezIekRIdlyZdqJNO2v2Olc6Crq3Pyk
txSkBUwT7k3BUNByxidTJ1VR0Qn9bneQeJJEzo9jPfashA5UIr8AdS/DeIa2nfasjbhqgFcpbtkg
w4w7dE9sP2xcqxUJ1OkQvKg9ixChXTmLTMFK9e6LWD8KtnoRu5fCQgTlktl8B5OACOBAGm6MBJ5E
6WGgR40KoVJDOGFtKBrsOaiP9rVRvmntxIg/Xpemks1n9lWIWo2dy70OHjRz/vMrv03jlcMGwgkm
5haCzF79Qo+PF7S/QNzYjbk6XbqE+jkvZlMLobKIph/ge4UJYapG7TSozu75+69evtB2FLl0Hc7K
73+x9D0ZYlTgsnKZx0YDQiJW5pMBybyayABrT52RYWkRAv7bmtpx6jjSdJKy0ohPSmVMrK9OrftQ
19ywqMKUdkouhDsTQFYQB4XL14zUYqLIdjwmGIQ9ZL6+sya/MgfjWurKIu/5mLP5wps3CfAiOFXB
dSh0v0VO40mvnC5/N0OK7FnRBfXUv/hAt5M9o/camuaTMCXkxPkw9kt9wT07fsSRqacpWh6IDQ4W
ymNcjzq0jTtNTtXVaLWh/PQJzxxFNp9sGNR9eWyjmBP6+UYUmE6/VJ1hF+2G1VMSU8t8Oh3skq+2
0zmpgpIiwqlDCA7PHDjbI5HDl0XmhWP6PB6mVB37TE+UmBSYPmXDUjknImT9ciRb+JQPGA9nY2mE
ATRnqNK1OVpzNTd2GqaALiX0STUUNKJxp4TVkXgHwww5mwiQdQQK3yDSm4DL7osNFdn35EApCH/w
ffhYCgHFCrWrI+Sk3/Po2IoGcSKGolce91rWMZ4uynmlU2OMG7Wv82UqghzHzV7pluSwoj3wkv2z
hDt48VhrmxmAkp4wdOu2BHMfIgVykZvH++L/mXdGCqZSUmnu3KwF0gNAer0H0AOpV6gjoQWcME1f
6rZm0sW/JpkdaA2BmPlQvP1wb251KvNFbDF84LD88zchgtFzSivBOIg/vm1dLpvgGR2L2xZnz2qE
7JlGZCYLhlWm8b5N48mdpLM8ZYgVbn9PwxkSwiYUacpulO1V0EHHM7E8Nhfd2ijo8v0O1+gCf1FH
fKzVA7EYr1DanTmd7sqyYcPD0d4qYzz4MFNbobDyfct9bJmT27DVnEILoxxRUh2oxQmrgNLbR7P3
qLTuwrJIAQ6BMSTMNP+/vRtAGXMOyQjKPJB6NJcR4X6jKwqfzEg0YZ7eyEor4TMIfiiJFnftg2Ga
k+7KKwRfrQpboPItAsm7OgaBdBpnNS9ntO/M2AVZlkdQt6HKfaBwlBzsKaY5wFXMNf8Dgov/GITW
d3HX1wZ+2XEV5ve0Jo+1ZnjbbS49VLkQY3/KaMhDf0YkiTv5ixnBAKujRwb3x8e/woIQSz32r19m
4VvZJJcLpuAHcti+m6X6Gg5bJSEeVQbvU0HzelbiQNTMFp4mr9Pq5PkyLX4x9UUkMDKLQ5xNJRVq
aK0PT0bBnpBc+z18q/B+OCU24bTVoLx4je5NsVntnFI4prO8TjulVEg5cJMEcMYColKYM3A8K/gX
q9bzogHlqx9lfR5HtlXNYktXwQlwIvXHwzVU9M2NLYycaRpPhxw8Jfx3b3oPrivvipPTjeqY8jd5
s3vVTleiv1z9JqbAGZvUYRYeBbxSgYRKvQV9xvbWKP/7T1jGdp44Dy06sDS+1DlZerZM+bdfuokB
sW7/5v0iiYb9x++4M8xgUyelBEdkYlibWI9q70NBzFaOgjbI57c/dIPUGDBATzb2GLifUSzSujw0
O6BoK4ghOF5t1hdrbYvSf6bMsbPhsd9QwdpXEI8Mo2tzLl4lzSpxxT7ItwlqKCuYZ+9xs6Fwvdrz
qvWoIXPQiz2nz4q+tau9BBhrl8oaLqkzglf9zpXc2BB1AH0NsRQPeMG3cU3BFklRNORGvMBhBHd3
0RqM9HIycUTMuVzBCXsQj6GQzPA0i43oRPnwkCHFaHGTjI5QOtZ3PWIJLOo+a6nKUJJ3xsSqU2bU
Pculb7KIDyPv35276mkZBzbEWZI+yBckFfiGlmvJIPDAcI5t0PctP2Xiew3L9IYYTCprQlA2y+Wy
eMDJ7FvsKZ3Qs/DIkwMx8KXZUeWXPdOzYW7Ek9K7XXbOfrpzAZ+W7DvZ+xPWxANYnOM+Oy+liyci
4KIpLIzwQqPBBS85UUZyKXewG1LrR8H6B2dU5v33OpdOP36avIp/KX/IIDNW69109FGpEL1IXEBz
hnhApXQ+qtlQ47ZBdiczbCV7wTWXerCDJW27BAu87mPIPfZvb264RtzRVBPxBnh5TsFGu4L1wcNM
uGxRb2nV1400T/DcuUYKpJ0ryZgdMXc4AEPsa8NN4o4DSrvAiEIMxzF216VwApVh8TU7QG0Fmiuf
5e3TVKW5cBHCEZt1MjuXkMYX03WiyilQ1g58Ak9fvJtTNyyoLX92UPiwCJgky48gtgTjMaRmb9VO
ufpnSRMrKAntS0lM7S+xNGVVGTMP+Ghk6mYMBYEtPYoElsXQk8r88FxbuRx8LZK8VCArKhkM9uwI
QLAHEPVgaOihk7x+VOIvLPLEcXiyXFUBQGvgYC0zNyH0mrYJi5XQBLMgVjTr5Od2rGgnCp6QGUCz
eoXJWm3gyjk7ZWK9QH0DpUkQg65h7ME2YKSFMFUJEtoNQpOv0t/lHofgq647xf0Eaeixjdr6k5p7
PkqFYnDwE1bCLQH+Mq4BbSNelpdX1XEoVPlU8CPy0akWU7ATXjq9GQ6y9GcdGW46vgiLmi2isWpR
67x/m4KhRxs/zWcEK7PwGjMI1zuZ+i7uIp8Q7dNHL6XwXruYCzTwQxHoOuLdHNE9mYAtMEvrS9gh
NSUI33SNG1XvukGc3P4zcY84O5U2op8fbjnsLZmdpgg5ghQmOms/VTwnTGWdrpNH0PnkZVynCPLp
wZ7/lN0jMsfn0LJo1gU7kiVuHjO7lJnDlCr8vggFcnGd363H152W2QkkmNfTLzc1bDQa3RXjcgAA
ka2VOxxpKzsoLmY8g4id7yiB5UqpZIM8Cxyazk9mUyh3ciL25sRk9pRJzszdTIVYssyBPLPJejhI
6dP6lpV1m45j97liZi1+zJWA3QAfMAK0W57fQlLxgmXw2jh02P9wjDgPjSetCVAIzGhnsWcKPqeH
LapppoYLeiU2nTxEFquzuYlzxYaGNo41scaOi2aCrN6fp0vLxUTjDtC2joreZJYbVFfNq9gemGHU
4r7BoVudpTeOTp+d/T/C58Fx9d/vx9NdMvFRel/mbYkMNlyrg00b/gSFSnFzpOuNMr47Bz+WwKHE
uceixqGWz2qf0E99xr11jUmvLObuFd9h8+zVQiGVrnvA9wa/6irst2GXYeVzXtIU5RSwMvwtPE3a
GDIUF4zAcxJxlLPjczXxpa5/GhEfCICYssxHXkx8+uhYWSk3anJI9afLSBqjupUSRW252hIQpjaz
4Pglk02dvQ1nve1iQbPh6BYAtMtzeoATGmG6fmlJzTvXjHHPelD61OmUTqW+k7Us3txZ8rCSw00n
NXelzg2TXzb76lPPDJM63KcHP+NU2ugoLPlKWUTfIYoTirYDJPg6vVPwlOGh1Jes8TR2OxNRzqgI
VJF7zSnXxtZvuFxY8f8e55xB0KxfWecYENTsqMbD9Zv/REn4EyxzVOWBI4MhsCgDo/4hWyUQC5WR
W7R8vJAvl8kuKUTeLQNOIU6La13FaTch8Abu4wLaDxbvY/NFTuQIAS2YUv3xVltuFheNg7/JJ0ZF
OWZ7xD9KhHcCgiKFXhe9TNaMd2DluLEYt2XWX1kfomzDzoLL1nHCJVKzsfSkcq2r0iRw4AuLJfDj
vhaQma1YY5Hkb1SSdJ33MS+qqqS4XYSQuyYaoD0hJtsROkvDwtnt6dtZm4Z0v3GDqjB49Bkl+dWI
kZu9dPTstcKG8shNcuPfhWMmZu4jjF2MLY8plO4U3V+XMtMEONhM799h4mVSU0zY/jO8lUbLAa4r
jX1/bgwELvPQhoLO78mj58r8KBP6QBXC44Ko2mSI8PXnKBlDD/DYtiYlp4CoJ9tJiHz6HxTM6pVX
EhRA1MTam8z7gcpdb/7HR5QjFUNOd3qAkpoUPEF8D2OEAnIQjLZ1CzyXGryENS9kevZz+vJtrTU5
Du2xuJJxPaYbYhXFs+39x9pZ0N1tit/kqEHgryq4f4R8j1fR/qg7qmQYaQvCbzB82QNGiHbdTnj2
F315/mue/EwlecNQ7HJ+gchnfyW3m/MliEHpZImzhs+K9N0JFMbI6/1e5ZBUCRzf6/5qtwubpduQ
QhxGWWwTfQ48Uo7oC3c00pToWjFBB4GnnLSZ9yvgT1o9zwYjiKMWygTYt6LSJu2Nu/4/EFgqOEPI
ujxdhs06MnX8d6WGln9//fdP05gzGmnq8jmgJTEEPG0UYqvxl/irMh8PxkepHVjAtSQGk/4fJq1z
aim0fnJQvLesx0Br5/GXeTRXVaAgQoeG+9LLzyZFC2d2N+vdQ10LjHhaBU0srU7Q8ZSwzOi5rRam
XeBqZ38ChhGFB/Z5CP2T+p+sZuGUJwNCX1MT20rQDx1EkLN8SbhFfKl/dXtuSEaukl4A62U/2jFq
XBQd+qBnyP8r8jhg4G66TLQ6Ms+/MxUrDCe7GJwQBStn+3kj4FZgkvzeCxWGg/J3ntY6cSNvXz4b
jbYN04YELaqZCXuCm/AT42qCkiv4bB/pV6OigZAgIo310EvguBw9k30Zp2oCsWjkk0bAQweFIVTU
HmfNqEwK+x+inW9a6tadBJ7BCAq5/jZlKqgC0GEGcMPXB2yHOL/Lphb8xVojA4k7n0QGL0PGE4pK
4JdruKh493Z24fEWtH/6bcquDIx1BhA9GdvmfGJbtiwv5fUOYcn3VAIrcv2+FGejlmL8taVxi62p
stDKr5PxLD5RBvw+iZivTHKy/1NB5kko+9G9IA1QUxUrlmLHVHO6f8h5m2PQqEbZCkMXiI8dSSD9
XsycQYzF4nFuS+zyNdqn0bOGe6Xif1x7X0AWgO2Pttx+xyC8tpSO6ps0JQySkSAdKAjVS9iMI2Po
zkZbfxfH8npnFZ/o6ngYcPR/M15GWjKtVVCMWZo/pLWeoZGEIE9kTfnwGPA8rxco+GiMg+EWKolQ
TaMrRlBREpMPDD0y61s/QzAx4oTUDLus2CPhkmAI4y5YX/zFsYEt8/IqtlodlCsFSayZzg3WMkgh
NL/aSzOcrE2R7BwtyOEGhM4zXgYVliqYiOLLhLxhBGqBc/s9+UGatJ3CrXC/W9BOS84mmTSeJJZ9
jWdwGnmNzPamRr5llKzYCfDpQgk40t9orfXmhUpuUI3vxHFzjp9CSZjzU2YjLjiD41+zFHOYIOz0
IXGAfZFt58joFMbJfItVylSzl7R5HwEIphW8LMADqRnXAef1yokGhtpEHmjp/4HQeOmtZJWzyOXs
ALA9LdCfqRKPJeWU1gkpP4i1vAK4Nep3gKdtJ2E3igu8uYB9Rh12UOqo+l3jmtIo45SAsX9bsg3w
xwQ1zwnyffpYZARvdYWAN2jcaXzVyIybRnlvpSiGquikcarsy6JJUEPIO7gdLthfVRyLjC6YrRae
8VUW1nBiDDDpt5B1PIiIHVa8MwKUStqt9oEmbYvTWUyTh8UZ0D7vXwIbdL172n/zxPnJQMDDXhNv
nq2h2/IkKOx5f2TswNAQv6TT3NBzq1xlDSdSh/+p2jcAIFaMDAHngjWbU1DLvFV3oCiLetvdJ2GR
r8TEramEFdx5qbRQWVCQkD/uZAYyA14cj2v15RLm16vhFR6ziCg/7RQPiL9bnGPOC7YvvozVA6Il
TSfcfFBSW5hjmwtHggUPoLssygPncUrIxd/yRIcnCnBlb1M6bpgyZEFuyJg4aV9nhX3RCxP2FVG8
Zn8BT2fBr9LhByqlF/IqgWXwA5fC5sd5QGc5vCmetnXttxJaQlInJzqXRFMGYF8jApfIwRrG3i92
22LuvAAzO9DAa53+O7KrfKiMfzeajkUud5O0X1sbU8VeFZ6/IVRPOSx8fzNKTEn34KlNyLhQR4Jn
skIwcYLTNvZEv+eAkd/pjD6L1xoGXFPg5KraKPj+GUAAnNAv51QVVsrPxHVoQW5fK+S+qk5/tNFz
FdM+Dx7pNwjFXl23lY1Wpg4ZaAGPzbTTOWOSJQAjttRqrqmQ4mO0KQAkc6GwPBm9Ek4H5AvZB9YN
yMubsmh0fY84vZ6Ysn1Unwey6GuMxVnFiUkhVnE0wvZMnTBY4BppP/5IKiNHDGGlj0ERx6NAZ8y3
E25TtNQfcl3QU4jVr10xpeshkfEapg8fPg8Lbbub3Q93/kRN2VyyQkOObE3DlQ3WTa+sSi+ip4EF
FnhOwN517iuadsnOQNB3mA3alTPe9a1BT10cg0lSfhaP0uEzVXACd7L5wTuQe2rpNy6jCA1IYGNW
D8FN1qUyVZ9VLeODSXKFoYFSbHB7akrnZvPQkePcAv+9PH6FgXS7mIBHgEKCIrSEFnnH0wERMa9n
li+s3+IKcX1WMvkz0+I493n6hviF+M8GFeDsousd13IkzqFyNCaTk7CFLAcmeeX05UHRiPmV5two
QHjcybISeS9nzwFRwD/QOrvwKgxaFL3qEJZKukMf5kau1yYeDGDSLYsLEMhq+HRx6LSlBEo3RpNE
rTaQuRW4Kg7f+Skt0WK4M3hTociwCxjmTngMrNfpL32ypdq4lKYx9diCBHfbl7w9S+fYOXH1m40g
iaJd0tG2motv/jXVryhQjh9M/wYc/81M0YR5NvNsybUhw+99XH6T8u+8cG2srVfAxjwdatmxN2iL
Lg9ESqY+P8yVEBXcMU4j5bJVP/tMEEIuNWFPeAzYVlmm3ycOPcPqbq9bSpWC7chcKaeqmCoXPCvC
Th4aqi5HUF08WPNXovRfm2lvd9MoC2ciclr8rHbn04Q8F1BZxK2CaaOBwnqGvy0wNKC3wRLI+Txv
SIqdc3XOfU4GkDLTg7hUA8AXgpwkNTwOVciu1o7IFZ81d6QiwSeSsdIiWIw7/i+tEgE7qXL8J94p
oNg5OhUwT59adXfWmVjTY2uKUPmJya/QQQC1Xz7ebYicPlwo3xyxqwoAvveVreXmzxkU+/b9GXuZ
85fgXDGZs73fYGU8J5olyAmlUGNJX1qE13tmHInX8+MxRdUCTrUkM4qRZpcF014QpeykIeIWnvzl
G8uul+/Rm13+WBBDEBjHs9mVpJVyH2WGxXe7Fkl4eHYTP49gzs1yeHyuoz0Ql0VK54pkaSuAKiih
XXVX2N91y3zgWYSYgo1Y0ghDphC/OA4hca8S8kyS61XMD+mmWgsnMaDUfEqS03GxhmrnpAvCnoj4
hHBMsBowWQt17eLTPOwWXNQ8ZAYCS4dUY5ZDFwDW6yyUxxjj0x2est2rGwxtbWd6iFrJER9RRfI9
cLZsKI9ME3jhyEZHIzLs0/eXNma+U/6mhyS/7Hyw3gv7DZMgQrC4tSI0y2GtX9JLE6ljjLGb8EDh
ydg4fATUMkQpmzK8wPfPTPsWU42e8hI5vfKMZz3prBiVztu590DIkcuAntqJ4DakzBJSk/mp1wV5
vMxIErf14+4xFtYzh66IqTicpYBxjayRb5xLTi97kKNwG3p2kF9Ezmm5eB+sbLAjl2iJ5dFlemgQ
YysGUUrjTx8A0QR0zC2MoRcI3YnYbO9N2CWoHXLI4PJaQFZwFsSuRtQWYFRWPDllrH/YNi+lEPpK
++0NO1wufxNEtflVi5F9HTaM9jNzG3KyhxYTW4wvZXjVUL3wijCR51NUYxJfr3yNRuSypQnY0x7E
W8+7fsy1IytKepkjp4QMhsjvFaR51zBtJjMM6EVY2/IRyiRQ51IiOb09cbCheeAtD1bimXchDKSd
sFaGdIzs3qPlVxx9SA9HPAkXBnbK1BqwWfu9pZCSuaOta1GgosRtpFKD6Sx7LaOQAHBBie/tECR7
mw0neroFCfKoKfh8OBz9AP85KklKpIEVFnpMAJwqp4RNXVGvEr19yujpVgGXK0JTGuo3rEWfZnrd
2vr8fzYEU3aGrmH7qf9S3veUKSkXXEXKwmNCbSJwskkfhm2LJzv73HOS2eWPPNTubC13z0gyXR8z
WpI9BXSc16YkWuWKEmcJIhtygPqYKFQe0f6M59fgdpCI8j1AUgJopBVfwL197RxYY4OzUt6j4296
0cnZ0iGntHGS9+/i7OC7zx1aB3yrfL53OfeURuEoHp44v/wl1EMogk+yarU25+I/FWtYYyOvBbMn
SJl0s9l5q2dcApbcEpdSjvTbeavIDOCGb4b2twwxxegYbpV+42CxeyeIFvJBLoLx6kEn2cGIQjK/
Rjuxf3ddWURv9M+XR9taY0brVUgB8BzD/G16vL+GSQEZR+DXTLt01CGYhRCd5D6V7pLB638A1SkY
DXSkdWUD3n+w8ew+3yv9Xi0WIzqmHaW8HKeJDdj9nsjiil8S+YFyx54VjphIJJjIso20atWr4P9f
U01FK5vzPDBi6bM8+w9Cj6tR9aerACq7ksuHOmZSl0tlzI+vsq1+xeKFwG2ZEgNTP0g4CNAAY+zj
AWH/m6RpBhejFwyu1FadFIvSwHhU6GhYKbhcd/hbFjQHjHkd82gegClVW+ORXsx6aKM4eWq/Zh0y
nb+q42ttOlF9uN+nwbOVxijmuaG8z44rDDkbXgwo6lHMxg/adcgBhCVsrORXA9SUUnOvaVR+HFEE
ExVsP5eJN30uIDqmxlOVxSpY55e6NmnStpU6M6DwXK0yXze1DApSqNJeVuO5HUT4b3X/yd2inZaK
01Mo3EVeFAWLOb1D+MIMdU5HdFDK6V2Dg/gDI94//h5LlyDc5sZOefs2EcfVpBQVddBgXlW+0QET
FHpv424dw9Z22zEs68VQxoz+lJWYvGouqqm0PtBoexPKAlqgVZiSWhKjaEI5Et02EsMdNry7dbZ6
iu4XTnl4zwFYtjMWxjkOo/fQ2hqjTcUlb/CLJPXuIN6LRXdy5PCyLRmSaKbhfBI7pfiyaEuq6qNM
pcOWWbEjhDoHZtjZE7nJ7OXp4z1B1BPh3cCpq+jdwXYH+9EiHO+liK8B3dX/i/4eC1Ggug+zEoHq
xBRCzpfmW+ubWMmRksOnEaLWmc42NDx+cV8FJs12BuKtxTwKO+2LVcSl/SPXh9dBwkNyaz4B3IZZ
t/z+AB4vyLG1bn1QGfvgHVydzVu6yckX0h+g79vHUSkY15Gtfr73YFV4TQ3X5KcUNhRySWj0Ao84
LnOQyw9klE4EXHaz7ak1r1cTyY1dPwdIL2YINvM8zdPypmSKtfc1IyGB0rqCMJCHS7ijmrynbwYk
IdNvhIszkRGr5CCp0u0ARpbFpWXU3nHEofDyJeI5lFOwljtZb5oUxLUwedD2VNUqA+OMOq5AK5nP
XEkOGYtnSEYdHOZZ6KlLRcta03MvTHRQDmTmDhTScv1mjK0B9wqZoK8P3atu6npA7iHw4l13wjQF
SS4V7QMUx8AzYXBNmxLhR0wlh1heXN3UANNi+H9X4Qy2gv8NxXYn4SeArMZMUDQonDb+OPhk3X7P
Etn6SC8LJfm9+QQDEZvOG5bv5Kga/6t4F6HvsJTKwQkOKnRxxcLxD9KIulfv3hGp8a7UrqtAKgoL
xuQC4NNObRU8EfUio0Qvhv5qlfcHLWSdBo3tSLea7+dPpnOUp55imuvImQazrKkz5R6ym/BPsK6a
lrPjtjoIWxYmjO+ktkkUprgO/djbMUJMk4jEeFoTetRJiwJvO25xhYCvayJSMFs17bNKVYYN0gF7
1yXYWJj2NkbEZ9tsls4LM3oaiamtMbzz6xODtKLDrxdthCDpixar09nxAqwhxtgsR4yiW4t3fUNG
yRp/mXcN8TrabUkRDFPrCdXguSmkjWFkDcMmADWC3snE213o+f44ylA0koa4kwCjun6b/Dyb17A1
5ytqTgJJHzoXqeHpZ9ouiQqBYrVZkESeWDD5WS/U+eRap4keBU+cPYFARRpUBjbl8LmrLBAQqA7x
LvSYMw/dOyS0jMN9XAFoOICnuXQQNCQ1JCiqHE9+rXvpMp7jPovTCNa6qLDU1wzf+QY2ijIbaV/f
L3rm5mFyiwHPOn9j+nyznHFgXmUSpW+ysLP0KgSLplovnIOcpEKPRAYnfa3Vk+t8LPi2UZQ9DB4v
94xOhvDkWLdkGqOU/ezrddjEjEzLVP26gQ2mXegSRLXXJE3VtQC+cKIrnOjk0CC6/A9rBBWoXkuX
G5Tt3lL6+gL2Id0gg5KprQJIdDPXymGYbe8WdPjCETAEv8DZX3HEGQI5r/to6AATdz+T9snrIGSO
Ht4ZO8RJuJAC4wcgrhicRpH0gmVWD+oXi7rh+e8llQQZ71XW0DS4aMR1TMsj5oXBLBcSA7k/v600
N6+FFtgI0o5pqltg4Z/Hy43IZqS8vDmAYWGiFfb+wHzuhBYavItumdqnhI5+chAK3MP1vONOCiey
Mk0DYyjpSA/OnOcmqCGbBcUqqfcK02WSzvV2ZcS/PhVqT+3B8xPqIkHJ0YNmD0dpr16rvvJ8sijE
iW+EjC+/gXTt/P96riTv1bstRh3FOyqEEFsc1sm8Gikw4BiNfFP0ZuWvaupQLBkbFMt7SCoevc4A
pbClTE1A3SnwYnIyUX5ZEjlNKjf2M935V1kKzV7w3i9IpPfNxtKrfN29zmrqx+OzTk4IISODwvkg
vds1cwlqNnZ1xs5yJGeco2P/AnSNtQvc6YvY3rR6lMmMEr9C1VT57U32JQtwRqLP44ZT3dBO6yQf
fEA6xfDmDIfgFGbZAZAJwu3TPbhQpsId/YLQn9j0hkbMaaD4ipJ0TVZcE+NJGzpg47fN+Ezfken+
NvupUQ/KAdD0oBZUDOsurkY2Btv2B+lG9isANTIWGOpjBo0+jNkE7keeuux7B6m5U8nxZP2azQrH
J6AMlEvrLGJ1LhhQnTko7NaoI+VzlOtNWWU4RVRy13y8B8UWrW2ZqsoxNBgQydGMc5o2iPEAiXkr
KnYRh9b9+Ue0+41jNDoAMm8hfgnd9KGk3kImd6EPmnnso4sPt3qBXWsC4PBgqJXp0AaTvh7vmbMH
LtffxYgvhif9pWXmJSbnvL7IkTDBQJrd0MzzmEzsc4rgiqbm96+y8Sm5GO61MSRuSoA+0Dg7i/Wd
2rafkqmG3geea+bBDRzaolVKlT9LgGDkWOP0J1DdbXvNV0okCPlmp1kGe6OZDPu79CzaDggAEav6
yXAcAQrIZNJH79dfZiJ+Tj0huFacvNDkjXemMSySD+q1uwlNcmYjSEtvGbq8hHF8Y8/xUiAaDE6f
GSltzyPbMhrs8dJCtpor0jn76HfA1OR0QW7/iX9Yqtgt17fIYBz689Jj0Yq0F3oQWEB5n7A1ddrz
VFMxcj0Q9GHsEPHTj0e/SEqeXAW7v6FjceajwfO8xe/PM3QMyakQhLrywgHvVaJpNjMoiXdCEtLq
2PGRuK2MUtGO2MMAQAq+mvKvDUcykusW+6hatfIPwCdQmwqIN3c2eydLvwQQou4ooet9da3vzf5k
gd+fwhB/r6xPA1M6qbMbmzm2aQVJ66gwthBqntOksnJWjff22FWtTv+u6mvFPigJB+XaWbEZji6F
VUwiBaVTGZ0hPSmf52so6d0a5WlTA+pkuk1eu8vdQMWWBOPVmlLQx0fPtALHXQ/1BHp8WvwUU9eH
POcUv0R/VK2OcAd5qIT480mKH3ZsJEgYXJE0LT2qXgHy66eqJdusrs3DGTxcRjTXUPw9iryIA1IM
ZQ1UTSQYel89voICZsDJhm8qvo/FuHJBoo5HnCkojwjkJxh3tv9NgW2MCCNoWlUoZc8mCs5UR9/o
w0inrCvhbrWA5hjjwtP2XOtRNPQ8uJk3YgofooZReqoYm4jwCDSdUbjhDq5VVCU/2Wla0tBP7Z3R
m5SBqmOYdvn7ChmXbkA+MDJMWYGK8iCocbnlHeabbrV1czh3TxL6tjsBKHnghce4xDsmv/ov3ly2
oyI9qKor9+aQ2rEfsqgkp/oYDdQukoaeaVBY1LNjTE7uxMesxHCqx5wXLjiW4NlleJVBZSn+rRFa
v0xuraM4KeSyUY1sWTCJjteekx0d2IT2b9iGUUhacQTQ9t/maGr7lkE8gdpQD4jhPsZVyW1kgzpz
iqTcfUQ2wdL4HP40zfWJux/CkO3zAyCx9m3l0Mf5q0oGWt5obdcuQj9/P1iHxKrl0bKybnyKpPjw
GgMNGTNUb92SfjgLhUgib4K39rBR1Qzj4Mno/dMJlii6qaRjqGOTIhFTVVVyEehl12V/L4dGb8cs
G1fgH6ifYuApILyZ7PdCCGsP+XtXmC1Vl0npUqcbmlOoCbQzD4aw/y3ikAJTIGGmFuXtHMRVkrIy
DW7W8jPbKwxY8i+BWBmXdUs0fm/ju3NkJHx/IVcxsp7fhpVsbPN+JNzAhJ69S2gPvDVOzZ9b02jj
F1x7kQ+hk/ynDRtp2LCGfUHvji0JD2Ja+E+H31Jcpg4dSc40dO0Z1mg3aNTsIk9VhWU6YT9a2V5n
yer0gJEcqQOGJikIDFcPIjDcH6/dQp9ywaNV1sR9cTpsMAFAHvN+4Cd7fW238E4bUbORkH5oA+W8
Gnq1H70AUVD9vVe8ntGjAnEfogB9aVSsI403mSX7OeBjCgq0HxwkG2KGkq2ogk1h4PCR4/srFTOR
HNVNa9pRfqVhGqQVkRVF/WLCgzKm1WRkarnoYrjA68ApJv3GYJ4ISFrXnj82KI65zyedYqwh3fdp
PnYp1opd3Bp57RyE0NgaOheY3AfBdyFgMdMOLWJcnuKVWI5ZjnJzx0u//GU9qFtUD6vlgT1vWDZB
skCkO7/T8xc/TZFB+lk6hDK8rKkjqEhDgOeSKg+vBGTbku25P1BwaRJGkuFhVv7hr/B992dSzRVR
ZP1KmqZX9lbyknu2vRwGBD5r6Fb9t3LpWJZtXdE9X/ezPnNVeramj57aonNWUQrgC6pLMe0sQHet
e7i2RMcwGy+4KjLJZAOyD1/FCattX+h9y+zmsjHEip2j1NHV0eJSTspeXK6K+QwWjplRolOoddwO
N1s+74e6zH5zMbN2iQOVmktAonqH8Xk5HcuFvUN4y8QOk8aoIPoqEzU359CV4tGtuBk0bvejP1N5
kk1wPnV1OjexWNUc+H69qI3mPcbnCFzZwEpAoY0IpeWvimc23AX+qtzv1BTxeBXUtciIdKNK5ZbO
6yZ1hQlhlLgZnJp3QolLEx2BxTO+t1EOb37bCI9rq8WvBt+DBxaswsbq+70ndAjRHy+2pacDnNMc
qDQJEha1abvzq9AAPVCNu5Pmj4iMhZyGwI9ugSyhcN1bM9/ZeMVFNfjYOKSQoYLXba45nW0KpGT8
FcsCwUOtGVTt/ajJ+tFJ4s46lgWjhAs3xJuV7Smb6WKVeeEEZEM/5mWofkd79UKfWmqN/dgf9O0/
EJYvCPq7m9gd0t/owAuuA7j8+PcsYaYfK5g2E6THk8Ohu6fIqNG01BRcmxG9kEIiXAVabN+Xo/lv
Yb9ty69gzAMy1QFmSd+TsBLcTIM5WDBlQf+iG2mzFS7xlsTcwY6rgWxnZs4nvEVaEZ1AqLCy56KU
qoy3B+JpEU1KX4abkzqiEa0yfnChOYTSoXBBnA/kIAj8BNWCmsEvzwhb2t2Kk+undUx40MKWM81s
kF2v1BGXDUP5mCUGTDHB+wRXhFEXXiPuDIDLUXSRJD8vLLQ0NNFvk7fBR00wEZ6EQXnfPzqvF8ai
S44/ctN4VEj17l9Hbhbg7sLlzCUr4EdcU8VXXgp/gocYpfXQKYqlnVTprKZTOAG2OCE3ptNLQa2w
aaySNsOlpRQIpP1h3C9u5HJomYHf855KlVHLwSLEnxK6oIBIZpHKsFXvA5peoTX1cwBfz5eC85S9
E6AG7KwqA2S/u+v910qzJt20PPZ9BHmK3egMnnZbR9Vtv/4KnwjKIFtouwwI77OlV3dTKCSSKH2s
xcCrNrT12lUOw3/7WMflydHY+7ua0uPZDQKGId3bLzJe/iP5FivVI6NNAmeP7qA2rmdzLY7XdqM7
/vL7hbSS0DX2HKpTF3kyThh+nSNodqMJ/EuY+//eLOaUDC6K/WIK17b2d+nr2NtACF96nfvfcDP1
eWdl7032tbjOnkVts/hsVilkIFoCtmdSX4lFG5qlhca/OM4k6H8BVsvmIUEjOzUKN54467SOdNxL
npci19raAHCb3Xt76zQ+N8gsizuQ3TR2676b2QqHlh5YI00ooWPrvH5ZZiDjBiLnSp7k1AGLw+bx
iGpYBh18+n6z8rvSc/SvSxIW6ARQoelUB4EQsazRfqnzqObuvDtUfABOWROTb1Y6BN5o9E+IW0PS
qmRxeaiJszybYmg8wxowmAaTpPixCIf/vU4STeC2xRvYvBLBFVva4X2sj8SmRaYpgHE0601V+jEC
KtfQE2Xrt8V8CbRmxWT4QooppqDZRxORhgPSMyTxsmZPDQYk0CnfOORX/I7OcSwlkyEpS4oFDYNp
epAADVPhTRl0wUXqlzcoM99orgvDxAyAFLsIjmq3iZJ13O16kENZokCuFl6zGzH1RMeXahxvU+qo
2AzLjnaq60CS2ieW5Of+Ge0GdVtjEAoTQ6AcHDMlkKJSmtBbWjx1rLGQZBRxsCRCZGI11g22KV1b
tqW7HRjKtYlSXoX57VcgaonQ4aNeNP9/EHQdQbz/vccKYZP5sTjmR3qENlXtLIl1zT/IVCeGXDOd
bZfBoB2MVGr4ykwazlgRL38RqKknCDx2vDohDimwCmFumpc37dkz9Akki4T7BCX58lavbpXjM1B6
HntftKzRRXx3CiUIAs56aJCy907+HfLqlTO+zwaE9OOwj5hIXZfRKYtD8iax57p4UD4TljmwX0Wj
k14Xk+vxG8A0DuszH3gFq5OL9xGm4nTJHifDbH3WmrFzzusGqQYqBzR3KWSU9B8tMQEKcOzU6lDC
I+JevFsObXZiWuEG5rCDww3XpasbXVN0Ie2YcwQxF+QN5AhkMdgN2BMr9ADex9tsftfAsTQM4SBp
Nc0LP/G3C4EOVVMvsvSX+czqFgB6JB8D0kJcVHcyr01BD3hu7OPHCUO9hZH4Bv2j5T+F+mmEkyCA
7T459Cl050QlzxZup4gEZUhVqoIteS+z+njBAECKGqev9o1kuVzn6QcN/YMSBdc7bfcplfTH53nC
zrnXuyf6mGdK0xNxBs7EUMmizYXurwWukr+WVaj+y0tXCZbWhiaDbNQz9PdY9wl7xAu9OjRcAhAw
vvyjP7MoEQPq6l1PjarvJ7dxYvJWQkawBIjXpLxzMuywpRoE3gwUVQBoue0OqaYePtz0wD4zRNbh
4AXrGtjjucJ7bq6Fg/BlN+8LJs2OWHKim6HEqIjSkZJC7J1miXAODENqDdKoEF0q+/X/eU+9OkMx
or/+9c8kCqVYLEK5XOWx4418/6yYymXfd7blrWre7/6k+s5NY/P4OKz9+ci3rOcUpu8fvMm5bpYz
PuwEbbLQEDDyy9bqf3m/4/FQzPUji1v7ph57SkwlhfPtc0db9CsdvndvgyfFEFIOUB9+Fy6+9A8L
CnI6uMi6aGOiV4TaxMcR5MiU8Lv6P/eekjbMEjF9XaL5Mk81DNFPOBBhbLfI2RBCYqSB2s7XkXU8
rk5VUTRbseun9Wa3P5yRRflV+Oqhg0cV6sLgNaZ2fhEIzujcmCfqMzw1hgL4Z8FDg2i1nW8qqJ4a
Q21/rSuiJf95+iPoekG12NAEH/dXzh+oIBI+8yiVLiVA2IQM8zIM/oSACs+9Sp7vnbr8cnVjEXen
PRE0BmWi+In9tLBdYPzRZGndiC5HtPEfTjbl8CyFJIUj8w6AFLlc6HIbmY0IzyntJiZjsgwcO0X0
WLUD5VvvNpiamSta3xer7QIaJQwNddMRqz37UTt/9Gb+/IhUPKRjYzyt08uddAbCJNiRWf+l9BEO
MtdW6jcG7xHRJhMxeD1e2PzRXcLK4tEpLoK5Z1QEyZaTiQjL36ZKVsv9YKzl0YjpGF+uZbjZXgOD
mRnFtiv5aZuQuhQ4DZ9PQdqPGOqCbOS4fmqt7VuL34vQtFBoaZR4dctzQ90SLYutrQ8wqht6m6jo
Pe9osyRshVE8b+pbmpFzeE9M95VwgAbwUL4Lh3DP092tdG8Yny+1zttIi+5toviuJVdE3ECAXqy0
JbwXYwLEWmqUB05gukxtd2obsdg2rw5uiZXVwhUPr7/GCeVGzoHfcJMAiexT7UlY+N/tuf+uv3qc
EYFsq8WKdFjkpDOG3IsYKXOwysrE04kRgtstflMRtcguEvONwhPAYJm/K/yM+KURBTEwiiaGvk8j
owKuJw+gKd5Pna2SwLT2JYZgXfEkvebo7GpgTuyV/y+Bxj8HYdBF6+MIwuCUwdeLAB/LZa/Gno7i
AW8Lo81AOU7qcTWn+hLomvyuWQaZ+0LCm1vSgqrI0AKdzt8MYLXLwAMQCTMKdeb4bIgVHbZF6eUh
D0sYZbMswXR6qK0ieZ36ZoKHHShqRlRWNG0IeIhhPxa0wB4IRd0Pyyfkn2iR22H3WnNT1/r2oMCr
MDKDLv7Wb81I1aAW2472lqxGJAYUAQd9Ib6Lk+tTeh1UJJ16ZgQxvk2GpKhL+MEnGmTFaFz9azOA
radK2K/ZMCLvKnZz7gLUTIt1ENSwHnaKpK47I7PoXz3OLgc2vbEh0+n8iCgCsfRCxW1Cadk4yL28
vmVUQPQUn1WIPs0gFogGYUcO669Jugrpa4aFAj5VF06z/x75nNYLHE9DgI1u7pP1fOtZjB3wV9yo
hosOfDrIqSyHDHXmuSnoGxFEKCXiEu4vhjVO8IWVsEza1zDBFDwIu7NazvKaiEbKixCLmM9359Ko
gbD1wO8VMszJatCcASIoTdxN+fv2UjBGcfDsy1RRMknkBNs+Yl2bTyw9Ppnou+pffbZz42i7on7z
kkgcilG9BOxxcEmVQlGc2UIwn6pEsR7nPhmPCR9mVEr0lSXm2k6mhVne8i0qc/TSzm75tyopJZ+a
0BuFvGlbSw1gHU1kNO/Pb+awSOaAzDWt5ir2KAHJV1ONCdJFnJWv44oZZOxRSzSxxObYWdhIs7ga
XpBctxYauCweuY0n8qwy1DXy4LwU4rIosuyPXjva7AoTPFI2l0KIhuXgQhHtkI6SNRPweAKo1m0h
4Bu/dSYVm+qbdDVqeIumDgNvHea1yyYmuU2kL1BPlg4uPVifA4/udZjE74+VQRa2dhZYKOf4i9S4
h92UG1K8el+fX2hWC9sYzVXgAmFnl3lv/ai+6gxoDVAebqzEnXRjH7hww+yVmsINgZfXxsCHbEGB
0Vh9obpoJ9GYNkaAOfJpBcjaueRAf7EzMFUeVFExjm4U8invB4n0vsINmoZhmOXJ5Nw+f4g6GP9q
EfUeB8lM3kC7X7EOzEjxeHzbfUKmhKipa4vejMeCLeRFP/uOlnSBivlrCLDnD0450M3yw6n9WTX1
nabeeWkpHtiXc7AhcLBuynGnuPhgv011EsiYrS6HugU2CdZ1fXWF4dosiQt1MZ7xzkZ+0M7Z6Lyk
xKmC0WxhBGr3u0IgRsu+e46Wu0BD4E7GcMQEn4YYxlydqXV+cEGv3RMCDKRZWAfiSHRm2BWgBsU9
PBOKdigruPa5as33Ge2UmpUlubB5khWTbgIEY+y9q7DZTlTFgKwBI7HczTwQXoF26a8zUCVz6SxS
Kaqo2+N9Tk7/ECEoy//eQLWo3mD+bPQzeBqEW4ESqg4ErH4uDZkV6fkYHkm1TFMUe6ZjKxqupQ+9
dq5xKUCFAwCGJozNNN7u2+OAwMYxwLfaWuYJzSL8wIWGWwSarsgSS/YsefKx2Bd0E5j5OXD5rEWr
R541diwrxhvF00rKvOAURdfxhpMyYz3yrInIO4OB12yStYiMelZGEWpk8KilbIZlpnrAOivKqzPU
EmJYSBmjDe8sfXkMObHcnT9eODN789ekltT7QQHaflsquFKG0spKZXAiZF1e+F4A9ir1/DHsMg1u
pJSPgH/cTRxYl1tDeSbWUjYG4oa0lMMjO0ntIkQOluTypIcLbCwtIbwoMDtPwb/mSAW7txxpxiKe
lMujz4OBWGbuoqSYcB6a5Hxm//1QNBR/x+kxYohL+defAoLY6w376d/gFuxt+7LI1ZFupjken9zU
LmD8rzxlnStDiXoT4I75JQzA47bRPGuHYtphjWNbWVdArSSfSltRcJE8aR+dbBk4VU5MtIQ+iGFH
3hRXEnrQwBc/ghTm4N7BGRRnCFtlnMcHiQ/IAuB7Xem85tOylhgSE3DkUdEqA5YD7twz3wQuNDsZ
S9N8edH3NvBx3PmOag1TnxG+hiN/Ooc/v+RfC227lKbe9MKaJ61ZxDieufo8S/CK4jyE+cCGQf4f
g5jxKugZrO2s3bkFEJ9wDOCZAjwFOBT21rviDVPz+i/2vM5p8TT/FklNd8uxmY/Tlr1V3eHLbADX
SI8bY2G4uLjXSu0Cb8ggtq24+B1ftHmdkEA1NoV/hhSprQSxMn506CoOune2iDRCi2fuVSJyOqQz
rWRCcW0C7ezvU9WCCKQM2rFM9R8jtJq9cJpIRh+Egbi426WUZg6GA8EJPZTZDh4t2/zLjS0K0fZw
fU8jBjiNw8ZsmGEmXwaQRw11+Oc7D3kXH3KjCfd7Vr/69HehAsqPp1uPQ1rMj38LdG5MS3cVMt3q
XfLLRWenXUBuneKCKAKxyUkuLX0kqtJ5ReARiwdAsqDwLxaJicNrDsZDCqFqtvd07HR3JOOCyE6u
+arp5wcq/GZrlQXXxp2LO8E7xjskN5S+a/SoF5VtH0/TLCQ96JtjEPWT7nIHyDO5+3z5CK7nEfzD
ACp2wVrJSCcnvDFIplxl9gmmRq9IKR8Y0K74zK+z9oLTiQ5NomnhbvvqNsvv5Yt/8FPMbV7DRnAf
Jx5oDqP5UydNeuOFP0UqzHIRiQ1ZI1puvDhFDAFquU1gjZ0x91vO4zEtr+7GsNDRURpkFA23UwoN
fGsXZwO/pgMHY5iUCr57FgFBuXBOv7GNTjcsdxH9hWHFKb4Q0jY2qJKrJcwOGx+uKFnc0YKahvSy
WRVXZwiForg/feABoX/tIktUrVuQPxooxyYJbwEMh3GLNLIBTK3DHhhSijJbz6EvXwX4FCuYd+hn
/+LR35Duy/RI9yXR/SVx+tH6alJA/weDn9XnvnDJAmih/OQAaS0ECNKdEYUbkGnmYIFdlTlX5Wgk
EmB7OKY8kn1MAvHhtB1HNC8T50wIcnA6BZW4rGd9UrIdbqyH2RYsIo9BlAIvguMoNrFJpr0RORrw
14RJ4wqd1EB9tQX4C34YIyHgwIu3CEiu/+rQn54lAxfosOrTDSxmAkkR3oi8hGjzMF8fEGjYWixS
YJlU7LkqiDu9RxN0QPB92fc5rkHRzMIszy3HEsliNrGGQzR0kJCSuvdIChyirtSFo+4fSBlk4GT3
4qG7rhLFwA1oNzpOKOP434XBPZXkQUiX1/srTAw4ii+FHQaycd3zmMEPNBxHbO+WPzDkWGoWnq1t
Ujx3CDZ+8sVITUu2whjga4hC6T7wF7SId/Vau4WV0jXFIiHpbsoFVBqv/MsNo4VB4nJQ1pVKq6l6
KvDf4QVUbNvZJHsdwv4bKMm5sXfwutiNIUlC12KjYZxRGgEHOt6lVbxEhRsb4QdEUIMwdu8llJOn
JM84jbDy/C2nenaL+2KSZMIz6w/o7YMkUdTsvg+aNofBVNiuviyOJHvaL44ee7VVzUDiuzLoyqif
WotepHMuqOteSOldizWZd2834XVIhykFRpY00Ko8lORrcyGqeYyr93s0g9FxW+ac9/h4DJxfeiY2
Ym5Y7V2YttWQFzXta6FyYmzl1WJPicsnKOoD0HvZqkHhkT72EzUDdJ/a3ZIMd4AMiwJPnVbhs+Nk
R2PUEaPGea57y2IBzny/tcnrrYsFYRQaj73T8CoPU0BQWhK/ZdrBt3Fg0x/38eCLSREs7G3HPdf4
s6VGqkS75G1Q8+8morGIUj/tMzGHAPxlNT6Tr6UiqjbsF4e18eqJ5O1O+gshBZSBPRE0k0diRbXR
3XYT6/b3HeXtYc7WTJK2UtIA/yAcM2551bHnmC1llDHSrLthzoIFQse7U5fSCBofWOF4szm99iK2
DRg+J/P6348Jti4GqTroMxNpIbubFr/i3x8slK/bA358D7cgaIR3Tr8vp/ZqEoiLWh02Y7V0jV7M
5aLhcs2S2rj08cThSIHapGBQZh5QAMiXmddaX0KCQi6pJZ+4KYPOe47gJzSJUvCVCEjoq8gGT28h
9JJ6IRywIJi+WvtQ0nriORzk3y3fXlZxflThglJYi02yNMxWngyFnK4EPu+n7sbi/DCY7170ZovP
E7abAEbRMZGVz0Gg9/RWvDPmTdwXWdNZnDRVNvmY3ge9aZ6O/TCkrTjgicAFnbgJxG4mxsnfoYiM
vFyhMDxKZiKbv78Z1exjdyoftDiulhqlRp1awXZtHQR9HD1axZeWJ7+mUGFX5Q745f3CEUWa0bEn
2kyFXYXncCvanJNBUzL3UuOTzALKfog1HVlLXcVGhNmzkUP2dsc9yKFvyUmYo8o9RFopfRWDNyVl
qjkLSkvgbnp8xSVXYuu3YEKu3D3LUprC1jTMVoigSKqJ57B8I2f9Zv+ks0Q5SIajAtJffdkVINbj
yan2/PfAUT+0NOgyRLu9275q/phCNCXeh+vb/jl2kuA68uBgICfBisdYRrzd6KFsEO7frrDOtiMT
ZXH/1TPoipqaaQ71J6XKBCmVykBMokxf7eHzTNGdwfvAdpjWqMEr3Nl3pudt5lkUu4u7kcnqpbjt
oXxk3uSmm1YDc6H4ihgC7fYskgjiv9uLa//wa91CcjjYGhxcFZQ1fmEoaui/hUh8HO/sjRXNdsCF
WSbBf1c2sy1EHVo+huBunTqpX1TeIGycvAPbCTM9L+2Xy0S7JTNgKBXxXgzX2QgVbJsw95CymvKD
qzCxA8MzF26cUzV+1Q/MoGL7sgAqPhwWk1YMdZcsus8aCdjnNLiQez4rkdb6KDaBDOitASvo+HRP
o424VdgbARc+S5vBbQc/sdHlo2/+7rDMzYJmHAZC4HcOsGC+22E+UT0ZgreCBoNyVX1E77xmYF+r
rdNkN3sp2tGPp3mlDRLRCZQoRmM4wj9u2lk4AHk6qlivOm2eZ79aADrDvSou0Y4DhCVV9/yOtJPQ
2rXoSjuB3oRqsZBzQEniNfoVGvR93OoJVEVp2+91r6rLD400x14fZ90buXWy7RLJ/Bw+72whHm0x
LQjKYX5RLBQtspplAPjAdDnJvY4qjNBJlnU3Ez3oYXaAknjx43PnVTMtB+wwVVrnfS2gwf53htOS
meC/RpFY2hRs3V3Ip7zgJhse1z0cNPT8oGYcziK95ZJwVmNwIsnIZWh+5qBqLgkA0e81jzl67dlu
yXBcpzmLszFqYiir01iZWn8QcV3F5XdEcwFiAKwEEorVMXKZnhQyHyqHLavC2ceFtdmYGKACdwQy
EV+rySaWfKB5LXQgVleebL+CzUoZoOZhQh2ewNJ4fQTAiRSwpf4ISfcElK/6PClMmc3rD/ict55Y
a95xrEuybJwY+wChaOmmSIdNLePh23NNxb8LsCL68i8vLZhrnFq1ihaUts4qnUqwSEmz+8IZe/8Q
JEu07uOKDBB0oMjerOvKmaAhbLwNutDgIZ0lVkgiBlELdm5Fzc30wSeOvV3GV9uJvjXlYNa20EvH
6djVKV7TjZsyL6P/PEDS07usRiKM0t6vewmrQ9X291hZ5+kU/rWYnSBmxZ/EXEl4uZUp/rByOqSA
szHLSN23e+JrUQV1UNBOdLFXmVtxyHhKQ1XySEQrHpL+ea6v/P4WoWBcsQObjr/ChciQAuZ16zkW
SbwAHo/Fm5vagXRB7wlUF3AEYCyhhw4A6AGB101PVUKDyLUIdHMlDiIU1ne5kpE+la60RjY9AUTp
vWczr12wDG4AZSvrjsskjcXKQAWmPw0xB+Nc0qqvwT8V1WqriIr3tVDDN5RzURfSuVmFzx32CtPY
a/BGNIy77kUn3SoNUOUVYPLCSt31Ofn4idBLK3EduntbhVD0T6rck1UsRX/qSeBOEzHde3WRQM7j
sakTw7e8JUt73rxQGOuQjH/t0R0+KRoPpzofetqujPVD2z9jWWD4xX0GDSmmnbQXQS+5P3TZ7kY5
wewIWAWu82mFDc0RclEUylYkBrmOPWo3kfG8YZ2nV4cLXsbe8Nj3fPP9kwBPIFNw3mdxENZ+Im1s
h6WvdNng8bj6EaxY70mAKRagkXrI2DeaF45RdbSL9DjlZmE2rF3GOmuBmkRPdm/e355gEM7412oq
3d0GcRTfHqSY6fyGr/MyuUFpHIQesU0Lu9OPfXmWojJRMhznOxajRCqZ+OLPScI+qObL5ZXp7+Ae
Ud27sfVnmUPYnqzErfPLlx8eHASS0pdWfxr61r2ZGuSlChAY7NEUk7eQSoiIiWt5241ehaS2MLz6
4PN3RU6o1DlKLri5X2dHYe86eKmIA3HOAaBNcVvutA7kYsfyk79G9j+wAp5djXjPujv30ZpySkx8
8BaUBeWZQI9mq0P112/s1fSPTHR3OdWTLylwm6ZnUqz4fu2rUHNXLeCy7Q20svzyaFaVXTLjqa37
SFNMeAPg7DinzlOKcyVTCLGqdMVsDCfzCG5JMVPyV//lplP+umOlKwlyqiqIQs+f+XaHqzO1/MWj
T49tppbs7B4a7PMJjKF1UICBllLX5DXZXS1v33/xtv3rx5h/RqCiRAKl+5jxFZn3xENjTk+h7Lhb
+lNmM9UOK1Oag6SwwK5OUzkF3sw2vU7UcfmhxRsbo2agCouX5XxH6XedxRVciV8mnISiNWzuej0T
YFjC7oXiwdTyIPZPX8DnjbSZhfSca6ofXypBta1QDdo+ErUMCbBfGQfLM8dZulCBY6iuU1LGu+cg
0S+kkVtl+yDg9zRd2fqTHBWSpsnhmr5aRuuREnc36pdfoY1yTP5JKCQFtlv24p9wKP2Ob705SWuZ
FHUlAEhySX664ZtWjA/XgvabUAblBiJAjSF+KjfnqJVsnnv14KfnAr6c9tKJDtD4cAZNrDjePsE+
rAVMEeRDr91HyMWG/ghPyggTQOyXiitvC/Ke6IVQ8kN129OJZ37/BJv5075X9su1kDKiLv1vjNck
E0And8HKjQjxYslV7HmOEeaD90OtvaVpFQLZZdc4O3V8orrwrYFIqAXCqyPCg0UqIAEawm1niCd0
nLpicaojGCwls0afTETre2K7T+QV5BZzknh1qUxNi7y/kq/Ifx2CO/87ltenLdmlj99OtcM3kKfq
rUr8HQXheohVr4uMkFaH1k6Bw6HEee9LUjc3fIYx+Mnn+utaZzydfo8DS79CFd09jvh7zRvyfWgw
n/sN3M3lQr/GoYsK2qMBsF1mBcE0rLMDA3L6khkWLWt3CbQnnSAfRJzlFd8hWr4rJ5Q7Lv3+xJu/
vf6nBx0LmDpTh8+0ksdGUuMUcd0t3F5FQYqfxlzrlxu23NVAngKcnOUNDLPyD/nhfg5Q/Yfh5QFj
xLaG25jP11wLa4NKLSFjJ46wQPjiZiOpkX212oePR4pWnfwgtVF9T+CARM9eT/rifm3ZdNruZSgN
v3FgCyT3H/6+XgtvcAE7US9JQhA4izkZ+9bBeRtVupEjRMhdQuIqjpFFRT3PyGz6iOyETH04RCe9
8KfrEdVBo783ZAK2n32iLIAHtNQ8GqN+phgxo3NiJ+5dSFB6JUH0X8uf2kmo02fnwTV9qpT7U9GT
d+AfOiEGokQ83jsW7DgLVl/1DALGeRiFLTp9KNNA6lTeb14gN+dEz56Hu9tKdkYZaDSMnTTWwIyx
UzJyWBp5gOeFhJTpioTRuMfSsQYAsNw7sEezNzueLtEgRZ3CKByg6xOZBPFoLMsjLq4nMco4U66S
Tv6958RhY1wgPCAhgEoI+hga3VbFmvt0Y3UsJ8xsHCX1bUZzl3Va9jSN/A5l1xKkAyFacFosBPqb
yXDkVuppuKH4yYH9mdjktoKNtO3XYGFJwzf7i7Rata0c1puH7TXTbOzdzQAyVYKT4YQYt3WaBIqy
/IJXm2GEay2VIZSROKTGhnH4SWDh6tCNmJPjS2335XjHf3/O3Jo5rrPbLxkGUKhwokK5ZQlfAScm
BMicmAzP+aMat+Rrnzi63KFx8HG6nbB+OTgA9MHKm5uI1PQubdUqljP2ZOsslrciYfxShFdQKG9q
N10ghKBWD99yd8hOyyjMsqoJbRSpxDghZW2BR5qcLqV5t4yjQxO9GEexB1jz85dIwR7u3N94NHT+
c7G/dbGaBIo4PiSuKWUYhL1GEpX1bwQU9Hj9bCkXHeNCibIGrJ4d+M8Z/GDmbcYmcxU4Gzxjh7zK
Z9uMNdFxYqXb9Bn06+TVQqocerHZ0k4sb7qH8HqgV3UuhlGbYgZ9OmEgoRJJPfNrc3ff5DQBef9t
7r7Hj203u8uFF2qszKqx1YICOyd3hsGWWDNZYp715REUMAPLL2Y0iURkawekqeE6Kzv7EeTAo5St
b2+q31oQiDkKKEO43IiHQdb42MY94voAEV9Xw+X2IDVtLRDwqmEMzChwKz8LYySRG/PgB+15wfV9
nhlszrtoeWDkK5nGKVuX9USFsRfR2s8VB9HVclQ6bFL1EGei89jhspjY28fSmhAcWxuFhJTa5evz
RKs/b98rK3JoFAAlYWsltU65feEn9tF1IUi2/GSZr2e2/a56kl9pApPEzVXr9nKV2xZZgpTTXrx7
fcoOLrBLkJSygAVCcB0oyUuS7ePtx7+CJfDlrvdmlUhrTFmQ+VgYRKuhsiaNb8BUsMIbmuwvShaP
KHWkOmV7NNolvBQKFs/U4TJnCLSzRkWRH6ZK9pjfpjOlyf5np13mrKVV9bmcwRXvNau5gtyf/Jj6
jHcpcWwOrdI7Yi9oggT5Anqvctj+1U9qelxN1IzGOP/JjfBXFiqmJiMwf1vULQD5ST2qKOGfqiMd
4jbbEDm4sbqoW5le5KRCv3u81d2eJRbZhVNTSCpCXdRKfcQRepMHmgdauDlP/J5CZ7GDxJ6OboDX
h8W2PtfV7hIVflIUFFwwxMz99jTgNbPwrsET/v+xAgH1ARWuXBU/OhnCwz7iycMVHdyW0ZvmHfz3
4mRRF5YqtC6wk7j0gkWuWVV1Yd5PDjEZoZmsXbmZhvrWl7NJDar6Z/3FN+QvTvAEe/v/pRLx2rJf
D4rreQAd/ruX9dMG8rfPYayw+clc6mCwI9STd+H/YzrrneDKCt6JOgLU7RizIl4Ut5cPjuwtLaBo
8/HXqHYzrb1GlCuWZcdA7wdQY42PKVuA0ADRNGi3k4EGGh0yJADpd5GOud6eR4SBAZxNlVUCuEF+
nxIfJgQecelsQ3zIKy8rN590F17PlN4xbEfm1OEy4uTgvf7wWp5ooU+HnHt6KbhfjUwmq9NrhqyC
dCpG4AF9nECXyFiPWV6oQCSX2PFBZX0ukJA2H1vpNXxokN67WZIdx1I9T+L/J+2pc/QblHMwtHd8
ySm67pZTscX3vMzKJjHbVK9taAOhlx+WLoUvMqHz+vTiR9ex7R3X71guMuR1y87Hv2ZjbOAe68D7
Df1ViDeY88q3lxjXPo786LyAtacFK2o8PVD8evW2crGgZLyJa9i9a3UvrDak3UB95qEUoIzcV94m
RPrVAoWz5ShDKCr7lfBVyeMlNAaU/gxTpllKA4V2RdXq0nZOxk5/9I6Lg6KEsXMXN6gRJoT1lFsq
PtrNhcmznZWUM0S5Q1KbiudQ4mUfYBoH9/li8zDIo8CMTcm2WCZqkI+jeLWn0Blf+41HrcDZr57I
5ARh5hXE15WmEj4rB7NwRyD74jbCtZcNcizhcNc73O0ZHiaaPMhBEZQ2doGuy0RyJiHn9sIplZ1p
p4IdYF3umvDbAy7X4+R8DBwA5z0/kX/OJ1YxwCZyt6FqCKU/d+QYMvPI0RDAjOQa+OxlNFYdH5cu
f1bzhAyh6Aa2Xm9ywkF07drZPPVlEzU8bCnln9pRfx+qPdPHsFKedSxjKFQ5nYLO6VNPQ9bdHQ0Q
/K4ZrWF9/As+lWgOCLyI3zGeQr8V0w4ZUSUrqHlzI/yP5Us0oj9hsch1aJKcS+9WyXfq2WP1giLE
yP4YpfRngM9hQ/Db3GKGFliT0qIlSiSG6q1H0mum8kbhxd3xosHF7iGKXPDqY5o5JkkkraWELYQ9
yRKfj7vKWVUlGlxJrVf3sG8g4C+plG/tppRKKYZNgIIn96jQAIM8uX+8v13dxWOjItielNjGcz9V
0oOMEuIThXilm+taalobsYEYCPUw1cleFQ6kKpaJk+cJnENhe8e66aEiWqwdQ+IhiAMnnxkxisoZ
sLv4UmpXpVTUPH89OwGLPSEXB/tiAFuWKKJaUkc8qysat573peWH4E1/VWvbOmIysbJvuB2C/2iQ
EfB7mofQaa4wS6bxIUV5OfdLS3ET0Sa1dVzFg8fp/exrnNewc7NSzFG7TJy/8X+a+sPEM2+bm81K
NjxdAKGcCs1Rs69wj2Pypvn0JYjkZx3/BRPAuQfX7RNGw9P+GyLoxCQNDphRErdENx5pV0bqJfFY
ZszDGvGsw2VE+RcP5/ldee/w7Y0vA+FS35cqORFrZHf+IbH4N2ed//h8GmiqgLSft+rYZZXUPRXQ
cWaVX9xVtM5MdOflq/n4vF6swllM8z+BzgtuMClbD8jwej7W34DqsPYgPvFfc4YLk8Dc3cRDfP8N
Tt0JR826xWyM80D5sEjdBEyorjCxVkBRNQshSWFAxb4YeryWFH7qgJPY8qaA7ffhz2lfuBevpFJt
oZxHmeNOavxiz6GPgcqs+j7KwC42Xfd1hLd8kCO9VlZbmjLFZP5R5Lybkl6KYf36hh452IWx2HEF
on+cX9MIPzZN7ILxxWXzQo4/M8Mrs6hkCMNuRHsjr0rNHTEu1gUt/x+MjvUn4L0M/+abUtmchZTF
bu6Got72sZHWEBHDCj5nN9c5+yzitoIp0qk49tOidA/pxcYeC2xKB/7FA2JSSH0t1V0zvsupnneL
rN7FPUim+ApyvTe3Coo6rOtJMrH2JPLJ9G4/X0ky6gsLmjK9HuXAeXij3O7EsTxeyRfHSkEl4VpB
//f6G/UPATaip8SD1BEQIcWP7nkhBI741ogl9g7xDwRNygNIMN0H5onkc5R0tROfaFSrf9sKcnwv
4l3h1YnwLhsNv8IaavwgDMZJAt9dNF8yeiwsrF0YjEJZr9hwgMoU2sHbnW0suKDEJQauUa0JUI8J
p9DOJ5zBvjroLwOrfxtn/jFLVLRSx+/+iorLa9mg1xiRXhTIgvNY834gIsuKGbe0CCSJ4GwSctQW
hTYl6lXZ8EJPMgPkDCc0MPzAz1I58x7O2BAOQbE/YiU2iByWGHOBo0gfc5rf5IoXpOmSsRhOlR1u
4ltwTMbFwbMhw3+AnSj5gtlNDRvjX4jGipLHI3L9rw5s7L0gV5NmkXQ3MG+MB6kyyM3EIldYVkJE
FCHdlMqa6bD9w4KRG4ocSaYBi2X6/mPks2aIls55NdWwdGt/Nk8jAet2F+j6EASG2wl/rVs+02co
pceHuoWpCpCodKjkCFg9HbvVw+hUpbr9N2XKrRuF1KQM+p1hCFa2+7ZX655tMvXyAf48St/GAt3S
wbZ/N7fPt4NaZpLyyzDLmS+JLqpgmmMMSMPZ+3s74VcntBcY4H3k6DkRJzDCSKLnUSmimkoAJSDv
1IVE4BZbzzm4txI0SHfJ03RaHXIs5asKTqTo+o6hVqY0DhS/OCUBH/+r68h4M5Vdu8luilVgEm4T
72PDRfZvcUhFjtZBuksRuEti0G307X3xkpmNuLyE07eZmlirrH2cEcienqFMRtGsVy8OsB9KmNkA
k60W8cJmVJwrltOflsdcsDLelFG2Vw4lzPtdIbAAgr5rTTKJM2vMNSsnhpc8kGipafbbPBUlPLfG
9YDaQzVD4J2gEmEKtktEhOvM5+hQEW8XHyqUfaOKHD7w16wA8SN7ybZIA6AO2SLtiz43DG8drEDi
+cTzXDghaIr1xw3sgO9SEbCBrj5UaOZL0iCFuqgaVOTAo/cmdmFScgLFkUJOSVxhA5PLYcLtSdhb
opouXhRvfSNa6xgVzctbu95L80kMxpIkBfbI0HUkbXfmCDnJiMNBXS06GiEP13WUswYwxkoLri/W
HWx6dtTbvsKDNVnAJjVDTLf36qGnNZFtbGJ/3tbj3R8+wZC3fnxttr6wxgMi6tI1IPv7ptmGdBYC
VO8FD7ASoNT3GjRs7zKiFjxfbldQfAN7APUti9xefT62ctfPZKX9+bR6MNdtP4F3bNTI4FvVqn8U
TIlkXSY1co3VNAZuRFhWbX1C/U2ibseARPCd1tYgIWtmfIVJF2fUP2//+7KdwdvVu06Iz5inI8Ud
CXx29qhs5+rw9IZE/J07brGy7NR713GnXcEVnc54AJE/5qA3fXUwGQOnfMFadO7VpmNAgH+wRtz5
+MOLPnkM0DDTjMqo9DoAvsJ+sjcayT+B9UfRK6SrgB+jy7mca/5zrXZpnN1an++d7Im6OSVwWxp5
GDU38P3hjNHX/p4sI3YDGMncYejuHqMTx5/P1lqXok92Tl9HbRsFhrmZdftXM+0kDFc+SbJH8HGa
O+KZjS5I0Ud4xwerTPjp+n5KBaYi6ErvjTOgDebR1NMmvVm0YYw1EWQ0mCCL96ULwd7cRebIlC/z
B9dPqNB+qefYWMFJ0r2Qh8zHjQ6d9IO4bXe8qwBU5fLyWJHdGdJxihIQJjRqmr+qIsHJdsR6FlCW
wPPXSFzrGkEbqIsLF57XW4vZhsUb5EuAVu1qUKciokkpHv/W4WmFWXzGpsxBWN7eRTJagix7rVpo
Wamr8OXXKCu0SbBbiyZ67UvNBhLwG+5XztRwwoHrRfSXEDiOiyv/8zjtjOHULD6naSaWyQekV6Ig
nUX/dHijXxJRg/DyRwwB3/PXiuWC1gW5KmHIhDsjTTqZjNAjRDWqjcIBU7+rtxdbL9Nd+v1mBRAe
IgDFZljWO33aGcCbEApwI/JHZpCnUnpfk0eMLgQI0+v2y8PxBdtchrtbBe6M/QnFfNEw91w0DEXM
ZRLILjEHVWzWhhCCS8lzDn7LJ+Zsz9BKpodj71yi7iPaYPMqP8Xvtqokks29UVSmtq74svG+JTMm
LTysniAgw8W1c/f6gEThd0XKzIVTUefb4NyL8BCPFqPAnQuBUaZvVSmzW1/qHnd6SdvwTwdRxqnC
Sys8300ey8f9kYEY8UTDjjq8kM5CqaoZeqkH8JQW0l+Lksft5ZXTCF6LvM1BMcazN9m1btFfYtCl
YcKVXdyfkLYt47n9JcZ9aj6+eyajLxbuNkB60XZ/bhT6M6q/j9ABVOg0K7Qj4zTbaFa1awkBgRAY
XJuv7c3NH0S7p3UoP0FHgxDpEt5XWSiNTfnaKxbBR+c+zs7KZJY3lrblXOHeM17uMKtNC3Q1tb+Z
fUKghnjn3fUjj1W91Z6kedeIhc1XFuIm5UMPGY/99+FQJQO1BILCssSCNiQMXXC9E/FLqYlTnMI2
kRrbEjrWflNlaHPy0sBz56BuIholwHW7bV//GfrYXFlzSELcvTRhjXlOUfZ0QWeD4YN18dof/yng
9FDzLSlSxE5MdAHcy/lyFT4Wu0k0g1CS0N3LwEMSwq1s0y9WqLV8rbuV41srQQkvdxW7ePLGtx2M
D9rbwYNBAHV8ULMdlOTejzz69l9MKqpB8JCC3seFhdVmqrfiAOUMsesDvR9QnKT0eHRueTh4K/Ue
yLqsHCFC5mZl9Tu/LhhgdF1CMuGdbJONCI9BYMzLb6Q5YAPVwRsIiZ8H106iMoQTcsELSTztfB5M
6JRvYW69B/lc8uwcKdREoqaygzufE04dcF46EtjVbY1UnLvL7Qhvbw/4zLtASSKySXLJtMB+gGlj
3prNYojAA9QQ3pvjIYV7v8Lp2Rf822GOgu9kne3N5cNNO/SpdqvBFm9FwR1XQ60tCrCm1oOWmGrB
A5CBvdKx1kkFFZO6eeLstIH5Onb/tMtVM/fxvKsdbbPQuV3QXNGcnj1PfyVek+rhaiJwNaacyZxy
GMTN+D2w00p5st5cV6XEOg54P9VgbItatIbCYBdrns273iUSa4wF6I3wWAzVlVaHtl5f10ML3k9k
1ENZbbq97C91bFh1m9LVEzkKX80avfovVCuUK8xyGxM19+TxK35Zp9weyx3Q0cSvz80MinKEloV8
hbvbdLa/v39Th+x7k1WWUGEzThKGsCTuf6uRCzoz0lmYBHVFDaU3UiQ2yib1W2HGTfuFuhzOqvAW
ySzZzslerOQQ5pMfNZWJJBQNS2UJhjuR7ABC3N3E2mwQTkMaorashb49nEfH+4R8pnYCsXYCX7Nl
RcO7/xtKb8Qmqa0+I+Bha3T6krfzRZXhH8XXpm5la+2E3nc4jrlWLv6SrnUHIuKl3jwVu0VNXIDy
QSnDCr/wCblHnaRaCVyWrhBNdKixzPFBD4mpawZDL8xjsKpoP5/ywdg50HNiVVOekuD65SjRa6ta
gxUn1dQjzuG3eFjGYtVFXgj8OF/GjRKMvqMXu0LIkzR7/RLZpjG+TUaGLJZt1BsU4HUT1kRnOoO5
vmXjtBt25wv7kegCeLyh9y7D1zmp4ocqKvla6uLiStAhqh8fETNRC1/ECVtQewuruiaerEciv/FR
Py0JfkhnPOpaQOvDX66QQyGqqOnAfnjXdgzPRTOMCegvnO6Ra9KFHeDtlo6swP9pn8gq9vafc3eo
QOVOWTQZphL9lW10WSB6hF6jyFAH6Vut4lUkbAY11r5fTqf8tit6ELMENz4CnSNn9OJ+JxJ0+kIa
FQgvdQVjeUDogUYjLKAujd4zzzMJoELVzi6zeXGpzgxJ58LmDniivQsp9JghgU+99i0+S0h8e7QM
9BsFRlz2gNChwsxBJRdaS3apFudG6JAvVp39Y/yLEsZuL4FnJ24pBUcwDupZ9pyd6s5QXzOJkRHR
DQXAFSMCCPI3fS6T2HeRsoOmeUhepJRoOXw2yXELEFfMMQqspBKS0Ms+MV1d9U2PUiUGvcONk8w7
BFTs/mvPM3WJJLBholPcDAQsk/r6d41qyPpuvSZHxLO2VZ2UfNioW4lv9Vp2jVoWHcQRAkgTLT7Y
XrA6+HLKgBxPiKBOqKWt3Dk06Z9gmPOU9HMkcWCCVOjtaJcZIXGeSu+SkJNgnnK+SKW0BbC99fm6
qZJ/S+2s+y98eFe/MJK9QavwD/HzJ+6ONIEmIVB5dy/q1G+dd+Ek9CAHbxPsK2cyGQwQmxTLoj45
03lLb0aF6IPTbyBPqmuHB33BwhetA/X9bbnybSZiKAxrqS3pawXm1eISVsSISeQdWeF66/AD+MBG
vy7xrMuATeX5n92H7rfEXwSsyDqNck+oi6AZkl2U/kiVVkjJ3I561KG0KLdCfD/DpgG2TuDcM1VU
IiV5iQuMRysQxrLIGRAbeTjja/rzzBp7e03ov3tfVRB/8okrKdwHdkKCWg6KphvhwMKfMVS6t6Td
W19eyUKGkgSHeUiyJ8/IzG1v4z1JCLCOw1olTzQBZ7Flm6YZmf0jYPtKrpP0puAaIaI5MtX52KjY
t6dKz8fZKNB27IaXhFujZSX3z9/di9BLaajNvKe9w/NmOCYXJinlc05BzRaOixSbKJ1NRcZXRiqq
Mt5gwgpZwRh8HmqDjy27eFsDBLoZqdov+5U8ZprBST8pndgpr/7fJB1MGgopf6G5r9Op2BcLcwNz
g/PFbieq2HdrlOxyUGjAUuwdizHME1jfCPwlf8K27BrauTnT+h3X91ZvOrpHzycYGf1ZQGxkhJLU
WvrHuPbBHTkEmZzMFFgE0LCK5fvlRRZiu92OgvTZB+h31HSsoY5gt1Wk8cDJHDWmhAW4iesvhbxL
Dlu6c3vsqnPZHmn5FPI9ozLFJpP49u4aJQDUCoaGMkTak3s6b2C1CSZHs4n/gdT3kXJt9aMq+SpG
zISsN1ntB3pPKRr6ct5+2pL71NtMj5LUMPh4IKAHqddF3fuIXvY1znpAMDnbafeeG4I7cAFKwJYE
/vpbjxHSbFQVQ/jb0KTAc9mGxPo4M8TblAC61yCouuN7Wcp0+v2TAkrWIfLJ5lZmS5Ev17bPI04S
4nlsjVZ1gunN8aHP5h8OE12Vk1FZDJD11j9drrkSTy1oXagvCUYFB0YzttUBBc8K9l96b5F7G3ER
q1WZ2B5+FeytIAl2wsKEg7T5VXQGo9T5OfqvTUyPBe3S/eRTlRNq9XBZdOA6h+Cg5XbsPqGwAjX7
nJqoCfJFox3rStLWjlfU1TwMhYx70pfHE7V0bTjkp1MtZXOpIkENupdxV4fIIkAmwpCqLO+B51U/
WiPR2+7AAauUPGzSHs+/saeKK3HlJ9Y03N0Tne5//gLLaD1O89erubd8tL/taWNBTpBWU7rYamxU
767ksEPGid6ENyn+64wKpGjXEBHSjLiVyTeuSV6beS74uDvC0ThmqjdeJ4/R4mbbwo2KPjvnOJBi
jHeAmjmRdkxU/tco5snZAH4vAyyWEFtD49zobpMnRgSxG+Io8b5fBQnoIk0UbmseSwb2PnWwoAua
zuP1UJFAI3mMwR4Uktw6jSnbxqR8NcTOwX4yWKxUTlfb4lHPTN8P6SiEbu9GJx9O0bEa16/Xwc3Q
vAArt/sNIOQuixHAY7AgLTSHcNA9gr9eqqAXidUzO+Z/jOB1G5a4lCditH7OpfPlhMZMD2IqxQxN
Om8xvOMS8rmNqQfvN9amY3JcwG7TD9LnLQeyIvfgulxchEaJwxOjWimai3XUf5m7ZACfUSoIbRBE
t89K7R4qXdYP+CdEaHwFrBGgwUlUpmNW967PCKUGD0apdEnLEaizyHDJLQculoNcRYZcyEYwSC9j
9uxsNitKrkSUTeD6pm8k8wPq1ntpOGffihFSEa+qN4zrRZs8jydia1lSC+oETKFN7DdI+juprADy
lbt+BmABtzP3/e7ZQssYqBLxeMZQzIh5o7rUWdWUIG/SXKCzhlicI/jsj+7SuYiJKQj89oLYTsbv
clAq/4zF6ot1w9EhshZRwIRFftrOQA1g6To00WxyhJ1nzXQl5Lx6zVFjwSvCYcICKqv0ikD/H75Z
/1rITup409mG3C7fgnIjVE89O7eDSGc8HS2fV3fI5W1C/qE2HxxuswL7HUt/69So6ouANP6yVO7w
PFcwxggM/fzoxcNEp3CrHbFjDk6sFDgL+W5cIekX2/LzDGgePIO5Haizs5foLKIyFeYOACyJ8zFR
oBVxSoteGbg3ce9J9RkoC5u4qgijBeWQ+U+/QJq0QlKNBh68sZOjNBU2ETn3qtcZijtU9A167PyZ
01Hb0FcTgvCgfQovDW2VpW7D/80SugCOhrR2O1sRpdjEbq2l8A1osGyTCkGsXvP7ImMR55YtW7sR
y5Z30yjMfcAKG094g1HONd35+c+1+rpwuX9VrmQ2PGeDTQBKVI+ZRdn4jWRFnM/cGQLdQucoPEf2
w63M2TWQI6XVn/OZhxgnkBqbVNUReoh3YV6Jj1xzQGzzRGroXxZL4TPw0bAVsg3S0zOxjXMSVcAX
/6Xvhw0CxYP1gje7T3nyfEDFQYvBufC0EGujVvLuNysTBjFtbDvmIwJKmqJH7IPPTVv/8lTUpzYK
dtbrq3hKVAnGYEGfELgBAYtFzbjgi9MmKrLUcByKCafFwDNdTnvY6v/7YS6ItSZ4gk3yS0QI5CUI
NTku4FmV+ZtbB8AacHi8JrkUtRNTwazKdgP/m4M7TJrTAl4FpaOiZZFbozqF14zVZuIKX0gh3ytJ
t7y3flH5DhFZaz40aUZtFdk17EMbUG3cqDrsmUqRvs+HQ3TuHrIAZMBQSJeNXKX7iJS01mDj5ByH
m67O8IAhpY3zaBwXHW0yX5SHpniwiwabmI1L7n4f1A0lVpse6hgJALWEHvFMyNBry/rAUPs4wBRd
NR20f7Imklcp2DsgnHUdfwdFv3ueZi3WoM0PxrFtC9ha1l5UAxGtP+WE9gEsQigIq5IQSL0qbU0L
zMhexzwRGtD3VRWZfts59lrl/VGCg9OrshO4pZ/3PIBvm2h6P8oML+FFDmsK6fgCaTJU11DGu+4n
dT2QQAyvzQHtkZzJXQKk7sc+MRwLy056txmnb0RfS5cMZLH7n/JnPFJiCO73KpIPQPZgu3SvDIsv
1nfoJs+OcMNxxUHB3wGL4VwmJ/a+7syuttSB93asDthzTutPaoU+jA6wEoDs3NsCuPXFam0cAYvP
I+deIXNKY6RxibHpGufHWtmXUX9BJtmqJ0o616w4yb4mxibvbUDUCaYq+UtrwS594jkmMgx4E6lw
hCBngcJep18ssyku48p6Rrv0tS4OHQFb9KPTG0XYCHA0ZTOkj63iboW7xMxNQOyFLbOLl70he22X
c/gocy5jTieSj5uAksa7IVlGZSLxn42s8B9dxj3+pO8MpLYqNix1ovBi3bsH1OjFgQggP9qWaumn
Jdq2VKcSRmfEjDcrT0Ud5wuoqveV9Emtz88ZmsW9PzrhQIt1OUeTTcpo4yS9FrUDc2KEDWD/kNxm
I9Wjb5BNQRjl+ZfBtjbIIVYXAsDYIOPqGHaps+uivVF+Sdu72wFupnDmOYxDLpPSznZ0OyLZ+fAo
3g75t/bZtIHjFARg87qz7VsbeO+n7lfqFebir0whY7FrAQbIZikp8UZaJDqM561+dR579lVf44lx
XVaGckhg+UJLjmGrPk5lNk3QGAODpuDUfIDla1qCNNOPfZgJi4gHnDd164NGglssVw69d3ztPW6b
qQSGPj6FgGtOg6hdQRlRPtZUPNyTtgh4zrhCD2RR6TAV+ABikdTu8rNuN46FwFSdvjdPTDzc9es3
oHhN6EidmDL391tj8O+AaC2R0jfzg2TcUnOrnPgI7/Ol/p1vacMVJihFIOCaf0jo2/kQHTcyZASn
KVGWHnMbl1WAUdEyn4AeVG9P6ER75dyIz25aEs7LWNBR6J/DMf+URDYKXBuhL0Rq48918UqK73j6
YnRLevwNt1sQzvDaDhJv7vKQpRsSyRChpw2MmV3KikPbNMt0eKwH/MoX4JEwfT7cewV5uSbgIDCg
Mgr1P9HlLFYGKHW9rBO7HxyupyGaaQ6rFfnswOXtUowOJoLk9Lpf5mjhZ3+Op5dfF8C2AbEd1f/9
H8m+j374Srig9sONju3D2mzSAI8TMgBm8L/9hVeXWyr02KCKuc5gZAfe8FXRTTngfqkyM8GtrYXJ
6n55tP01UJdC8MypshooiG8ILBz7x2R8A9+jNQNYVqrz4PmfxlobOg6mESLGChCRFxI9hUlTIkSJ
I073odDG763FZ0kBXL1tpnp16WoRBZLhB4POuFoKv2nc2l8lF+uIKInHRQAVS9F8uuUO+nbpO+MK
m1gy0HiZFuPFV+xQ95xmG5WMayURB4fKfgjo0v06FqNKOEf1X3Y79vPkqUC1znlgiqQ1UkFU/XnW
AItLYvU3yB9/be4XZLYyBdpq4jEWE/oVejEobw5H7XRaiLlAULasX8ZjBLNoIwQnJBTNSlz3DukW
bMpX5afstCb2/qiwgPFDqMaSElTafdkaS3q1p7GpcguwugVe5DAorb29mNBNFeOpFSDB6Q8hd66H
9S/UxF5xARx6K/cm6Rm3dHi7FdbQeYjEYYaVm/BtoiiGP1rbjWeKVLYxVMqVD+3lAM3Qc1Et/g/R
QaXkiDyPZoepSNnyhesW+6Yg0v0VW1smRGLxtm+D7fTgqdgjrwcgHU4IZRfPcrr/XRYkvkyuH0U8
MXjka87loJZyTxi8SDcxeBUF4c03mXS91kpHPNWOcV1E195D9klGKXodos5G1PMUondpl/9CB4a9
CKQHAXpNbMJ10Yp5vJL3EcVvDs+SU3zY77XzngGhHvlRkbsjThhK3QreIfARtwJEhL/CFr0m1d0k
DI7VzjPtBsdZk1Nf3kWECO9JpkFgjj+sY7UHQXkKrpHjkgjhKXRttRwv11ruhwEHa0m4i/J28Q1Z
q8ihjIWbqo9JefLZvn4Sl6zajX/zEAWVWuU/bzp0ijJtorIgZd3aPCVcvlbdqo0AGKNvd1MOy2t2
zlD4TH/4BEmVE9VQmhG3hKtiyDpxykFx9x++AMm7ohDDFb3NdcFA/qzq1dukqWo3AmA+vqlX1UEI
qKuNONQhJFWpJEezmcoSS/890uQ65isZzOgF0zjQiyo6W0KRtND5NAHCou5WpygRK1iaWm94NKXG
eXfLu1VyQH4AXf6QJzBF6x1UEX/gU7voyBdlwxZrMJRWt9b4Enrkpt94LT+3uZrVBR5OyWk72EZ2
Ixqz2rF0lOnFNnJLBt7p4qoF3ob86OQ53ULD7GzUFJNuz/6p7+0lyNYt+re2XqU3WDz6c6JeClmi
apGAiiJzx/Rmr+cvhMWYu3D3Vwo+wSrihI7l6AZIVWDnA+SFPH3dWLYfDD2NMJ7TOoYHtTP8XcwC
iViwo8l2hgH7TsQwTCjkvYFPLy0Z/fvuDnQApqw+sJfNmR3xiQdiBCAnbj1kSCjxY160nMfy9JeP
1obWaf4HmR/EUQRaRcbmBHB4JLRL5H2fEY15eBkcdIIDNKVXEk3uTLdhGrv2w7xZBcSuIyTeSE8O
K677/bET9DVJO8WcOkvRccpG7I4nke7AITQdPBJalrOQBtrC4t4zQ0pMB2E1AgorVtVJXpWD1sNs
PU+PqNyri08yiS+ZIsGhR6FPlWbXcxjPi7p4diC5g8P0p1fyb9KaxqUwcaVLOQuIWTNwxtxhyIYe
Z2m4Ki+K7G5RQ2WtZlSe2zAdflsTcb/6u7zuZKs8jQasVFkPqscemdWcA0b1twK9GjNaG0jcpcMd
vQ1nFF4Bwc7ESF++Wzfv4RxxX+nB/YlxUI+EozfeRg9AV8WtvSgDvfVmJa8fE43NEQG9bPBZBBYW
Gd3cVSf1BvQaG6VUZn5gfYt5Rv91PgHeHOwOUQsXa/nyGHGu4qPo6r41MZu1WBQeF/0e5wpAtz8K
j8HvdAl+mnqyeipJG8ok2rOTVQlIqUgriJt3fhpx2gU4v1zMjRJPIJvGmIOlTWkJ2fqQmhuz1Bgj
SAnAM/QFdxfJbWRRe/JaCSnYlGFI6xjeGmFsN109WjEa4dySTboQx/em1RQxvw/8jSJl6ixeDQ/B
c5lmS+pRUgXjLj3geyeqwsf/Wa7eFCUAPwSEDtecdN0Vj7GMZCbS8adyCizI2Ej3r6UPukjg+syW
uy6os7EmkhJz+503qgF6OecofJWHNbtYgQwW3ZraeYjSxqmCGDJk0zTM0ta08yuHF/eD+l5Qg7ji
HH97NIRjV4kHFpNSr2jPYGqszTTZXCF4gQq8LOGGgpKB+DGEgf0TxzhPjjaesmAD01DCcuhFyGAx
BQRrUzSr5y2d9ESP+IYrfokSBTAgiqVwSfB6WqCIKmGjMjnM1pXIxlNA/To9X/QawrVPlsO+v4dx
95GTqgu76tJ6mnyTloBiks6o1+wG+OVTI+fcnvk46dxGMh7mpdQH+6n5mc1qqMd9IKNrwx1pNx3/
NFuWx/dNdtc1aL7XAnmejOC2Pe4N13l9IinTMVUfOEPW3GU/qweUQI38dTjyvbelJikVCAMU0sXu
DCuTcVk4zPU7WXInb/wY37FOdSVipHLS1zfkq8X1YY5q3NkzBp7ij2C00pTwDdDIwXiLrapsqi3O
HwX50cpD8ofYYEif7KVnEYoMDVuYOixQHrgT+94KjKp/WDMmBQcyBa6yvCc+CD4Qy5/jT2COehBN
nFTxTd2EFVYkBpAdt5Ptbz1Zg86yyQsjpVLhJmBhhkHz5q62Lzupjb6NTzTsiBcHXbZ3kIS9k9wt
THD2cacAOLrTpyPdjVz6AIIrdPNcw+A2kZDhhQ6g+pRzWNovGHh2B0X9J4vVxEdAaB0GxBa5zH3a
ZcM2epHUJUNA8Dif8kTvC9XydiFSQ5KsvORvs3aY8yGu15vQlljeNY3qRUrIFj8dDQOxhlmvI5rO
npyyxApyENSf66AO4FphvhHOPpaC9FXrayGWnhHosRtBWeZwzfIJ+sA8UmuPwUBTJc72kqHI8u6O
mb5ULPXgxQ74QLGl4XmpjRIZTsc75j4wMNfkywHilDtthK1lMICHLqv+Hg5oE+AYKAZhWz2cFtdE
uL2dG1HYGIbmoJeBRHcmT8ICTYT9aZv58k10+tgMJLQClfecVu5ZqVxtAQ4AuPr7bx/UBqjRe9cc
CAPO8sV+atDV0fvIMnqgxSDV0hab7iT/Epkz9etwPiF6HdCzV8ukOIViKAv3NpB2Uyl+CbFG/LO7
DppiAIDjEryEOXjBPPzLZm2cpiMMmYjUhvxrFg+9CvDukhstWVPSudVKsTVyNbg8ZS3VRQhBZOTN
B7HQzb+4yqul8Jh4TCX57E2oZp8gAypLgXxidaUTTnNJPxll5DRHK1TEdJg3ymO6R5GlKV1/NqFQ
1yHEcAeoR9QB7BvUbGHTB8Pp7maVD6E99aYqyvQr4MrTFQpVKLYkNw9Ru48iEla5UMmD2X2w9CAA
uw26iJad7eVWzklfAQTR5aVXBi4HUAYUNeS4pgxuug0Iyn9fJWgCmUGdeaXqEAxBbR/7y9XmC93Z
fut69HiW5zryhymJH4Wy+I/AbsHPhdi+UcSE1heHiITb3tCynBQO3Qte0R8kxsK1d5yyNTw9F1GI
hycHGJH/GgPaL6LsAKPREEu8ZPP+9mrPjFja6ZH59Bqnun/Db+8AHAwyUtCpWBnJvMG2Mi79AzcY
mNU8V2BFEx3EQezix0qpSYt3RSusQcJWqXXavPHwUz/7KGogeKT96vs/RLqYWruMiM6jJQsK/IRF
6Fc4MKFi2ONIgqaDcURLAZ5wvv8QI5hrb8+rUgpGvNH8RKXmfVu8C3/YjmD6L3j2U8eVS6b/EXHl
LhCYF7WNPui75Q0zbGee2HeGRek9EgMhiRyLA+8G3tk2GTib84kmZBezheSc0F3nDndSBEjr7q9r
Jr+wtJx4pzDEl7Y8xA8TS1VigFMKg0Asm4PMDc7E5vQFOIdpAQztGBFiYFyLzAHGs3mJHonI6sHD
QgTZtgU6fUSJfjgEPvROEy07Ar44m2EBqoRuWBVvsCu7l2esSTCKG0yFIqFoFiFQXrLj2qR3FZeO
xTL6j31NbWv2omkt7xOxJju53Y+zCRKBknE+UrNIVy06HtXtAWla8+4fr/nN7l8WtXeWUuDmfBSM
MhLg4HkHitkpz0euC+uZcxA8JJp9L/vTY5va3cFhFmezEBUrr4y4f0d0znKyFI/1FmcUb+Qmh3jV
sAXoqZ1igo1jvklpfDB4TnZUOZlWG9RkqMwcomcthuA/1B9QVnU+i0sL+tf8yB/T8kiFLFax5JAZ
yot5vG8IT9RunLfWP+zHWJDZ4cGtudObXs8YUZn+xXwQxc/BjzmMbGmuSJEdQdggrVlq9lGCcGET
AavHV8t9qXyNVHH18whlGLiKlu4kEH7r0iIkjNGBfbg0YrjDcFfUVPcIteeS9kVIOFDK01P20rLY
yTd5jhojJ3/c+keCBT2PMLM1Uzh1Hehx56WWyumihPJYOkVEKwPOfuSmHkxXX2dYeexz8WCprGBd
t8jPeBJ1SvvFctlqHaLAOFk0usDeHCK5SEEHmD9ZCenBw7H01VRYiWO2yvFxO5DCD7mGQtazMeox
WIhVIourMqQgEiLwnXz1MgEdoqy/hb5qsSpID/JouK4jVx38r1/JYshhHch0+BA6/J+vacRIzcrB
dZzqP83IfrEymdVaJSTWIzQXxbET8UZkkb5gA388/ErGoq8V5K5+tRfB91ykDpxFXKQz1qkqTOrn
tHwefZkwawvKXlfLabHuEfmAU/5v0bTtZvSGPAeEw9Bpm31WMtVvK0UWdkgZ+wy7eiqFWPJhdp69
R1Fz+76iUZGlBiSoYwji9Rk89Z/8rgeTW8pL2D0Wj1K/fJZ4lmtOCbo6sHQAbW9fOJsePk01ajVG
hMqJgPwgBsOsbRYZbsT61qJomQOnRdJqqu6M9tILZFiVfWM31wMi0Qf/LT7CzRyeWaRg2d7dLY7p
rggEyKqC3sruFYT+9Yg/MFGUGb1q0+JSdloG4fC8ejiC1EGIbuHdnczyF37c9LT/uaJzJNG94jfx
zgOvCZ+WGx6DN+38WSPhnriORsrBAuW/CK7U3cWk0D1KctVRyUl9nYFWWCjh+wuzdhf613G5Yb+O
VppSua+/9WtAwssD7ldqDeyeiD2yEJz4dNFhaPhpCEqN+cklkfT8H5axTwMEl9p0EQUwpfBD4fqR
O8Sdz1tK8k705d9oU+cbNPcZQ9fL3eDJ4aUdXS/z/h5ZEov4E8/bQPa20DcQ7G7s92TgIPi3kTa1
d8ZWTgmlS9Oj+q2+I+aAOpao83zGNlG6y8t7G3IiBKcw+M1HDDMJKyv2FeZqSlNfw3M9Sj1sUmCB
DRzfX+fLxzVkVe1BWIrsMrPu0hrdG1bqTKXHamcRh4pyc3yYb4dDuWFQ+EgixhM4kJBfSDzHoiJ6
7n8X+w37jK8++PjBmwSPLgKkq23bkYFGmNKOwcIlbxApFRpkUlrx9WiNttUW4F4UDxqpGS2mKYeM
XbEyRTLgikXl0BV2Ze4pB5KczQHChSGaSUUWXrH4JnkaOeUfzy0dz26KSVLFuClPM/s8n1ddqWZH
l90OArHyfWDh4NpumZdHe5s11GZGgOtvwsvNK+GODTvWgEQXZC4/bAMD5g4DbYKF/YDoyhYziiU7
ChGUkchN5sjtA/w/xxckp9Jb89z8kA+J2PFaLxdIzOeLr77WsADEq5svnNHOXCn1qP1bF/TxmsM3
erpiSH8fCBbPo73/OYaNwblTyYNz5DOBSsemosW7GRWZdwUgtqYY1b6a23yVXhCugX6cmc29vbd1
UsUhUAmMzsNhuA0t2CRXu1P2i9/7XC61xb5e8cwmcaipHM8Cpz309AsvU1Q8N+LHNLf7BrmTPccz
X0K1GkufSRMtRugrZj1hnKt1ZPWVHg8zjJRYLFT4W2qS/NbKvbaWj/rn9os8XsPokLV3pCyn7bKp
tmF4wnFXG3yWUZ4mQOIZAuSCF17z76kypVZuat6wFBJizg0cO2963mCQIfOmoqa5KA+SW3AbKGDa
NZrBHuNa7RJoeLjdd0DETINpFTxkkGX12u30IWQIFFA0GixgUf02SXhS5P1D6q1jISwDhHvUUiUn
4FLMa3BTjQhsA0nLOahv+PXxR1safU6RtqP2KTyVuW7aJUpNG2+do8AtdBmYxZkicj9OXv8XWjoY
XOlg9mBkj3xE9HRAIa2sF2/+8IScPbewfgFodZTRp4bMy839FSJ3bIRztT5M7qyCYyFNCvtIpofh
wqiHnOLm+9lipdpJFH3ZLa4ExatW9Z9mFMZRVATaVwiIsFSP4NKYo/DEeKVNNw0KpfeTMjX/KdLc
wzEqzrHk4wvC3DF1QBDc6KK2DM/0lYDy17UDvAWWOqJZ/RAMOpnUQ628VkcLbubSVB43FKZMiN8X
B8i9StvSO9mU1noOOMnOw/PO9hTspEnqfMLrxWHuDqoQ9umbE4nFTmYEi9GJZ1MkJidIfRW3ihcO
jwtHYMNwWxSCAmzszkm6GVNwVHsIbACNo/oIUFLNSZqiBP9o2mwu5S44xbgOECeaimPq7WgMx+n+
KGmf/JdHyv5Fg9hpYdcTDxB8aVznZtV7F4P5CjtQ7wb16rsYJhGygefzPQS102f23l3feNZS3ULE
sgSAQl6UdQL+wWwYBmJJv8+4aRxMlMvGbAjMMZFAj1ZkVDprJhfjeCpKT1gHrm3+cpfxwnxnO/U7
mQxpmKc8ngXnGvyJtG4iMANe3SGPHm+WAPfuSwfHjtsL1DT8PDhv/GuCUH3Ci2Fz9iaJJjvVJOqo
NSp3c8+dQJlNKZnfkC8zMpdNCBFls+N2mKv92Z4auSzNGmEYaF0KY5ziOnL2OB+tTyWzg8WGiGPS
VocjWJbl35xNyR/Wr25yJqiZkN98+vY9PKhScWYuL9w4yw8tsJE0mDglVOfkfdP6zZ2vJSJDEVDG
QE2xpYgmCRmwY0/DnejnX6q4D4X3oaseRClKt7yxn+oIroEDRgmw6FE4DZAWjqGhXECmYIyONGHf
fuW0WCPQ8ZFE0jmNcMH6ofmubOq/3Eg0HSpJ4SIUVrw+gz3MBoqSs40TYgy50zcpq/8hzl9WZWiJ
mAf48ML/aCd5Jhq7IxnCFldLIK0rWkXEb0pQ45MfXxftYR2ESTOH3+49C4FN2u1AUbIIMHYpkSwJ
8/zP8hLAyu6AQfNwwbk17mFnntYRLHJHc2PQs8PBPuC9E4/ickw5kLSEOFwoC14cjlS+hB+Ikyt9
PKtCftvGEEL54kmlhqjxxF6JS4FBjIlpKAeyiaUplkCfyuh7UL4rGvZWdA72WG6wo6ezyLbHdJx/
csGVY1db+lYbYmar3+YBYKeaF46V6lOP7D3zGg1+jCVEMLr6KcpN/U6gdIRJ28HLTcLOQRb1vXtW
p07RxerxsykApffL/ywapl64nBk1BGEsSpCjO5mQhNjvMJy8PtUM70ZN8JcF5reZE79hwRs/VP2t
2QTR4uThy2bg31vRhVTpazgUpME4ktqNsBZrst4IUvMB1dLhJ45s1rSq50Awh6qr594mRwZV1eYa
dd4UCL7Kciyqr9p2GNDiYhFwkHIVrANTYrNLENZjdKzhyxB07igo0ualZ0o4b8AvdmfNfts/ABGH
idT3TS+KmRI7sY1EsESU/57Ez16GMg84QhH5H84SWBhBY6iOxeg7PchgCPmJTcFFYiM8bhedztiA
OiVzC3eMDtmaWHdOtKlC3k7nbCWdZZJc9JOqy+vErCZMRVk7m32lnqq25p0ktVdyUgtu8InW4wJB
7mUiAH2rmZxXHn61F4YrSNbcpS1HigNJUZtR/vTR6AEfZ958/wFb2TN/nCauXj3DV7Q1NGvtbFBi
6rEF7KAZqdgP3u3O2/oWiAqQV6Z56YIEiqq/dKdNAk+eDQGZDvXwMywlWWg/QDzT07c9RvL7HMEf
uKGlQHNGy2IaO7jn1ufcwAku4QQovlKBI0kktOnNmOjyq9WzTGfzG4wK3XdUBn6M3sE2tZGPXcOy
fhiBEKDKMPdqUURCc4ysRYjAx3X0U6qPM5pHVmBxDMJBoiglzq4qjW9fydNhLs8GPe1PlFwHXC0j
mIVMtE5AhZnBeSsZXLEhTwzHiOtImbBydXiXX9Yyn8aaDQ2YgxxSpQ9jFDu4rkWy/kuE8OUnE6RH
2Mv3xji/koT+gxDYn2qe6FEGgKUn7nSynBn5R1JGOqjf1FRVBfUNKzckEHQdlN9WCS33tEAT86Cz
zd48VDWFUVW/qLoXviNfpdVkSKR8MIJtisMQsavGTmPG+3wdC/tIVppPuwQ7//5OlmPNmwwxUM5P
hDpv0+KIHDrhp8yplB7F/KU89NRPKzYAwn3a8WFapi1/kzdYXzbjRhloZNiI5Hxt7ruInirJKjN+
njijUbckzDV840BgpnOCd1fl2vC20qaEHR9WDA5TGoB6wtEBVxUOvevAB+d6cZEUnXGJjQoB19DQ
vMRN5ISZKDGAE8qTvcCFujY6JrdfazSipwobaJeZOY5Vdo2ErkNa/wumeD2dyCvCrA5Zjnalclwi
mFDWnk/BexbbJQTpLnVmdMnuBQvY5XuekUb4sdbVobmu0HEkdGVyjzhKleHM/q8PisjFDY8r78ZA
7lGZgj9Dh/d1VMIl476kdSDe2VPMXp8ffLf5O/qIwvssollE6Q88o+gEs25VmGxMcMZCA5lsjDh2
SCaqJuGO0HXEE9N4pqlGlWLjrjpMedyDAwpk3KO05Hw6puGkuRkGU65Sqec+7q7mFjfhrkyhfsNx
8Y6USFwER0DcR8d2xyjNNbOPXEfOACIJN49L3w5LogtU7vFT9v1iqlxOAeggpNr2Wah6K9yabrLl
JMnNSDA7mxD8hliMaV2Re329tfdDYWAU5xkmB9MEoZk/SBlG4tJ3vwqcegD7Y0T+aOgbI5gLKXFD
fgppKAQJnTmpsTd1n2G1L10VOJLd5QqU130p1kJNc3T549dkGEz5IvBas2MQp17OZ0FOmX2qpo4U
6NdLYYZeX02YOlMKJkUe4wDScoXqXqGfLO/dh3SjJg+YWf/QCP8BNc9y9lx1iAJPSPJt256FiuN9
RgUsml6WSh+W2myCob0gZyFRtsaPaopjS8D52CbWrr+zGy6mUJ3Tepa80/PI8BJaSf52K5y8oL/q
9sr+E1hLRkSrZOoVtkVnAv3ejJcJ3jlnrxVEA0pZcCjvGO9qjDfQIMrcnTzvcfKDsgEiJftH2RkI
8HeaeWNF2vekLDAtAu/Ho+QopfBJQaTidIRYEm6xzneyfKTi5GvHS8U2TA2prY6XzTltiT5Srl55
DaRS87jo6mp0fc4yUGLovzD1gzqgA9+rAz3hzLNR+r0H3IrXJHvbvja+Y1M7pIiLkbNJzEnheWNH
KpcDo5R6zoRv3wAKgY8aAvJAHQhmKiS5SqjCHQsKBOWTwxel5l9QRdXHdoicbgYBr/MkO5Sn+Bx6
DurB0QOmYib9zMIK7iXFqn6uZdhcMNjokThFr/w8xyoLgPV/1wm1AaYjL855RNDjr2cLwLBNdXly
l/wHdeXcsCoJqspsop1VNAwcDMXVjd0UHSNKdz/51OUuuOtPSeS+VA4RkIXPjfvLaTPbTevwVqNJ
2QTx069oREYW8H3tC68vnsfE7HGcysMaF/KHmIrnGzJSzfONlS22dqIpZZxk4VMeQUZ0GkVs3bd0
HUDxda1UlNYnDrht04U5pnigSTe9e7d564bsDI2N3Pw0plM71gRVbi7kVHmGVv+HEExiLg53Yv+l
YhQajB27vYusb5hqUyQyPF4GP+JOEm9gkbgH/8pK3vPRNkZZEFXMGyJszDiOO/D4fQ46xrAMYxdD
Vanas8yh2sZNSv/VuDfdE6+M5EId4W1Xgztnn/ywyMerY9u6uM46tUNH3lzvUa0hJiXK6mibM+nZ
evXr7GuM7vRzsCVqEpX62f/W3Scm27n4IvYaz+DDGibnJ3R2QfTQghPAcILChjNlzY920CB1DkSG
Zlo8hMDpYofHbSNyZj+hlc1SK25BskAvS1cX8lmoIzUsT2TZJe4ciXSP/bSOFo53CDOFXX1VOKva
x9mgMmoLtZM0wEd4tNlSiuqESLOQ7HkufSGF87xfOOBpjVL38EK5IK6HakkYUnBvk865NSTypl/T
UvWqw4WsYMAo/lrSJRn6DSqKx7/LiK6BicOzyeUrwd48ASbMPYiulKmxVMtFBoT3JEGzsqah5l8I
ze0Rik5mM5ktqtMjMGZVylzVzlcyWerKXC0rwTTBNgbRBXIW6ZqAUaNt23ghHbLlU7jz3Wd1+qgQ
1lLJhUKu/zNTyaoJDDKtJbyDZQAN4kIWPQCXgZ8pnT5Z5WWcJhrsBO0lE6rBftS5V7/bHFgbB+Km
DUasHJzwx8TtaAmbXzEw9rTHb+h9b68EB7J/VX3WL98cuyoDy5YY/c3ttIMG7Ua1CVGBm2a1p7nF
rOBRomLGWBXD5UnI/aTG3FzF6bbEe9WNHq8FxfeDs1IAdqMibZ8jTIbqYvoNVf2OLSH+pAKq97iW
JS9vy0/eOSWaWclNBmqIMjPOzO266WmHQnlAk5E4jf69H6x/vx3NBDgHjnm9hJ/c7ndjCETQx7xo
72b9eT0bkuR8GRbn8MjCa+rPYVTTxkqX8dc1y/okTQ9kux677msIuuOBvsZaWFJGclLf9v7zeyp3
3jwvz7BWMY/JTFY+m1IZRr/ue3LU2X8NubwDIvlYnoUC3593tMHZFA26SvpTzD9+qWagYaWNvg1H
yHKb8yK6Q58aX0kTjx09ce2Ix7Db0B2WmacBh5/k0kCiX0CEJeBiqfAqB6aBJfewVApWJZbUvJGL
TMzqs4pUrBRSng0zMVNTJ4E92sJRG/zLuc5WKTiYRV/cYzxAb8xBrmEKGErikTP7S0zcj6M2np6X
p7aJ/QuSAMUXFzQHv2GQ/roy+sfOIROlwo+imYZDqEisOYFvpnuNCSh5P0cXeyiJTZtFTRj2DIIP
qPlCGeSICmycnbBzJkGOW1RRQfwNf5LW8ugwHwdu/UozUEWl2NYT7JaOUajMRuhCy2SiHhh4tng6
ln2TFtuvYwm/Djso5Y1ToDiY+85W9xmPLNVf7HZxEUJtt9Jssk2Qq/9GWMM4LSMl3qhikM33puis
+r12o01ooXBZqMEIDw5X/33ftC5l0yXSevnKkG9bi5iLoVHaw+Dy2i6fimdWvtwvgKwhdwkwwzFB
xk+x2P9OOJ9rKH+it9j789sJNIhCTnuvbNMz/IZ5w9mimGQiPpprtCPUwPSahfx8fFHg2hI34omN
kYsuaGDRLZAOlQ+GXarTeFQrLr4MNvldqve7nUVKSSOTvITc/6h4Xj34catdgF6nY4RwlFDlNbAs
xgA0HeBgHWHWYL9qjVLtTuEtQ/QI0tx9xcpmTTDmt1mOHnMCb5UKYU2vselIIBWxB+hcwLuYYn0a
Vohe4utwRDL5KPTHZtEO9X6oBvFNKHW13b5ScDp42IGRYOWrrWEn7VJCsWyFioU6LG+1PCkMfBy7
QsHE/0OGeHwk5pWaMo5ohJ2j9VyATboDMOph6mCM88/TrRj4/ZmvlZ/CucIkdP9ZtTC8CU7C/YzN
FnpVNbFIS7RWUSqEc9tJwTwe3WD+A180Z/hcDk8PwfTCDdUYP4KwkQFKeJ95B+ZUXv4IWGxJNVc5
lA36mEmYXHZlQ2ncEANyPWeUKvUe/Y92oeTx3NJl7taFc6vAIEPnQbRI71Smtw2KRLquoijr7qjW
R/SCHCqOWy3dCo3ruA94E/YZt3Szr4gUi4fcV4aO108Vxp5Q+9P0RDRIHzX9j3LdlBUcPFK/2rO/
c5kJYgmxmX7umSGmKsQb8HXzV9qANqlZYAb0AnDCRpQY2Bw9Gbo8g66VndX2ft1O1dkcmJ/3m3Vd
VbqoBQ8NgUydxPYbVu3LtTJo0k6Z+zJine2pJNcjhFY4mcwm3i02RpuDbdchxTcXPsAcQhGhJuu0
2bV1egwteHaoBfIgFWzzFV0E66iWzF2mz7d97CjzgRk5HIRUSDddmwGtoegy5fVUzltXB5io1ZKu
drAMm6OoRnOFDgmGurrYFoTxRmbrctAUr2WC7SbAkP34atB6W9w18GuuqzbpS9Lu+sTGIXDl/qEI
ZTSPOhkmekw/MC4GMzzrPFIUllACyBU65FawlUAJMpofeKZeUXglDuq5zRjc+U5BIYnhDqLQSJxT
znrAsfn0WFuY1OF8atGnld01Egh9FtHT2jWedHDXujdGawJArC+SpWueQKMACD+MNjTUSNFpoSEo
7fG/Y2KEUUqzZio9uGB3aidf2pLZW12wnmSv+evJIrWsOC84act6nPVI5zJ7gftdRNcXWSjQiQAI
j3o48W3rXYcpA65orknFbZpFjRLhgoApd9WC23Z5Lia6ac95jnMqVGh1Nn9lDOMm4nM2YiADF/1c
zw1oHniSi7G4PGZvvhp56cDJ/Yk/vVPSlYWsz+jpdoi6X374mM83eQYkdeilIVEwZ9pu53YYQ9eT
pQTl7LArvuvi3zi8dKo0E/4mrG0DBEU/kHrE5WTYBK2w0l81AkAwjU1uPPpsd3Kz+BcxoMSiku0X
77tpydJyqage1ssqSR+V+4WanW+7MWxPlNmfapOOgQRzJiKe2af9oPriAO2DYPLsnuj9nuve2QWk
DPe2zb9EKO3FW3+ofpAzpazun6olMg+aF3GH4w3w+13e0MkMnAa2TJ2Fy3EGLs9hIExSBiuVprL3
ZJQb0GDNvFS3UI7CXJGxbu+lAZBbqzrBBSGMrLxm+XkpM/M3+lXiBExPkQM2PGb4Pp+bqlOoSrSC
Z5N7BaN5TFjghmWKUnIlOhLglaoU6r5oUhZHeQ2UKJaUfi9fb+Tjn4VywukioMn5NATt3bRl6o8C
b4qWISp752YpMvoQdHDrjyWAN6A2i55WE6x0VAZSH57eKGmGbOmrgtrDXRXYbLHNRNzSRZl4pFU0
YZi8Yf4rN9DTSS0tnv+lRc0dUFnti4aRQkRqBSzKDvpmS+Jp5SXP65zeHB7pC+EOMrg6sAfGV9Tf
NqsrkOSgnuOWpEmaqQleEsuarO3FQEsdLeSwe+qnbB6Qm8FN5Y10OGpxLA8pqUiTZEHVTxB0Y9Bh
QVgBDi2nfr134vVStKQOJxVkMNkMzebXE5Fjz4ui1ZrciBB7944I/KAGDhM+PPk+E3Fn6KXVvXjP
Xk9HKBW1gObBSgzrP3RrTkaAEmZXCa5vcn5hcsHF/Ev4tRKi75/5DQaA32tu9lqRf80Ivf8J6f2P
1KtLTCvXU7q4VQB/Gpmph2bVHaK1ePkVpRJLozdo2Ibg84JRiGKFX9sJdbBDFuyvltEeU2HtJoJW
wfnJqFDf1igtiFW9QDNB0sJlW4uFvo9/cl3vnBaseowEBZ+SyOKKlq+Ll10xfSX+d5UKjMC4XBY9
ZElrvg6l2nSUGssMo3vDcgAQyPFX2Aqv0RjkfT4nJAcbSqPZmKzoI3qurDlBaWd1sZw+NZJHmctF
9J/0C2EArbPLPhmFPyo5l9siBNtwW5kPtxSdhVaI5XtL/JdqsFOY2MpagYkmzeLcQZb/iZUtaH/w
jpU049EntqJvfDuBE3n+LJ3vCn2vxUMtmp8A8ZgjrskjNriYA4H8qS5o2EfROn4U0vKhMxEBJAwE
xChjOW0NRn8/sHJ1iHXlDig2zzlfn2nXG7ViE/WGxaBUT+QgPl1sN6aMSg/y2NxwqazU/4r+nMxW
zWsWs4VS6KU9l/0EMjUoIgDZArcWh9BWcw5dC4/SpzOwRrJTDqDEvbWWQ4wKk0JS99A6xiu83HaF
9AJZ4jg2hrjKwJICNgnL6/gHW8N9R+87pkxUJQzI1ykWpq8hEIFYlgP8Dr3bPBUZvyS1VuVYWRGH
/lj7rBGKxdgiRLqxoq9Dk1a1wr6Rn0vvW0FYnXjSDG8urvFg1vn1Sy2/81xx7yabGRq6DdDfLlcp
MoKQSFZatkzwSxdWSvN0LKZ53dee5s1OpC8UAGzDpbx35c/4dZ5rsgbFzfB0isqm4kcCn5GsboeI
wBxGbMDV+LX4wBbXnhvcdD1zfvePONKoHoJyII30a+R1u3Y0XspWtsjTxbMpeK/pgn6jGfi3oOht
IuAyz/sXc709qyPG3xtzv5vUy6ZaxAzcz0S2ABl3WXtRSvZrWE30MPgmluXhy/RKzis5CnmTXH9N
QeYO7qkQpaE2Hx38G91qXoyO8x8Ddb8Xs6JCS4g7n1LG71REeqWacCLTSTjdujlOSzkjzXY/3GO0
EUp86hDKpHFvrYbth9BLbbhA/tDSjOe3Yj2yaDCSwKGeyEfr6N/OT0ugGiacaLySb1QLSGEyTVmS
miE+MYkhDCMm0iHMHa3+cwssn8/9+kSb74pVURyZMVth7xX2Ju7faHyUlq+QjA0KYzXjJ81//QjK
h13FmbBq1xNf5UcSxbe4EjWmdMix6Sf2pSUSqx37cSU/6rPeIQJzP44WXJMuOJTO1ekjvKeR0P65
w4MCIq3rlY8YY8EFr45oITZt8tXkCMP+dCfAHeCpyDbvk7OygsfQTyJbClNNITQ0hn1gu2W3oBb0
drvysh0WyKQgNpYMhx6ydnh0YRpg4kJQ9UGFjhYdXotpv3a+UWhhAr2Ta9xozpwetLdDP5JyuIP3
3f0h+fcB/bYiT4dZb9jKgz3FpDCfujgvMIKcbPyUmQsS7IIYLJpWjewsOKv74Cu3SVf6YBA6uyXY
601DtB0Gofmu1JzsXRPhiMBT1E77sG4RzE3zJ2ZS2i6ywB/rdP/tcfGTeloytBHDkqMeDDgKJBr0
hlnKIhBnTo1RpNnH/LVB4irYFlCcsYm5qpFqLcnDP+qcfb/TMylZeugBz0ibK6DIpk7jvc6g8sR2
4bwlI+rhzoLIdY4bJ/a5xQ7bOnS/Ct6dQLtcaa8WDyu/SeWm2l6lk6nn4IOMy1gXsQ2MTCLi3eXO
1YT87Oj5IYM+4ILGQUfCu0i/c3QRfnPDKuGCOFqKK9yTcGTJ6m7OpIezvad3AtO1kS4H5G7fIwqh
WIFNQh/dsPSJQk9mECDPu6LNWJv0EsNM4Z9mGfHKo5LjvffFY3e5HGdYNde0NkYrMLZxOmh6gkzw
3hWEzODsq9gV46nEHi8gbJWQ7NpoIot2MkSEet5fSge865aBKI8u0pSe6bp6icizDnBrpQGUO+dF
FDFwVVcBu7051SbcTJwOHQToXFMmqoV5tb2KIIQZdfyF6SmahpKiNF7DkIUc/+Tql4vreZtWFywp
obGFWWdkk2RrfS6q2zRDXkh3nAoyLcUdF/71fmIuerAPFURCHxVOQMua8Om3BRI5gXNhP3culdt5
URiPLJlnJnsJ2xYkCmj1+20JgRgnJGwFS3JNQRGArq5pRxXXG5PkqIx+SrGT7yeK/xmr4fux+Oob
5wYW6dZ2NPAczf2uqL8k+zKYnE4d6SMuo/NUOz73VyhPQp5UEhTAQ8RRAOe+UDSND0me/eSuGWMu
nhai+xE1P4uGsBJmy6Mv/fbrcu7dgiE68ZQJfkGULu9zs4yIUpZAOwFooV+Rl5YkA/ulz58Qp3eQ
tqrELqDeh1anLt+g9//Y9gWnyXBldCS9Dm3uzPQe4me5HBIc8AmFA4iZxE+CIIWWIVeHiWO5LgL2
bnN618We1U38FR+RDAx7xftjVR05N0XP/6N5ZcWfUYRWldGmp/Y3anpjlZ4BPAbwQzDetEsE4n2P
7GwUTK6VBo9cQWtUxlDfnZVcXlcRT1EavGnG7dMo8mzV9Jobn97LzhhUvNCthFqZ7p4sJFRAtnAB
cvCGICN6SWMuQmVedxBjTXFkjk/OSyLiUtVkMztJH+0lYa4zZ5QlvNyq/skpA6zdor92i/7k21wA
VxQ9smV7x+UQ99/Y93R5pQnP0WGVF5QxTE5kBOQoWlu2IS1FuVqKscoN/dWHIobOAV3uoSSdCYBZ
AZJxGEDPRFsJLh25A4aTlTWTXV73+5NSlBxgQ4Q0tY3YRWR7x/z+YWyqWCJLMGNg2hJx+TwvUMdI
+/I8tQOZLl/fNbzYWmBuJaVw+eWBcJAQsxZDxU7LN2n3U2NSuQALbWOMHDkb0zPmpQ3fZFQ5/RsY
jmk+fPxOavtUU3Owj300WUYcm/Mn0mayuevlTDBKa3AaMVm6HHc7Gt6ZPsDV/O52RCFGa9zgbVa0
qdjUJTnoeug298kOnVuCLl56a3OEh+qJVM/FXBzbNr9W4M9tTm8b9ptzpbxryM1b8rzaqX/sT3Td
i0MGJOM3Pcdxdr0GOO9Qt2YRbUj6/i+FuPVNj3EZt4a71S6NUgNrHZZARtn9+GfGFlmz2aWRMeFI
L3lq4iqu/D5cOdzCN+PvJ4POc+XJO4jS1n9W/bn1SUst2egTAINLttpj58jz5+rl/YUu5vPn7Ixe
vHNRflfNGSr0lha8aBrdF8n5tZtuPbOiuCI278zo7sJ1snY19g4X5yk1plBGTJCfPhU8Y4Se6bj1
8WFrNnZWPHSE9dQxT1PVbnccmJ1vwjBTtj4T8MD1Ul/SWcngm9dDuboyvwJp8V3HcBKdJn1/VWZB
i1QPKBF+LFPbsCOMGcelZZB0BePmnSGpEHcc5PaY23EFM+WxdW0BM2vYEs0zpf1pxY/mSccd7Ycr
bS20Hx21wn2zl5krKWNDVEqINvcQRERFr9opI4BlSOHWS6iCKHL/7+uwOuFXw/hOLBkVHKaATVnK
tmS2ISH/UZw+vH0ZIom7vKo9T781AgqBgBnwU3M5xO0Q8/KB3P1HxDIVV984PkMSwciURe4nPxI/
tjUFORI5LsUynY5Y/Gjzz8x6eTDdXb0Ne1LS2BnTIa06/u+57tHhKVgL6zcYnOoFfQQygJghVfkv
4VER+ZY0W2ddpo6OY/LstE2cJ3l2Z/zFTgKJFgmVn8g4nWZ+F6N5Ci7ALAtBIOXNetcpuly0G82y
Lu0smizXiZsUegE2tdaViytJxEOrnTLKbKbYPHOvD8Obpe1pJXZ+2Fbf3dQM0pTX+dlRgSjvwtfE
L6pvjeik81X0/X6FP7T2PN3amzGN5gXNlgm6nM+Gfri1xa8mLMttUEZB+TYNbzbtiK/qbhBwVuSO
4A4KQiNfHMf+THJXFkhpqHXuyI4VLhSGSsCqZLGJCeOkWJVILM9D4QNBmuLcY9yQFWN1OJn9VW1f
RGxWyUoi3siWA/bWC2AHTuw9icCudDhFpwf8kT/R64SGr5A+p7LF157T21IlKgdYitpHT60DNr5/
b16Sv2/E7FtvbF4KyakjIb6kgnYFVOyMqTpucn2Dy0z1GOT0H60l/bTTMv6wyQIpZVuBJ1APNPTW
/V9sjm0rG4kw+0P7ZIiokYYln8T3fs3li/d8oRYYbsoe4WHHtOGWgGV95XxCaFfqhbxRSTVzM0rX
WuJeuGoaTw/LqMi0tHAdm9qaMWOZ734jQVV4/oEgaNqauMrPUxmBZoxWGD3joNn0ClOkmThrjo/q
MAd6Oicv7r8M/kJGzfcRW1aYZJ+YIhWCRgVz0NGz1MRCt/z1+kzcjFSzvlhF4ZnEt9AIQG7ct1VS
AXHCKbbhDH/BkgTB3xR9nrYGlmSez140jZD2ClK+bqMbycXL33hrb+RZkFLHz4qUwNA24rtdEcjX
Osu+eBa90+aTqTjjqxbZvh6B224y4d7doFz0k1KkKr/Wk9/OrR6+F2Vt/tRZIUs5v6eL4lgtM+5D
0rQk2denKIbQIpx/F3lOpkDi9TI2pZnmrcPRsUoUxvEBP9ZAUISL2Q5mUIvdMmYtdCfyhhHwwLD2
IUbmu7pBmmXRuUM09T3V4ZrBZz5IdXp9dksqkEZoQ0DmYew47hH2aWuZOZKI6Gqy47qHGslzuJl1
pXWxyrINEHAIRwk0sZyJ0QleUcxPP3kT9egH3p+1yAlSve8ZaIoi0uElhCgB7W/20fvin4d81lmR
Ot6jcCwi2g4de4FreO0is4O5P/e3QizObTuA0EZGRE3kE/aO9PGuI8JxDHa2xZQvwQucX3U+jfzt
HxerFa0VNegg8WzV3BV99ErGPNcVMGuwe7lGSHMQclCbeqYr4hKT6UybA/wMApRZjP1WIiwBb0R2
Ncx/3Lnii2bL/x/EOKLLDmB1BJh/9kU7/196NbalFQIAQ8QhrjSJ4l4xDgvm/zyvN760O1Wcj+pz
/QN/LgRMF7epsrq8p+oSLevG2bejUYIxtxQI/aTHNbVetDV1KaDwxU5K4rnRWrmj8xyhkksYKmmw
GbVIsjbcn+//UxUZPoYTM4+Uf+OUKRjaapPVNldiQBWZ1ChE3x3DzE1pvwQYL1X/9zrDhBHW5OV9
iJeKXoNETAC18kY25ZIksuTqEgOMuezLbLF3kMkktFKTAp79Bha9w/P7NR73Z4CPPpB8Kuf1Ok8y
WZ3cuM/cS2pzhze6qm7fYHkcOaay4pMuZcraHYayXsF42N1RprDrq4sfXCOnHoCWyDVsJSgVJ2qT
qS2c4hFIfh0pYD5QYtf6oqWj+q51gAojob8Td17HePPete8bWXj8Ulq1dQ/mzjxWwNB6Z9qKok5z
tAm55LUmYinWXktllj6LqlcC6zXvR0pkJ7ILrTMsLMkAMNHAwUqIM0vsQ2oQbyYnv9/RMGOCsUi3
q9MXvMGJsdKMSYBSdu5WxoHF3N5MlaItLipYxSFj6/u74+Xuu7e/hOmHpgcoyPlZLpAj4khABSt/
RuXV8MuZFTZccDrlpGrnJKo44G7JW/ELPg0Sisn2Bi8Brr8zsWnXEC0Hr85BoS7S0xnWQUZWPCJA
GnZQM21YUSEIIudn0Hicv5Bj+y3KWfnbK8pPN9A/zfB+6zHWiAvmtfgf6mVv9o1tlv1+zHZz42Sv
HpceHXkxMAmqExclywAuqwqmqm9CA/E02jSRKY4gVANbc7k/lNvpXNS8QmDxRvcrZ1LIy8ZaPuSl
Ku5D5/BfgbbIR+CA3TBmn53bajvlJQ4M7r94Qtv2On5GhETNZsMayORl78q4qeptDe1VNPS415gk
RKIi9ZOQK5+z5Y//pScR2nX+DxY3mULPB5xMZFkX3NukqAn4SgRGXoclwsEox4lonHtYQo5iuJca
pAymA00wNKW8JjyMpawKyn0GpUEsA0mUZHPI67my574BEC95wus1FhfKg9znSE592apZzWig8xGN
6342Q0l0AFaqK5HYzWEieM6yq8s+lo3ilOt8s4fR85y4Bdwgiv6pEsEZnvcrz8iEbVKjFHZGJGdk
H4ng6okzitH2u2lffhJSYtYh+48PZKU6Qj651pDSkrqmr8BuxplzT/TVwKL8JsbS4NgZ56kqZfYn
z2xPAwmh4xtMDejlp58ImbqMaUDeJxFOrRIKG5EVj2/ZRhP2JJe1pQSIOK7nXgmj2I75VEF4zXBc
IekmlhtgtTbS1JPHpDpvBQ2+Uf7A4AID0Ce0Guz9PDhZX5UiuF+9mT/QB9l0dDSg1SEbuweuibbU
f1XyQnYubodv3iyou4t5eR1h47Z8dFhWomztZauuZbUn1NAnqZeZ8lQ7w5r5Q+VqGwNIAWQQsPCx
NqGPBV5CKGQQPhh0g0GOTxNsKHY2yy0jdDY6/2VyPZ46Etqn4mEcSeEYfmG7E4r7Z3uebK+oUdtV
tEJ2gLL4Lx24tPk4wUfkNe9S2Hq2yXJYMviV1GvuDLunQsL6cOKqBAITnqM6IkMqBNUjiY1Do6ny
Cv+azBsrG+5K5gLxIcLwgd/7hxgj+/OyDosxRTYX8Wj5Upjw5HgoPMgOEYnfJByaI+5tskQuUcrj
bM33daz2Q/PKPxS8i9VsXUf52Sb7/IvAeiApE75aqD8vdE+sWALlaOM4gc1HaVq+jIXRA0diNpUM
ozuSSiiHHXkiK0fgKwrC6aUZH/tf3dNuWdvPoxRQ2tB0ySfPtmA5soEXWqV7rcMq26GEtAD4TDT1
cBh7ZXiHaN8BwD+rNIOy0D9nKnPqnB5tkdrH5ZMLP5fxphO1oqS60EXQNsSOYPuQLzcci2Xazqd+
yZcXwATk9BQGjVx5aGpl3FyplSQ8THuOQNXGTmOnlBUpoRsb0Te8H/aqkRWVl58RJbS9+mCRAGPT
9w4IqRuXMnqW4/bjwuAAh0G+Rqu0NT1ciie4kfA2KigCEVyYh+0oNHtP4Mv566AGZRmbtRw6/Vrf
4NNAneAXzmYMTSP3oPnI3e1eXpSGE3XL1rQ2JXxlz0E3bSngzrpz8Sp1aQwV7oDN3eE6vVOQJNzx
Ra5qHkds/IEdGv4C59wIsog3fiYfD2ASoKjlTyh6Ho39OADMqTAcIzjF2SdWp5tD/kNT3jNFm7ok
oRiq9C5JxB1mhqxFKycQALm6vygCUSllRG/Co/f+SPMF+tsQMaKYuKJkicRWBrVQWOF4TzosIEc5
3HRTBMIN86Wy/i+RttfBeRxGgZ+rgQoRKESANnSIYY6LHHOQ5O3E19i06eUHUed4jMkDmKGKm5kl
4IeS8iTi4kW1TusmET8xexT4A4m/27yqkFgZEcZgHY8dBhA+4FslAdzXwb34WDAEfuORauwjD807
ohJ6oq0mpcq6ACC5iqzHZhUVmiEbiQe1SpouVR6JjDOEEmapywpYLibkzDbGDdmFBNBYXr4tjJee
ZIQ+uOxz+TlXNRNtaDGiEpp+8DGx+0BspN3FHyWTiso7Le34M0DmS+PbRCB2SyqJOML1jiQMQqv1
Ck2OypSzxZCBGW1dBkGMr9bZ8YudILQLuQrkYI/tL5efNzVcHFzKnxBNvo6vmnL2PyCwHMpLZWQb
7rioPCPVtK+fekhA5X189uAdDfn9BEmVdDIOC+l7a9le7io6Vfn6CLJ7lFdItm0+OBdoRS0SEe73
/iV1E7rAl5OhkENn6wJlZZOIe85YxXnj4PMjzofK+wcAC+F85HAZ/i8dAVdeZ1HO9FCNNBml/WoG
c5Pqjf6aetjzGnsALwwGinNyrXe5+FoFTWTSoNUj63qhoQshkj/psg4icqowPKDfuzmz1/wLxei8
JEvKNhTYqHPR6RYDSJJp36+HR8uIEd+mqdLSOJmNVX/f7FYRRfVcjOQpSAFrVvKNJL3rRjm1P3dQ
xJcNukHfQ6Cu0ygdc8JGegs6HlVyqWsvAlvpoTJFdRJMwV+8OqQgzyxi/ogIHUOgYODYqosiJJ0M
VG6i9lYPKTe/oEdx4SJarUcy+s3wi/PE34SO+vlGMXWIUVWqh5swkEqflulitwPBRgMNNnpeZX7I
BZpmASCLUDNDwP5bg0ow/LmcdVyMzHHkYc1vt2AeyvOvJouxewkzAzJWsiurgsssGRK0yTwp4Dgs
6x97TxL4VRH7x9VDY1y+L7TMFgw/795w38IdxZG8pJmDzMuTmoIG4fz8ymgTLkPU0iDV1xqA3Lfl
0tPl3cbC3yzBkLpswGg2NjNc1JhLCghCKgYASvV8Auw2TU5Ayy390lbS78pWPMkRofyVf0NSHVkO
CnaK/oVl1Xem0XcpV0PIuxZDmr4jWf8g8viT+Ty8Z+ydcLnj5Ewzhlwg+Cxd5H/IHioEXjzb+cHr
CCtM9+wRXhu9qXH0HKlfS0Jwn0BV7ltqnfNal1RS8Tpyc330PlnVRAiYCmm15oGnge1LoU4C8Pit
l5W2Uej2hBkqLFEIR0CqUKfyOvYCVRBUvJcCMHhH3B/ugddq2fQjJ0xwnHAcSZPbtqwwBCV38Iau
xmDgYICbl0jRGg5lP0MtZHB8/eVZYrOzroQHvhVC7Oz0L5kOsNTWxniqqgJZF7HjI8dODfbhCx0N
GgPScsCNUU+y9lys9IfyUohVke4mXu42o32aXiB1gAomhV54WyIgh0auUlCx2r1oMF41v5T0xgAl
HaV8cf0lJ36v4yH8eEIHyf55j2+9I+lgFdUeWt9xwJkSW1JPrfh/mOv+8pWCuPwIMAjc8wLWmPLF
lV6w1USZblXx73z08inow0Cie04pYbI/rk8G0ftLC7GLmZJZybFmIlOaS2oQRMDOk8KIZvMy8VZO
8QZAJSszmnxfWqqZrqttC8hz2NemslOQLvoVPMiL05De5t3u0ADc0r+u4p0Cq4yD2Fys2rZ8GCNS
iBLTFsAq+BFChlORBLmv3AMGRjoqdNK3xEv8LkoFj4hUUqN3Wp2OV2af19hPOauWaiGsLVT1knys
ssk3u7+RBjz4gAxCX4a23eyjWW0LR0DbmkKqQZGAv6CWaLB2ATgHgT1nuhgLQTDymG3rKFINrzev
paSbyPlc67jRcpgvooBa+1fXZl0XTwU+LBWjnBZ6OCDAtU3dzk1yk/pE2YwoeaT10dxC2eaCgfPn
tT+wqEyUE9vLGo8frDTWe4Ibpmn9uR4Zc6vCVA68x1ZtfUG1ptz5hHVcCkne+8z/AVHwRVObwe1I
4nK+Sh65sG9NLLhp14qxqshSuFiwVkjF8ypDE6hC20/BOnhJl7rJ2e3OcP7wfaxyV5Qz6XSZ0qE6
Zq+ZFbHa29LR72/wa8EpHxW0Mp7H/b+l/XFvrPFlwZUc/+db9fjFYBHrR4GZrQYuuo6OE/M13tgJ
HOTxGmygP+7pZwFQFD1T2T39R7EpvYhY0HjXXeq1nWVqxbD5wdyD5ezObm19u9cZTmLLwoklsOrl
yH6MQvfIBNHEoDHcZsa0L3FSi17qUfWQ6jXo08Le5wpTHWApWraA4yKSwfzegRZszgim6IyZAnjk
9m1ifQ0EQmLWr7kQ6ST8COmD0MTwwoVyEx2INz2TtSyA22+6rK70a3P1+qITVjGShzEsgtaTwNJH
UErgS7hyXEd/NxC05Ohco1XyFVgRX76ek0Le6RkNa86Z6++YOxsYHBpMx+pOkFExfmthvqolFbdQ
ynO6SdwvhUcXDupu9WvrSjqDnr+VNhyhY98tI5Ls6bspsu28hEB/0mWU/n6yjoqI1fB0pjFyDj82
S0eN4sR3d6COUcsHQL8fRJ5TgSAQnwrkNDaBrjW89nugJE37NBwMg9eMVKUA+rzwqlb02EMp6Bv/
AhYJ5YpkahvurwDvmdaC0tJVkIygg8lMeGjHic59KuM0I3RXNgsEcIcl/7xFXwxAo6du+FlWaa6x
m9wK8rPeSh8CFtUzns4HN6UsLz8tMF4KgdJoM5tfL05s/jQYfs3QD+kJUn2wiR62Yu+ByG8wtWUZ
ygkZb/nlstD9I6ql8Wg9W7ZO99ehWCaAMq8n5onhWZAt/tPlodCld0HzWYK6/OXbFaFqu8cIfqTu
4t5cMgOuvqNSObOL9Irz6wr5LNL6vTcFx8jEYbmAtPJi5mmJ1YzPK5j7HpFHuw/mysA5DvSAlz1L
/p9YMlzg1S5HfMjKZ73ClsQThn9dGuc6A6/tUWnTuGsHVpuUNF7KY3++kF/c9ZRxwwzEmzHvQuNt
CYLK/PSWYpo94HtQVFrC3vQQrGe3IayUCKFVkIMUQqTFGnl1h9bwSgDdck3ADySvD5LOz7i2EFiv
6JXWsxNQYk/weJFPCyoEpVRIAgqi6MaYhdHlkIeo8bRetdOoOkPQq/yjWfivHnrhh8H9zrR92FAH
gpF/ERxMrui8DK3+r4B3Vwm1yoCGFxxLzrZ4K6QxO5V0tTEPKRl2Ki/6HxEMB3u+3Odya4bEPemr
ea30OzqEgpWsC2QOkEw02Sap9wlrLG49yVvV/8CP8zp7o95CvdwG0BFIq9Qwef3hHWSHADnE0W54
FDP1/FvVVdvccNJ4GRpqnQBRWqpckaNPNOYU3NJ+pzWMGLj/W3br5b+6cNFGkIS3hgUsQ42Dy2M/
ftwP5yIhlggY2lz5p5qtFk2y0mYnjuJcZab5+thwgyfdOnxHJdomEltMCsmFMi3rcGg8SLhljxOH
7aXZuavWXPgLhcCG4EMk5Z3OSGg6v6d9KVANPsPqf+R/eFENf89eYk0IA4dmhb0ce9gHmTNa/qO1
ih1Uf9OHcWgGdXxuIE6i40pPWa4ErrB0FrnBPp/CYPx5bbVqyqAZ4uwF7rrwerKiXgMsK6LELG7y
4MUREUhGCdvTp4XOFgyvIDPzyJDll9aggWvki4+ps2MTf7EKgIe61C/lsHFkPUSGk2XNLg9AplCr
qhcny5kOyPclZ4z24lcOWoWOxngShdgzgHGVE256/zyWMMKl9BCzBjGiaAYIQ5KddgWiH8HmlUI5
seZLnsrz5HamW7u9KHZBaTYaqZwXSoocWXK06FL5DbDGsfxrm6A/1T4IK0naMm5CSBIDIGttHMab
ECHjo58/uhHQa8dZt90s5SKrH+9JtOjKK1S/S0Llp4M/jO24g3+0WzoXFD6vvv/PjRmKla7NheU8
l+MdKDshUfUyfJgXXWWm0Ck3pAKDNw81n9/x+7mCsmWsxfKINAhCHXjtCjbIuJvoZQdzvETtEMlH
ei9L0lXx/sC+M+jufsvbjCbHz++WHc7ywulcz+PzKHSIxMIb9KmFtSKfHSq+icr7qoKKVf4kI6tT
LDRUl1bj/mIGO4hhFzyuyJF2BWpasxUuvp/NnyBdWi8GOZrTqBqfqBN8DlnhV+h/fDwg74FGtELz
YW7XmWCjXbjzL2pvdwVfvk0Y0rPLRdF5BaDQ2oOKQby3UYu8BV9aW0et/UiCx/t1yu6pX+5MP2fJ
iTJyv87vo1UXypaGZ9Kxerdjtjdi8sN4SW4dL/vBDfzQ+nVx6LvsqZyjXqsKk6bxazfmUF2carsQ
w/eLUQfQqtzsL/7xQAl0PqIAkxlVWlIKTZO87in3lHAPNAxWEcMcBqh4dQpojtoQ/6mkSP+Pz0LW
gYETWLKBINvB5W7aY44c9CqmZJ8b6ZhK4q0jgZRTGeIo82K7U9uB2EvW+bWURW3fuCW/iHMk8viu
h0188sqAPgINm2Sx0o9OewnLg1aGkHV3ZvYaHsLWqmfyEzXQ7UqhEG8RHFgcLFGBgvrbRA/vgAXl
XBpTFZ6LQlPowDWBd1zXfKk8zMn/Dp5W2bq4k/ioRUQjbeKx8neUtViPiQGLAjJsVmYgB2H7nCJN
i92JLLseJ0TCRog0vU/7j4S8lmpyMBt7P4IJTdi8mSCypA5ymvxyccRJyRMyRRroGPd/AwQzPSri
2Nd9VQKc7lC94e3LCJ/yCoxPcQo3ByfnjojzGstgpmSPAalxs6+5xUDLYDT7PJgk+FQRN47vXf5r
ErBXBt0utQsbzXuZq/xeWxwWYC2padquEVl0T3WkE9g3GTW2gXP4b8PDVW8b3iGhFgW4S1l9Wpa+
QYnQczY7RBs0KXunX9F0wScDfsKi+SN30zoPVBHft2iv+FRx6mQ1jrMcGgJN46gt+ghRF8LLz0FL
bLYbJNt6c2JdzNkGZ9uBq/83iu54li3OrypOv7y5aTQ+OzwQiltcEI882pr4pXiJ5Ch4kh7py6p3
u6eYKtVZP+STzTTqTf7wns/sC9X+q3Nt6PTCF2XplQG2EqvMndA4nFTFwO+63RPZ4FG2Zis44S4w
PlJCV6l9o9LX06aGg0TicahvXhV5TA8xpnDf1C1vttXjEFIIQOCNipbl6Dqjzl0Px1cgrqUjqGpT
bupiwH4yNI3KlIWMTVPpPej5cjM3Sl1n0xaN/aFnUi1QRe6pDFbPvLcjXwJiQKL8Fecpl9mERsXN
/mIWn7ktwukudRjojPQbSl5P7UrvdzbLICIUopWmGpkViRqupVpdpYDq6LoNrtNQzdGO8AC3NefV
w1BmNw4xZxrTKkp4dD0tWPGGjTN2ccMI5iSOJ4Et8dkvSxCWlWGY1ShmfZGSeI3Gv4Ho7Ud+tjq9
HVs6qxPy27RLkuhbLvvOypX/p+8jqHYUyHIttHF1kyosYIrTnsTfItjPtibYWPt7nLLvXImcg+xL
1lMZEGS8HMeCRL3huNprlXzVrWYPnaYACxdIKU3l1cbGzW4fq8M0K1hqzdJolr2Akk/7RTdIGbb0
Ow/5LEu4BlSZHBV3n+usyT54GC7cKfVwQpVnFbTsaCX4Xaq7zmS/oY5oAGIVkmdVAR35VwBe4is9
zAOS8UxC78p2EwZj3HNNELwTV1bSRtT0t87T/yKsGkHHtWotUHvxwbwg2iLGOvOeYiUevMPiMPyr
/nwaYT2/bY2kUEphlMT8o8aZihc3+npMoeivaX4xIoVsxhe6g/5AMrsnj7JD5HCR/huxho6EWqRb
oAVaVLLC38skNixpkitKHokYJlSpXX0Nm10mQszaq92eQmljOjSgV9iS/DGDXzqv+wwtJh6tkUiI
UT9+nqt6GaQhe7HPvOLoyAUCF4h1F7ewZ2J4oWaBTdVItAyL/lb6w/P0+H7r0BvtUE4GdnhSa0yQ
A5aS34IozNlGJCesDx1lk58yDkKnoO0Jlz9BoWqz59m9NMlQ5BqAgefBW0Fb9JbBZMtPuJLmpfqJ
4H0AbJhtgje4wIDJtmf2ERkVSm+S0ZqIIyqMWlJyB2VX4OVefJjtkeCf8I5KEZ46xq0BdmLsnE+v
YLNRfZSMcWgFVhm66e8z1uFBf9DLYdz0dugB1lYvFYsGv4OcumeG3zeqLG7OPU+4z6bUYq3V5aHS
vly7D7pUe2luTU4Rz2cxu+lFOxTPYLvYPeQ20NjswA7v8oWfDW/Dusfa/Z1ACBXNf/6XxEB9OQZB
khbzq6/jMh4w7CknFGP7MweC//J+oH1BKGU1C9Z4EG/TYGCL6enIuRMEpBlk6imTv+8Ae8C+6L0a
WsnkQD/SoZHdXEusvgqRADQJz6nOJSgJa1UhON6sFbZvNPadyUmCE94427OEIrTmpa6zfThwBDTv
h1VVCXsawlyTQ1hMsMWv0J8uDH+itEz/GJrKWcj86mNnV9Kw+z9Hdbklwt9MjJFN1e3n0kOrIG32
kJZYvR8TNShYHHwWTp1B+fbx6Fg69Z6PP0F2+9oxiMI3oRf5GmZY/5kGeX3FOjz3P3oxNR5P18+C
ACMCALCgFcvYK76tPCeqn7qCPkCHsdiYALmAt8+mSaCwXmHoOzilWhemjkJPwPXb4/x2NYmQEtJs
FENczRJqc53FqfLyteZWh9ZJBepaZe2l3z/I6w6q+iydNhWh6kEL1RfGrzOvBDxQSP06jsoQ+Yfr
v1ccIH+a/nel6+XZyFyfUWfI52Rcnmu9RWzEnbH/4ggcm6Pn2ija5ro1ORc8XUsxdci2RrZu1LTg
dCbNMorjyumBVLvETe/Gx+5rFBffSE78RWqvVvKDgIBFwID9JxxqYj3+2IqmoQSRwCsXruZb9Lre
T39WwJnw/WQuj+n5a04kxR9Jh9IdW2eOZCh6OnXVkRhz36oqeWosc49ExCE4OILQv3wrti8gKB1/
N+s/rNBbXxxzMe8R8MdhP9FYPHVE/i8tsn7BWRs8/WvXCxbGVTPjB0noDvkILmyKFY6f71S30uoC
EoX1D8EBra4jTxRb903pA81SjUN4HQymBU+ux3PBWyL8d4r+h2S7K5s8l7AvuNpmKajd+JednBOv
PAm2+exy8YbIYv+SDym1linzK79/VdfKN0ZBQjjQM7k2pODKeQuTvL+Iq86WE4pt0+GuwpYuR6Go
ZOoUmzd0lI3MSOC9cPvkArzeeninNhGLSGTashJP5xlHsRckOV2IDZIIIR6UjauWMft9hcFQndDv
UCjsqT58hS8RBynKXiksYhQS5CubRaTewLwaQTgNcuwnxuskuxn7NJZuhxBWeS/tg25t1HHSoi/p
ZrwFFIltGF8ti48dFfzs4Ysv5dCWzCVZkQGsu2dXi9SnxVF52XtwnAfc2MWCmI1U/eir3rsgBeoW
Ilp9tu6mGOfrq4eFxal8CGgRB2ZDn+eV3ri8q2q77Lx6V8E59loLIt3rIgOUV3AcPIGJNA02+uKG
n6rmPTK6Tke2wXWFahOEIjbIUr0PtKVCcYQA4noyVPZ+jTRyR/r/qLUvsF5KEEOD2tqMyV9GAV95
5EtbGbQV70drzLUXy0X0V4jbF9CO/QBw7FX+ailQ3m8f5Llz5O472hJuKc9bBijuohrdyzNB1VIz
ymfNFVjFMWhEzwVqSoGQjtRRe/IrCysFmKqdy1FCFnrdwNtqgNctL1v8CxX7SRGu1IRdlE/2Qgoq
tynsjwbwSsnLHaRlvdEtnS8u4SlRmmWS3b/bCgX8ZLnr39zJEwteihmElTARyK+vpwgDZPliWGVZ
Ln3YRX6UstszQeXSt2eLzPVyemxM8nVitngEzpETIY27Be580kq3+oTyDY9JhscY+JLx6buybhj2
uhUWSmEqHi+BVMUg/nMRc3fbNyNrU7NPtrVf3+C3aCN2FH6GP5WISC+qALin5bg57zgmTTHd5Qve
536gmD+ZIeWqfVglHUFC2HHP8f0PVnUSPyfSV7kknvPDXSB48FySHqlMCINk1xXE6MG6OnmTya0F
Ah2XGs5PN3w4pxIlqvosuV4o6w0L8wEfuLkWV646ieWTYQxDzlat100wwoxDM6Ai+ckY55kPj2Gn
ll1PYEC+eLto8OFnmfRHpQly6ScHnDCGZlzvJDSwSYRQ/JfXEBP9EnY41uEHlWLvczo1D5WHw7Za
QT73viOfsu4vfHwj2SDjPVDng3PuCi239lC7+EG/zL6HvKzbqCSbOJyQelLhfRB8YO4JZQaUyMQf
TsogNwMAvrd13bZ4sruN0LUjvzilysuQaY6Fc9prTFOs54zNaI1R+7GaadJYfYDPcMfHWKcQknlf
/AlKq589Qg72QRKRO17Jh6IhubkWZS8W0UTttkbN/x+huSC3pxUCiN6H4lqxpZxbhnQzT/4lQXjs
wRkW4D2chCh99TkP6vA9Xe3z2cGOY3uPixLGSSvSdgeBMXAUYy6D65RkeLkbgDyv8yNmObA4+sPf
o7Sm6bjIUgc6t9yPyrvv0wkKMD0qqV+KKL+4SjTA2RpGtuYJIBu5iDbBs6Vn/iI6ze/D0yRd3wj2
Dhf/YiodBGR7LYArIRe7PqlDozrH0eQWNZq0tbaYdJy3FfDON/nd//oEzE5EBSwi/YOq+ggl3Dgp
KiZ6mV4yj3PWrW+Kf17Kxi/gEkotnVJ9AAln6K+jkY2ahcEBi/edqOxrWWuJ8JhaJeXVhJf2U85b
t49WpuWnNyqwioRKjqCvgLPyN+91zaBauEHF/iRYKIa0+t2KO1olvCoSPLVCAcUjOdQEQmgMeE37
PhJMlEBYRRiGY5oZyukVNe7f+5tgj0HKPuqRrlt2FpUmjbWP1rN1+7j9OJ65QRTTeWjHxe10a2NJ
W6o9+W3E2wfKubRZ9V3rEYQkAPxRX7keIJGsZgiEu84bBJZo2pCLuEBD9XLVbgvfATKAREswUCv2
QAaijy+icq/l6+Xlyip8ZGpdw56ilWLPMglnjFrSJZ2DhpOJyP/7Nfllsp3EbtUYulJQxUEJ3FnY
CNzlw8wPt2kqcqb2VRcVJ39P2hWtA7kyARCUmA1KcE+1lkxzKU7ZFPlIVsVEau+JthzkfSTnqgcE
+2ZVEZj9L2EzLI5Xe/kdYfkOiOYJ1fSXzXi1TmZovVKz2hS1Hd4//Nigv1+1S4sOj4x6tEHa6od4
QHBmPh4ZF+YNtl8EaXC/P3zY5A+pj+GIW/nfSxoDs6JNTigw+BqSY3qQwEDTkNqOM4J2uDgFKQQl
m6uw9hVpv2CGi3ykmYoO/vNK1ewfl8Kos84PWsi6R6dnwVca+7FImuU967qAWQe8vzkgw9dYxwoo
tbwkumNyMY+bUxPEhj70Yd2rLgc7aJDj6j5jXrch6MGB8KKeQzBomB0S4iCULr+LhYeE0BcvHl7Z
HeYnPcUjd6P8ju9DH3dO8i1MIHurFEl6GGxCDuqS91/zVg1GZNoq0iuPDkX74fRlttK27RC8PnxQ
uyZAnqeGRuGi/nFxPvsCuRvtsN1pJaZfO9Uh0JiGf2T4vrYH+KqhGTiTKPp8nivel7NMhglhojW3
ONmRBd3ioDyGRb+BRuWwHH1lzjI+SDBJNg5Y6YRe7Rmfa4EMEYkMmacRrhtD6vb5wF3rcxxcYNrk
SbTw7jFaC0bYyjtA9p3UX1V+NlzESIFwfWdD+k45JNfUll5BzwR6D8HWlV9oy0jGWJsQTD6icdKE
2ab40obt/uuljflgzufKGDu93qV/McZjCyQVn5z88W7niBij/R4oEKMqjrevltrUphOr1g2LDfAX
iX/upfFO+QNfVLAun0wsiC/CoGMP07ysFLJIIT5rbZ0op06LgV79kn84OzDMJxD2XcCJSNBtkfTj
Xo3E6PH4ias4esscJkVV9Cg940VNtUQecuc/yP0xZynacQG7JoPXzh0Ras2w6RlpMGssUPN5SbNV
FqILSLQh4H0x5fR4xX4YzZDnP7bMf5w675GzZovf0uhoRp1rfh7F3KMnbtRK2xWhGLTGIj5WATBo
J0L01I+9ndl3qLVUfH5l44DH23VOSFOtkU4YbCDJAgwq72KXQahuEC/TfUSlh8/kWIuwnU9jkw3o
B5Mc8FGnUqUsPiECPqp+2CYlywCVpbS0MB7YtLP3seomx7WGSo4ZoR2Xje0SeBrGnhAXZUV7+5EU
jGrAbVsV5QwLVf5DMUXqktBzmh1z8R+PL8XNZZtd2EF6f5EbaHugRe4TtmM0osBLishFMtTIBD0c
DNvU5gcqZuiaOtX41BakMPVrisiePXqFtV9BOtLDS6wCPoA/Kpot28z4tca7w+nktZHplQ6ai1co
HwAl7yUZlli+GL1pMdJyBmZ7eTrE41XYmjb2FqFzbPMwROUpQHcEFOEh4BDLF0p+/bSm4Z5m7hVA
I/MIWKwSpCxh+RDeHUezzL+PcOp6dWLHmUK5ms/Bixs4fvjU0DzJQRnnjkCw3hVoDbjiNzoijv23
XFyfeSJgv0mjvCjLSfMIbQ2S1KICJQ0f6KwJkTM+fK3KvWyRmadgxFT9ux7/yEurLjEtUiDyEi1k
CbKBZGyGk8tjYCq6hT3vnr5T3lgtsqbU7FZYJjQGIL1ymTdUDcgeMZzQu/EhVr2IIraEOsY8Cavr
YHjxqtu3I6c5xl9WQRMqWDt3L8LnOmKhIS4h6+DpRjm4M6MkRUUWq5vJuQ2KUGyVVGKonZ8tFdWv
39lxWojNc5PBQTr21Q3GOepK5wNt+W4H2Q4Pl4jjUMBIstvKjL9vzYjeR0cg3+xaIffcy8uWzjxt
7erGgqlQYk5dI2wC/3wIxe/JFRkxZysyPXoCHkIkvR/R3xkUrUbB6Da5xzSjS54oj5YzO12EjPdO
sXYforWMNl40WGb+udLCqGKLyJv6ZdRXEIttVhfDFn7dJs+nUhikFuAuIeCkvgCWaTAhVUWbg7kg
b4k23Jr5vZW12Hh1XTmQ8u42Q5M0MUmlpMsWY1KinOeI37ANGe2iiRU+8sycs6ly/O62Fh0oiWeM
Zfvl6THXGqefFwSzirznjU5PxfsAf+o9epfaIctHctRn39efnGYKALBZaRM77u/3GF3bO76YX19D
4oOalUxdxBPd7MwJBdX3EMY99Lzeqx8Ssn8y6QE44O4xN5gWj+E3yQQasOrCL/31l0BLo/8t3th0
TV272W9SAVa+k4jsm2SvspR+0UFOCuPGO29Y982klMhZgcx6kPY0B2X/EFWncH99D1bShiCHBfpM
KRxbnaSHFIKRDAV+HBcV5O4vVtjcgwx08hU3kIHWyJxqDXL7QnU3QzrBT/LJCJHcaMuVVuK4c8yN
wkqygi6mHsU/IjQDrb1SoUeJFOD6NtrewvHGNL3Ztc73SB4gR8J4P7BCTlyEpcaYK7t0UbsaRcqy
RR0x/EWyCJkgiKvgXNkYiD/rFxvilxwYCcdLxtiJSEkAHbQp9boshHRBazqMcmVY5mUeNIlFcXT9
cigEXbYl0zOrHgkUOWJ4EOQfPfX7ZQgaUFcLDWUH5tb+fDWFlG+KTN36JU0fy+b/quzdmX91tMZW
bhJn7HPBt4xvdN8qgQbkQS3FiU23ZNwzoOYH6WM7fj02yFKXKwDtKPnV7niZP8Z6CwSXX3DPXsrx
Dz4nzSs+QJbgsYcJnqbB6MetSyysOtvwV7PES2c0BYAOHa/GgVoOC4rEmTk0b21DFv40Z+EE6YVO
iZ6rARBd3GsUhU5+wB6u0t4l75uVFHWBi0d7IyjSGLx3FFVY7UyVe+5SZGQWYRH4DEYl+FDuXVB3
y20MaWuxNTA1ltseyUVJW5x/qdhXU2Figj2NBle5b7oZ+Fra5lZwIWSmYCa9atuVTFjBiPYUJPkL
MF6sXlpGrG9TXHvhWWcCw6wMVzA8ZAVN4am4eUQdIqCWjWr4EuwqQGrycRiTHixw0XeXp78eTTsG
D6ujSLhazceCY516kJZBENWRoT1vZcwt5d8QdEc2fKQ/fMqiBpbqvPsqBMl2oasq7XIZ+CxYMgG6
02sCubFG2pvgn3LHq2C2l3HRohpTMigDaMYplb6RZyj/I1zgN2DmjYF6rRNu+ghnUnhERvgIcGRn
3pDk0UOT4XEwicnqbBM2XOWVEn7k5GiCtOknWoi1Zg82kEE9Ui4pVmS/botrJ9cpnMlu+JlT2kw0
++9yxdvm2UyN/vK9wbGaluzdfVDcv6ZvwqfALD3YZ+aLfDNAKuAm1xH5naoLRONu6+5rbHtmDg7h
Dzt+KsxTcvvxdcTfqZHAsqERs+iwk+7aIL9NBOvh2hSZFkiqD11Mvlrg9K/OkTNsmcB3+Y9KuUqI
E6TgGzTaAdHSzwDKmlmNFh7iBFAt+9Bzj7iAMGLDIp1nODPfKJ5r//oiCm7Undemt1Bf/3271w5p
CSO1skglB5o8KoXxGNwGVQsMU3qyauWLFYbqVtrEvIXSDpFGwLT3w9npzpKl1tCW5mFLuOr0vt/k
ZEb6E63ucnbQIcRVZs8AtTSMcCqdoPiTwTZmh6uKABVoDDK1rbe6wrHQUE+/jeQiPyGiHzU2prob
bk3fzR7mt3DRwYYnuy9Uo5uhbjVDfVhVputHvTOCPMwP79eVLpPavmdzQh6Qmbbo1F3EeU/SjIw4
EZXtWtSmGgFo2B1DHI+Begb8Iy6cuiiMv+PcYJP729nqzBAfbwfGdedggrRyElQAbxcGMJlE/134
SYPS3h5x6WD1jEpUc4Y0Dx1VxmfpAl6Z3dker8C/MYD75Sudwdaywl9inhvKvGTw4s2Bc+dGdKe/
fzrW0L9z8Wov5DINYyeouzVn6HFN646bN7Hu8ul4Q5gWO5EY+vD+adNgJEoKKLfb9xeesvNZIp1K
y+NDFb43r36UiYAg8H8+mNPGcW3uhY7gMClqyzZH8rJTnYNxDaZBlkLmNvh+fYKGNagStnVy1UAP
tThMjxnYHj5i2bNZ3SuTzwOfwdwKfGQX6dmMWUEvsnKlkNaZTEO/W+X41Y0fEjAbyVpBJjqEbA1W
ukrb1pHyWK6VeXNgcjuUoB9f0QxIWS75kWj6CuogPJ/ROKgp+ymiJWnPWo5NLxsc0tgnR5QQKPBD
beIjagrq5SfosK8T2/FmgoujoA9xn7O4Tt5BIvKblVnKDcyO4/+D/qNjCkhXuVjKPn2ZIJqsEReV
aMEkUuUPVQ3lfa1T7z7gLJ5oX7dFc9hSWi8I5Rruyq/4ehqXmL36kRY6lvQH5q7ICq1zExirb0hg
dfpILOX6OiyZTdk6YKX2hPUAufA82xtd9ZuvnMAX/O8vj9FV1rgiMdcq33BytTlkmXbzpg1Z13lz
gRxPR72L/1TOnwtnPqbJ/8RVPj6nO9zI5ipiUAWmWnXjIi4kTohsoDfoqAOF6+gzj2E2UKNvgcCp
elXKoBTeWQxhuv3XOOd0Hs+DcoDv+kQ9sbm1VfQ/ZaCOX7I2Xj0hSwmG/LNhBsGd40Tw/oNQntTH
SFtOHN52ZSccZphexAE311cc8ykMMbdDQL9FZOBmcjgFArxQENl/KsD3ymEyNKbKvDxcP7J4zMmB
Yinn9uTIMvgbwilhF8U6bbS2xFRPB933eljK24ZTVQ4zYF1TPDRugj08l0X9Wtrc2QqyNNKTv1XT
Tv9vhdCMrGxOv3n9IQjtL6fRVRZLHgvGe8UsrtBhAWgKCppohlRJMFD6MUeoN5k2PbRnYkYLal5L
xyjCASObLNPehw8/Xifvetef2NEDHiqfICBrhuDqLmsfLjQlADszttq92+1+6J4QMR08u3AXkCh8
qxXreG6pw2PTw2qZsuB+FZ1cvdEX21LDn3dbIziqCBqqKl2yj4ZWAJQQPqQf1RxWad/1N/u8I0x+
UmTYkXHylsa1KAOp0wiIKMz92yGx7yMwlXwtElzR1Mp5lsbJ8qQXFh7p56VvNhBM0w5U+cfiu0Gb
0gRsKDXvvWscn3hZWe5lgs47pkr+/j5nQCNKENs9HyzAe+KywqC3/YSRT+WDo4bInoTqAtJMJJMt
SmnUB62s65KPhnI5+OC6FFWYxSPpNghK/UfR+SxW3rQaCbrEfqkUB6ft1ywLJtISDzXR7jCrTbXJ
wBn8LmleQmq11ALhT5mjUIaU6gHbiF1MF/by7LhU8JyMHiZlrRoVRt7+X7c0NUe8Ugvh+11dH0UP
dVs20jbnZi/NBDoqoORQto6f6GeYop0nmYiqhdkVkDP7fRfvVKXiXvo4XSBJIABXpxN7H4I5TjC9
4X9vVMy7pzj4tHoD+jD4X0tSC4e9rZ0VUTGNEKhSqcOMzNQd/UcoR4jkGfM2yOqy242BfvSDX0D9
NDmXW6WtT+Ou2aQH5E9Q38+TqlHKXiJnyO2pCVwe8lTHGDqNVIt5mS6PiFOM4E98BPsq/nAceLNS
f/7urlUWQeO7W7Zr3J18OgZtrg6qxCbbHQxkWqvQ2knbiDklacsW2PsF2tbSMrev9oSDsKc7mhml
6deYNjpOF8SvFnUaIWOzNl7mmPsBdXfdTIWt4c7mfUD7++ZWWjJkWh/Wk2Fh5gc3v012AuZeHs/R
nzTrpMUy5GiNrze1pTgAahVO+nxb68Cckvo+p/dmkk51FVqDaczkue8EyovvOJR/PKL2RmV2oqxv
a2/ykVYuGOsDwN5niXug1vw6HtWMyOfrk6zfH1JSqrSvTqsZTBP/fa18fHrqNtm37DuOTC3w4Xsb
yQtJhkHXzQeV3emM4GLBAzUnCRtrEXwVviGyNoD0GlLlkdnidCDRTY+P7b0wmSZLGuUfi7t02S2B
8GWNIxdryKPlkYb5pmE55CMoVgBIzPTQb+bUaN9qrs1BvesPxe7OnL7PMM26OKCaoFQ57cVmKv6O
zCF8G/IBaX0Uu+TlSMTlU2bcUSR+4SaMWv5ZnyqW1zHrEZkaSZ0VIS+tMY9r9IOEmKKbXKtnA1Jx
+IfifkQH24Vu/zX3OkY9SubMSBksSk0kiJTsYyuwMfrE/EbTzsyqLrZ/D41buuv3hh2873Vc2ILe
jMNSkvPd+Z2iRH1wh9mBNYDvrjoDburRi7lvoslr02qeVKFe3zckxtcoI2+MStUdnTyg0vWJMb+C
nQR1NX5mAbncli9caMIUVcnCd01J7XdWSpKjui3GJZ2A6U4+CtRxOTCvdZ843mfBQ/9qmy1Xvbvg
r2FpYFGh7rIzYtn8gOsEtJJI3xsov1h3ecwp7EBdm2bUQDh0ow78wFUY0SjaU0DZjQsQa1cKDc62
tnSN65WiAdBmpoRYZimd60FrV8vbYi5nVSWrwb6DUgXluHh4+AGnW/lIIze3FA/2xkYisW0T92ph
8GmalrD2PRkIPY0SdahYi81BzZH+VpQQmb4857pHkOODmPfOGbs+UkNV5DIDh79AXFjQac4ZBE+w
6CC/l3/S7kFTdOh+MQ6ZSIzxeP6U2JX3aFt3pYqThd1XY5GVk28QA/XMQ+T07mY4eIdvjcoX9cOi
xRWqVCpZWPcmOmzVdznpxaJAZGSUHop5gh01Z8MdQCYXwRTEm51QK0mQwMnGSQUEc+7vL3yQ5cDc
HGWFQhk7A/snTXJWrGaOnX3p6v4e/AXA7huV26WbsNUbdHQi8q7eikjlafqR2h72PevBT+PJG6RI
buTbd+yDTyCkAiYojgkYpilzOzMfwVBsHHECnuRGWcsTLapYYRMPMZ+H80mdmawCLHTuJ7vbuin4
hlkatW4XpdekgLCNpsulbSF7/7Txab/icrmxVALONWWGBBwRTGrRClQ+6RNL1O2qZafVsvralrvw
obwGcOsddJC7EyIoiKPEgV/FTibClE4i8U7L9/YOoBuNPsA5e5eFU8lcSp0ONvYxY1nBwgHc+UbN
yK2FBxr7epJqs4jPjxIizqw3ZXy/X/1ZxJBOVUXjYTJ2+MiEtZ4y2awKyrNXU6CS0VMDYTSvSuWH
ycS6jkYcNev6fYc8sd+6A13McykItFbKFH5nKQC1E08sTIxpVYXPicPQK88Ci7gApJLGI7d8TJ/9
P8tPnwq/1n4Kvc0+amcJztVSmu9pCP5ysxHS6mVLr83j2JdnYE3YnwmXSxSDu/DPIAmPMs1nbYzs
xqvjSdEpkxoq7Vbu1k3QH3eukQU79H6RXU9xBcF+bTuG9O3v7OedGGAeOWL2m3l6v7ne5qTUwHH3
c+o4LinSi2yoZVXADbKN0vkrqxTP38Wvfuev2s3vMpuIdEmhzRAFBQty3AiLrhtQ0SHlBH8cx2KY
tlaIe3FNT2vwneZTN/a5CMnLZxgoRP6QhG/EM7H5MPBGGpRd1v9cmushBDvEb7Qy97DhgsIOLLf0
JiVRcu3UrJxynoiuGhIKq1b5nXBFjhsKnHNZhP0RwTvZwYUn1vDvOue/fBHg2ha+QWh4cGkggR2X
xj5h39Yn8IUqgDNSwuDxWdpb7zHUcf2vrh3N70HVYloWqACqqEuaBNTtBkpOsZ7nn5pJPpiqRbrs
z/29Uve0DXsMfIIsKpCQhmtR76f1PmGEPxFKwcqobMdoOH3uAG8WIYCOrK8rKGQcO7JqPe8rvE40
87BtXq1zrK+TrvM0F6MWtJTJul2BmZw+isJdwMOqTr7f5B5HvSogwvbFx5Z4XkupQ21sRyaZ+4Gd
QgFoGJWG3vtoOlY0Ntq12UnP+YaohpJrUISeTxPQlBQxqiKqNGGZdJVXAb9wrnOX5avz8631Xo61
3v0hXSWj4RPamWv3zJrWEmBfBKFmjO0LlaL9mAgDzwi7rlnk/hkVkwZjefrGY3fkp0qQqeY+dD1w
wtcv0+GIe0F7eoozsrWd8yBeIPqPUvw6iJpJj3b/B5yqSzUlpcxDrWNA2VuTFg4ZmbPrC00hT6AK
VMYsZyGm8k+E3Bap8iHnXuzD6jKivMco+HZl51FXjngxjft4S3B0Db2RN09tea2t30XcyH/tF9U/
Qf19CXrf7AIzrXvXKT3VEh5KzUQ3gAE8JjKEn9J2ZE7EtRxltcUmVwkQM6550mPrcQLlym/FjpNS
bzPSLwx6jnM6MTenjT0gzVJ8UWdba4CHMniCRPZxeq3HgaXP7fVHBQR4mNS2G97+tKyKXV+PnKO6
jjqyzU1n0Lo6iLtxG8vAgMVwxAZ/07tZB+Yd7WhqVuTCGsoA8vDPhAgpbAkfmY4FSA7dA1S8gGPh
lCcHk/gujGpJZOj3kqZKXqux+Io6mGhMCuZaDl8oIbzJpsXjqfYg9gSz4fg/dPF1+6MPgT3ByiWX
CWIIWszhRDD6tBNy6YpnEGkXsGKGCkWrxgxql2hAwEJ1QtKInC9rFiz9Qf6QTCp3mTmbIQceRedc
IQyG6/sCjOzjjRlJF2LSFuIVHhaYMnFAi3H3t/JY9KEOby5QJ3Uv/PbCx/JdIr+imYEoRsGYP3Wi
F4oMpwuxsY8+0m0boFhEMimlfTmP11P2o4tJOln9cxUtJ1Z4LEanF6hvP/UA8NhDr+cGByEWNRaS
JsRAmS1DJiDSJcf6DwmLMhhSG3uvt9jmcIYe715CSt7jta95229b/phUQrg89zDnTEMAbx4fR6F/
0ScJurPFjvU72wzUWbhoNUyubtt2Rc0zMiQAiMJjLX8oTdpKyRZuL+KJwT0HISYInbO/bwuEyAXX
fC9et86MHUC6BMBBcHCavfLNu1KzTxyee+Q8dnjCDBgjhYBJqcc+51nQzfvLZGXz+EBVS4oSBRqM
o5qQeHgXAsloC+pPPav1yvu+zUn+AhqZ4n4pyAkGul92t1q4m9RGK5pZUSv8qlDWbCzGA/mNg2EC
FzW2JAw/Dsy+lEWHRsio7V+36/nr4whvTVYdRzKL2Iu9yOkbaopYLwewIMmXD/ucChK7Lb9r+/2C
sq29UN/+wmo6Ag3IXHHki4fhAfdaStbyD5qmEFjhvYsDiCd6aJpptjF+5mGri0WF9UIhY8zVEJDe
CcrjDS/DDVDlOReORRZVH2KtfP3Bk7EyDso1XCKyAffcbKKl4RgPBXDrTfb4x1r5ffWpT71UM7/f
4MFHsuAa/+TJBQMglKDjH2/XnALoA9EzyPd5Pc1aQffLM91RAmtzqyKDx0BBW4hDftrI3Gz6mv4k
/6r1Oe+71I9QJ0YKXa6RmLUt65c7mcQ08TyE/HvaF+BFP49I42VJhgPfTe4S7ncdnYOlKh6W6Xf8
yU83DBlouaDp2DBuEKaD6r8Tn0SVMc4008TWSPSrBl1c0AKX+GwnK9TfFc84amK6+K3OKiZjiRFc
rygeZRf3KOggmsU2WaC5TC8sq2iSs1G3bHcyxrR6hGJvmxG2ni2SJqQJ0M2zZLZ8IfkHS1vH5SM7
/GFqqYRTdcPeqP+dc5fezwNyN08hStdzKk1/bD2qnnKfKtKt02nFNzHTg3GHOj/3IdsxrynwOLdF
iAKi++bx05G0HpPS3wN7ERNVp0UEovLMTDwS0Ctf6siSUD4yZyZBaCDz7T2LCNgxXrzZ5BP4+Ekj
C9EzkbT65SeHZ1oIJERjeheCeS8XCGjMwD+WTsUdxtYi8md648C/+URfYuJac0RFkJrYWBWv9+z6
zy1UqDoOapECX5VDpTojfUBK/fkchyV3K8KgBJKAyCcvtpZPLeBIN15J2ZbJO5ghXaSpQZo5gJCR
C4EPXXQ50XzH+9qp33HFNTLPaBQKtv292ejowEQ188fec22AA/iQDRNwjOvCnCUDPgWpah1EdvoK
5HrG1I6yrBKqvz3ZO8MUyX3WcklG5aGY/NMwCZHO1Qu2k3aSsfYU2Z5iHGYP/5oRDeWbtIiuyCmI
7/GBiPZhydVU0lFAnfa6h0QmyvxCcSZEbtL6YLoZY/AZyGFv6Kws+4xHjuqd9f+Osx8HVdcI2vw9
sw1/JZagKEHmAau3gFKvDaJmKMhLc2f2E+99uCLfIHmGuGpmmgsX48hgWJij4njZRIDFA+XRfxLe
qWM0ViDAfv6b/0FmPrtwiOUmkK3aRy3pMjOcimu5LSx4KbgFMKZw1nex30E/HICFwpRoKHiRPZS5
joUvjSgnqd2L22ujH/Pq+6YHB2zSbJP1o6rA2IWchygOQ6810zM+raX1mDnrLWv7bM2bnYGQtQFI
YFwaCHz66B+5+JFpdXA7sELaePWng2VEkPRDd+Lw6HilryhgEiUJ2VFBL+isZvlFcsy9xLpFwFRN
gUUtWMb7kk4OWjCq2v3KTNSJ/H+FvsrquKBxCJJSrCq3xay+XOZxbcrggs8fvfz0wB/EGbwGfB0I
18ZxI/VxwHm5kBn+3EVIUuA1Rxz1X5AzgIzaUnIOIIvoZ9A2O0xcX578TcLWNDX45gMjsPcYJKnW
uYdcJf2iINgSW7+HzAWN9Bd7uor5nl4YoQuw3ScKgTJYIo7ez3yDqdZXSVUgnFTBwTmDIwqD2XNv
J7JiZ4FLzXbHNKwsv3GrR8cdNhnvqr9sG/dczU1H7zXMWfsr1TdUGuIx2G6wG4qIgbXLeXKSNWTX
0eBxSrFccrIox1U9DHmfAcpfU/yxy81joADxzCv3T2iaWskzkAdwMh+qgOGQ1H/luuqST7DNAOpV
/Xgyo0EWHW+b/HDkO1RX0esP9BHNuq7j0kCcmvwap6oiBvPdYfyPEFwf0/hIIBCxi+wiauIdjB9p
wfSY5kftFlYvuFWEVaNIJ6Pw0gqbjk+NPkyVgmpEw53FXmIkWC3BaHnKZedvkURhqSodUyhjYF5T
lxBkisSFU0cptSK5zY+CeUq5iCyVL9R3QT1jjKksPqAYggJ94gKwZjY9+kj0Z/6ptjUG9+T7NdC7
190offjhsbNLAtPMAdTUMo22ExOqDrQA6qrI0OEOmU4vq8ckwPGkweQYqPtCRPh8IVKYD7YR5O7p
OtRXO/Ewwnheq1o0OwCtg6kfIL24th1KOGFc1DgB/Ia2VlBOJQGofIPJXgQbWWk0BxgF4MJaab/M
HoZ0Og2w62+HHiL3y71y2r5dC2m0AorwANkHqjrtf7LTrMret/96XGc/vE+Qd2Dr2UNciXZZZ6Qg
YKj/Jb79OVv3HQUF/c3STVt8fmws18pBmzImpX9v9T2I1gBTB3GIwkKvq0FipHAsjSn5UEcPLPpl
7zDG7sxoBF01AWuooZuzpdMkXI7NOsXq4HNcezfk2ESTR2z8b+NB3jmhqUj9Q2dNdAPwiSVXLMVW
m/OC2B2T0ccRl3KyX+qr1dRM5ccCqnB0rJvoxXRG77BknD3r58PNWHYBo+mzMdTOuAcRnemDIm5V
YLaulco75NI7mDfHkcV6b+Lx3Q4sgD3JxPRaiuH0SOY79GiUvj3EbKDuch0OG+ghbKx+dXfPxuWR
6SEtqMsiaIbpefKSHckGcRyglrR3bPJYFQ5q0Vb/AH13KeLx9zn+p/MrHEUof2tJ7KIQp0+hrbei
phVv2hGRIXMzy23WutVz42KZtqGGEDdgXeQ5KAMUEZ6ZaErfV/fJ81FIciiJcZQqj8WnXC8LVYQX
3E37oEu0qGAQ/MxlcYsDpJ7MXhVS+1ITkg4u57pIrfRX335DOdwqakaqkKjpMUvBl6Qf/lAIGJG9
H5KckwtYt66SvsxkmhpmjixGQ90RL2cM7NRo5h7LJu1TYCd1gXpGuqh9WJXrem1Vd/IW9Ftl7PVo
ThHvU8mns45A8NjqCGe9koP1oPmM1a8rmCPH661g1paHcX1htIDm9ofQ77bVbzRnVk5QZYeH75ZS
FtltSelH2kVibD22rqwN4Y8UxiEs04Fs8x8to2dnJ9Z42sRxARgNnjjwjNyDFBqk3k5im48a/+QD
P6qZIMHS9aIkUnATYnZ8aJ0s4EizjxEbYaMcUiAIoiTMapOi47/4Qy0jSWIW6XC+qs1ONrS5nGpd
W3vZLg+YFLnBrTt2K0aiGUpQbMXh2ggxM39ETqv+66q5+5Ht6ZLRd+xqLdO+WKk7aV7vx0zo+XhF
obJAmma9jgIvo0S5DeBddsoYD8uCFjFNEjrNBlp5yJJHa6H6746NVe/jgthUbWcdcbbQFDdXFNzd
gG8r5ljl5OpYZZVsrsL/iqbujuTiDJiAbevmaBzoCzYsyZS+Jnzd2d9/jrehBFS2mWJBnep3msq+
gK9KD/NnjGsSa0y/5x0sqwOTgdKVqKebbYNyyKi8pGk2quWUmelDwIt6dKGoN4SvQLGZqPH4ANYM
WPQlp0vz0fUrscL4KDnTu8qRgrOxj9iFIodzoXd0j8H/3n0oDbz56twi4wP6iCi/0dLLIDYhDqyl
JH8Bwlwyd5SJ4GaYEdXbEcySEFbLajEQy27Wc2s+0laklT5Ip99eKoQyjbQD0zuWmp4b/ow0EGAZ
QROgw3RoC/BGOnH0NBmW2DWu/GzMiT2qiW+9XQ5xQGZUSAFiOTeLphv0UwgnaqbpABX7qCaoRbaU
U/Q5frATyc/YbtHkCMuPz1osn1JFb0Rw1MP5it9FrQRD+cFsMofc9KZpGkj1eMOPCmV3dl4DAi+V
fUgJu3Bp+6xMCKXCsk3YyVuVd4oVCSdWbVwu38ibS5xL+TIsaF3e2I8nXGLyq8yS3F1GVQ3i2f+s
55teC5gD/XH6tgoArcEjOWt+QBEEHc7ng0zNTpGabv74kiheREYK+TjCKdRCwRUPrvfLtPpsxUXm
B97tVAKhX2q6n1xQLbDSVDWv3z/1x+M03Gvf3Zux4BLTCiW+/H0n+2hgsBwgUg6xpo4NHwm6n3DG
j002P6/2I+XEsLfwsxOcM+EBXBoUcvEkTWID2DHYP1HwOfF+rZ0hPfift4X++fR7guEaeMVfm/y/
f/1ID0DJLyS7t5lOq/3IxVwaFul0tUfKiUv8rNzbpzJfWVJcF0mG41DCsMgxyDlWGj52C7OoEsPn
+8H6NLXMB89gXyTJcOSXPbHPPGUF0jO5SyZfVL0nnGaijs0zFnjj8nVHJrdrTdVTSR/EIinJUmbI
sbg0EEKP3WmOJaKD75udlVo9PBRF1qM9hocMlyHhO9wHG2XkWXhJQByVFa5P9rUOiduBxnSB6Ukl
8MgZuafMmFWlHGg+XVMRymB8QjUcoC6pFTvHvgVZx+HhchasYApu9nyOu7lhCdrTz1SvkyqYUvWQ
eYqDipFJoJUARFxBzeUPmBn6/LbVS3uMHVk5eyPM6wEdt35SrgTdGKgh4uQdM+mD/tjyCSBdW3hb
eyAA079X1h2XDC/D6LljcJDAKSYP25OduCQBzpHe3dQrxU7LZCbZXdwmyVoKz/WAwEhF1nMvJWQv
J71h3MfQbd3Ba29ABc0JreDwDeysOy7KDJnXzPnCiolTGIoVmM7t9J3xdFFZ7bLJ7C0YX/LzhDLh
PYP2/w7hk8CQ9njWDottcLDZ9OfmBt8L7PpiI/6oMuuzFNyDSCCOStCdTbiut52k8vkPL/RB2s+c
EG3nwGBLKNLTQ1WtS++F+XyO3xBSyjM9y5agj8sGwpiDIEjaIFhVhhRK5hJa1bsGsLSjB5Rv2hHE
XAFiPZZT0AQKWMaGdayxeAk+h/He5pyc68ByfWq5d2ZpPk6USw/uN4sHDRkYscL3nrotCqCX0nrM
MD7ksGMJjeiIqY98aZlMYvmXB58SQ2VTQ7B6q3I1JUqm4fNDXK0k6PUxgMf6ckgQ0DC5W3Kp1Qzk
Qm/XALiaUMFwb72HDU5kQOVXOoWyQTyuWLgjYy2jg158UPz7ezbZFfRlLXB5imp7qVoU8ujWhxKa
TljMakGD7mGALD3BBCZZV77+72bBbmTUoeiR4zn/lQunJrQrq2bEQL41dgjgw4vTsAwB+JWfl1uC
PXmjtUw4B3LYr3K5jw/DQFJ7khXlQNBYyhQxqKjkvWc5irf+Y8+KAMM/C1q4semlG7NGSI8+jE+/
FqRVgiywxOnXervL/pimcsuo9z5ZZ3fHzOFUyH8kR7pG+UqMtakuF+5RKAPHCUiGPoU/29ZDbB2Z
NzBIPwAjrKP09JNTAwUeQBsZefTqcEMjweBxUg2W/mZQD5ftJ82jK9I5u0HRrkf6tBnf0VsQC/ve
O0kkCsZJXjHlRk5/8kiPP6u4Mt4fiA791yWcsKLe8SQLWmqvjnCMS1nzQub7em6S9zYXHKBJqm1v
ijeycNq5DcXXMVtqUTJ90J2+Noj24CjbCcRTxNjpaK4+rY04vQ/HiSGgEwLhDKURslKH0solHkzO
RuqfUeuJgFz+5S/d6fYQtVxXeambt4gxj8Ol2tPBB7aH856ZnB83PxpIMVsc1VEmhosLF2RGedi8
++FX8ZUKn48uGr6UXrj4VB+6hkz8SR3O/tkZWU2dykma6BJRVJONti/x5T5aFX7yaVIf+nyeTB1S
1EYeFUAZh5QBfYB2RHCCwMqY1NhYaYSjukexFysqcTM/jYc0BZuiamaKmDmtAJdFkkx8R4nVydHG
H4GWyWmV7oEGjWorCvYczdhsZSwrOqHs6xl2nBTTxFguk3gOn7yETr7kjlxuZo2ulcRYcR6G8bIo
NugCKaPd//8t82jip6evCrx7ygGIh7Jp/7RJo/XsBx2zqSgeBpPlaHuiUiW72efRHX7F9Mc36AoN
GGQrGuY43Lk0EUEvWUdW7GPPcLIbVykIew31jyCCSQAEnhG9Jew/QgLATaGcazCIe/grTOSNNbUv
lJ/AkOl2jl5IgK9zERY36tLRwfvjIv5I5I1k/4aiNAJcJ9o/d4AWqVDX7DyZXv0FJ3+LW4XuYjKf
pMD3t2zHm9joY3rAFnlZwRDA3c3hS0COWKsPuo7/dEdyVaVGVL0+msD7n/HvqeMWzHjf6nMrOudy
m0HsqELuX/daymqiUSfqUbt8aM7KH2yIG9zdiQS/GfLnE/T0JtpSocVXzTfjFyN0ny7saYRbmjZK
Tf5e926XjTNbwoBuuhcYqnleAitmjxvH8w9qdQMAGJnfezCFHKR0ss4logMGvy0VjqYeH+Egt1LH
7JB+UCdqF0TGLAi43SFbVjy6rkQLs7wbUECESFmH12KCj09D2p5EN+iMDnLlUXnB04QfKPHPokrj
GIimiGQ2q5hyZkOobwAx0N9fraY2A59WqFSKE5X7UKn1zEEOnY84HcAUDPIUmcsDRq0FhdLqPJX9
dGHyIhdRJCO7J5m2IwhmSe0NN4NU7f40kzx59AnnFQuMloQfS1HMsP1gy1UzYrujlWo0aTr2jTfE
IOZEpSXh1wUHMuvigxiHArIT9cxl8mRDxylC2jxux8B7elgRLznANxeVi4iTsIKu3aEJKvfotQJ+
WI2E82W1XwgejPCUCTuXPR/Z81mmVIrgrKlDf59a+bnKZIiU5oqIb+WzHuf+K6QtYokq5LOtgoPY
r5IJfR/MCQ1TKyf8qTxiIKIOn7HpywfrJSLVBFaamxUx5UQMA8om9j/AC5oNkVQQ+0hhVnT+9QTT
p+Ui6bRvA1TCDt1pH4GeEcu+skfMr2ZSGXx2uoay4PA27BH/PikjVlxkj6f4zvotOQpTtwJcWXRk
JRQeNd7EEiRcA+GmRSoKmQ4EAJVIEvtvZOoVgjcd1tHOlRlo6iFt4Cf/4t3SZtkNR/NugaMgtKKZ
JrloOUtgvq84DNtxmaBuwjEtf/vEIQMXxMfYpfxIoAnRLVntI0ug7OsWlM9n7EYCJkj0fbIgR/Gd
+YiI/nUptuBhRlX1bwp0FHXixMLMZqVKACtLwB2OXD+y6otjXJAkkHZZpV4BwIV1I9i5DX8F/90o
ZpSobLlfu01NgVkkiWMLv+5tIg9zzq8H15cfPxmOvGDa+xdtca7YnG9uWVsvyz0O47sd+Q7n9K3h
2rzWvBqSNDc6cCWvmqjVhBJLSbtvu015lWKgCs7lcbooeP3Rn6U42jHVcM7rqc3z3Y5+Be68WOPP
Q9eDr9ASzHxgFJqqP5xH90kPx11Nn53Gv/iZ2i6QFt0WAADZlUAgXT6CwZupCpchY07Ed4a5qjeN
RJ1dm63bSyZo52uZjKL+lGZ2aSJA5p+COaQmPQoAKGtrUwM1QbhasaQ5z8Aq88uUbjgZsJb9nw0n
Tpd+c5nJbLOOwZNFaKtPOc2CQWccRiuvUuRDwtd4n4cvERhcVWldN7xKZgMy/2lizsh5N0x+ZxjF
JXqzDBzTSc60kg5/Aiyg7IeuY9DESM129+e8oIyN37yZ7Xc4xdc717sCTndp7/gKlU4xta6ZLgTM
f1LFMHzMcZy632XWjIWPmBR3IPrCJ7N+qVklvBQbRsMQ9wcZmuGhajrr7LVw+hv5FfArhdJK+F1N
sXZr4vAMUhyiDnB6tOH8AWRVqbkyv9sCdfKQ14DVF23BXzpPcCHEE3DRkPIDO4lxwpG6/2mxKiGW
VCzw6s8xGp2DdxBfpEE9y01ICGuueEP9/F/E+aWDZaW/g65wh7ofuj/pggg/ccQq9TCcb02de2Ss
uRTbVYSt4uXRAkRii3EKKPmV+Xp/i+yCWJbWnVPO9Ax05G87e9o9PAH4oDNnUYgBAXD7IyVI1h/v
Z4qzKMpArXV3dSywJSquxXIRd5MzSeFabaPN0GEerZnZn58MWh1CBpq7KLVnAvmT6fDySU2S6yuo
2Scojr51I04LOKtnFtz2xzmlgVgNeY/RDytgS5FLQrhOpzpVQ+bv0NEzUJTkTZKwhKhuIHuJ8+mj
4oCDs45hdmBcYgINJ2lUTkyZ0390Qllx0iIjrCgixv5S18YM3PSdmfqMgkXCWp4uinW+CIwMr6tw
Coe3VzHWVlAom2rU/Zffq3fvd1uGYRPnKfLdRssWenDnOE97wg6tBdmutHYtbKmR4aGQ6qqIOC/6
/Mv91LMrJRow1j7cWXd9Hgtq4CZiZ0YAmXIqsYh5QHpMtk2X50TfK4MQrrOITltweIxPjFE6kWp0
SxUpco1Sl9iBSPZb8q2JF6K8c7IA7w36FVXnx8pfGVWmYkN3u3+r3tynwErUaiZwplAkeGIXjnky
bS9i+bekxXw0cuyszRojc1UNj6dnfn/kUOOyAssBTnWAQw/nkUuOGx9vSWfSBk6KrLIQxlu8wrRr
8kHpquInZ82bryLzhZg+E0npHFv/f2gNAkyhp63nmZjmOapaohmynW2I07VnZtTxTAxJfki8oXmS
810tEh+652z4PR+iuX+07spcBsK758b023q3oU93TBUdrXziM9QWB343h0xYX4gcaz53TTdcIH7n
P82L1eAOUrOpCs1FNmvi7gATGZ/Zf0vPq568ssNu4ndGxcL0uAwEcvJ7353i6gkzCRiVB8Hc6JCn
kcgbK8dZ84aEAlLMoHNJ05bNEpAeytuY7HDOTKF6VZdqdRNc/CcHFkzfkjcwBeXr5J3lABm3yQiJ
ZVFM1+AEC1k5HoCJscuwfU7uzoXas0yU/Zs8QRN1vsQlLStzPAlVFjZwW+sb4djJhWEdwYVTfIx7
kUGrUVMFNxm4QoJuIv3MSICGq2B6mwSQdhlP9TYJUJirXX502eOyMvt6ICluzQH3eGsUk5q1oEAH
DhVKze6zIZVDP6bwji8MrwSH0uH4dcc7aBORf3FryK4oWvkqFlcribuZVQE7s9kvb+QdcfmPNc0y
sF+CB1KMd0sLMVhCfEpRCNGwi/8zngb+6s2A6aY8aHdEYpVguOTajZgXtY2H+RnzFx98UcQF0U0B
/ji997C+9i33NpeDoKnfkK1xdzUP1XbzHwGMjCc0myIo1cdQGG8Dzy3zd3IJIaHRB7Clt1vgbpJ8
n7FzsbjS75ph7Xmeee2KqoalC5r/vHCZLxmayzAhgTfNPj2CiVkKA+h6PDivohvvGPYEDp1GdxAc
xWLxQBdI2/pyKyE1z+yztLf6Kz8e26K0scHdS2nQsnz0uEvD9F8/G5gGbCEi+lgCVGyXJYeBpYSd
V8wpm77mHGqGAvPp0/rOZhZmsNaVC0vByb0OKps/5DXEyaC51r2DY4q21OooKgPqWSTem6YIBc/c
TQccp9tNJDqAt7cXmM8wL01i9Tx9M0c7tmcthtig45zzd+ASA7xZY2BvKa/wmYz2j6NRQ/6BkcS1
BGeQEZXQ/cEmgwNw16RdFO8w+8hINu6NG8QtHSW4SLCJVA4jYjaXlLQ/X+5AQ8PPeO13dk52wGZY
kZVOz4IzjIPUE3MI9Bc4UOHfUFJVC7dNNsD5m53UAvgts11wZ09NQvPvoHDPii2NY5elCoqYS9kJ
YDaEJ23hJkBUp8vCAw67myMFwgCNuYZtHWyESlzwxelR+G+UIbjNsLey5fRYghxVvwbVjjOj7oCh
O55ltmWGGa0ZvFVVI3FKvquOp9lUKm9rfBshuiALcR323/eM9gP6mglcTmxqKYYkoeYxiZen7MGb
wlv9l/ECVKEtVPdLeKMUquy7XE2qkdEC4uUNdZ+ASfHnxCf6QE6fTuuMvVMMEORIR827xyc7mMeI
ZeczxgBAM2XD5JORCpbTtQvMjUdINFSanSYG71ZULJxVEpD8xpIGlqYVyj7TajSqOGAaDtTugDA/
wwBQ3ZScsT2oaL4/qD9qzdtj/h6UkT/zP9hglL+osSR+GVb+ffHcQlYVqx90EAPzKD8bOwnBxa9a
fVHL69ksGk1FS3vXtG7+t1jMD/0+c6UaYEgacR0LeQOXldyxaPAmqjf5rhY1fNTy2gYWzYgyYG96
8j9kqxJPiu/iDz1UHnPYooe5GMeDRfaBtOhqpFGGfa6h94IMqtf0t+GNpFaDSaUYYetrW4pesbk/
uTlZYQnsTIuqcgs/gsgxGOYXbMyXEfDVdza6eHRabyNcbkQ4xZXPCYG4mN9Y2ms5CMqAu5z/YYcG
gvyzZ067VPlPoK2B1+O7eXUPTnnBvytrRU0aRRKhBE8X7+q1ni1SxeK03DtNFsvXoz0JJ4IeM9Dk
/JcG7PWNxBM6/rv4hJ9t/kdUIX9FZkXv1lKXyi9ntzqUHKS7w1Og/6uZ2f4f3xl/ZLGsC1H0qCPQ
aMdS+ZGdCUOVf8j0WycOzf/6u4LGwjBnlAEhbVJ/Y7upt1UwtIg8pk1g70LRpanARGmYvOxzkjN/
SKV2swImlmXXrlcYgJoNoTdUrVR+/skm0teRLX1Nyk2Lu/GX/ONeAYucCzrVtRvFWVncBkG/kA5+
8891YXFcbVbyMKiQqlqF1YeQw7h1LTd5WZ4f+KwltZ7yKTieR0gHR9vUAFVMYQT4RUfL0/ikqdDl
hDh1VEODl4Jf0ydAV4l8UmI9zIsTWYcjmYwbhheH/O8c8JDjosmtyFm423WKTFFFYkxPLZWjwD9y
3J0Y9D4VEsWPCcSJU4Lj89KK+RmZ4DeTZp3PjabcgCxVebllN2dA9wKXxcd9eqAM9ghY35MHhdj8
YnoMYsCURo+4EuhFx+L92+AO+a4RMds6CFUcs6nD9YBsi/N9YRwsKL/RATiS0Ae7OGU3JXOW7o5G
OOWBxj36leEWYOqb8HxQTJDSk1m+7ejDIbWEDd5dtco+U18MaP47uEuY4bGEOQHU8BUXGoBzEcjM
MzSWjDAZRYOlrh7JLvHOxyWWRm+b4Z+XmRNMPlaP84d0g2ILkmTzzMXnSTvajY3wyil8tDCJnP93
pkWCukp7maRuB2nhuxF/uphRHansceh0MD0YtvBqhtLj3I5bvFZ+W1i+VXUmrVT1d8YlfA/0NwfC
t/sSWD3ns2BXlu2qR+FImJ6dgrI+0HC3FqrT6kcSmNYGWcukwMmChaNmS59K12ZcH+Guy/F2+p2h
zl+zNkNQSEEeKJ6wyu+kMS/VOOL4SgM1bhWbYMyZvnu51ke4jz5YpkVFncFZ/353OyvDL1JHSHE4
J08HRlGCMArvs9538vFjIH1+jUNREkBoWEcB51hXwRM81PX4b03KvVmJWp+It7sNa0EXrG4Z4DoZ
Z/buNZskEEDlpXYUAwAmQUqLZenGikzvlIiCYQPReeqHWwWj3KqXnsoJFDAo7v/lgIiQuPB4lk6d
P/TNkZU3zvzekA942Y3LGcsD2uckPGN2i3rX7Oy+WSLdlhtpGz8io6LbvYJDkRE6GiuQwIq1fX9c
Ao1xBtykaUqlZZ1jWEkEw2FaBT23sGWRjihBj3txzWQioGN3UDUEP3goyZNUtXtH+uzNfPMRL34n
bIHPPzctKkut0p0ws1l4NnDruDylYgZytrTuRbhkUvPx+YSZKq8hM6tiCO4CqZcc3OV+5X03ek0C
wy2L82/CP9GG148PldPa/4izOI8DuFBR0immwzeFVRfMQnbiJUqe5CW+zIKXMa5KR/QxEkp7mLRv
Th1Whe/50fedP7cVRnZKNOrgAjTkVa9StZAWEO3Mme0VpKCkPNP8pp9J8P3Ig8ALngLniOsRsq34
bQexdbQ3feOqoPN5DgjieDqnp45G69S6Jjf2CH8TwFgsN+nUOzxU1BQ9+mIi2viBO3vRYQpkPGBe
4NXWUoYpSgynipMmNFtqlmBSsvCfEhusUxb23rManSGYC/LdbU1ui36yAnFOaaAQRympKapFK9gm
Ee7HmP4PYmik+x0wfp/EXqOGTXvhpYvmBCB1k3IBQzZw6YtCnFjcVJXx8Jn8eGhz6yloFQatU6AC
q4ILjm4yWDRXP9pkHEUImQC4uUhrzg05pqs7OWVG8RgDxY7nyPtVaaZ+fQt+VhallFA9eO1lYUNg
yMOYCGAl6h57i+hpF/gya/FJi1zeRubzCwaI+nDCznhNMwHLvWceD854wzWbPl4QyKeVAzCjVx9y
aVSyZEiaScV/JY1bRirMl964pvMmwFgJcghhB27XwcBRHcz8grBNAAn6+SmC3MwJE20pFSMqpdK/
54fK+as/MS+X3EiwCHnsxavIYi+3E0FuKxGEYWTg/+7xFbGvUsXn+v0SxF+dxl2fHZRn2+ZbLWM/
/OrQTTcuZKM8onH8FqhioauWcNtqBGnZUCXmnKUWEEhb/1T2eCW7DOp/uMuEtUkRLtsO9xDtQbWO
cRWiiqoxciMMYxmvNo3HKYwjcTCzLfLcELO59PrKCPR9xEicHZsM/ulDUXXMQWqJjZkC/X4+zK0E
ILQU6X2lEv7Qlz8btvUi9CKO7/9oZl6dCspz1F+aZ8FuM/tPwkYnVlEv/0ed1i2SZaMM1ShBLCK1
EH2OeKzAuuFqjlwtXlnTvTQtt9dj1hBoQQqIDs5cDUuFQ9SjR9DRz6X/LinXcK9Z5jMoVIqHk71s
kuZb9NVVJnaRxr2IPv92X9OnEt00xbZW1PtLYnZExZSDnc+wuQUcoBRaJJLkTpzfIa8Nqneih+n+
pd9fTjpdo0GHGGpqFEteS6mjSZh6nyGOto77fWPVbLMEudlVtQmTeZ6xnbx1bSZ2dO7QuuhJPh/N
0L26MBq0RzVLrY6X4xVurdJTA2qa0NxcbttvXzOmfRTBan0ocQEO6Zk9vD3b7j+mtY6SNrhdZJQw
QGvADSJfbFRfn8A2wJsk1JmyaIDLeF0FbsipRMnmDco/6JdvbtFm6XfWFx2gMIBsO3nQuUmNb9b7
mM8tSvfPMSfbl+UasMDugqrvz2hfXD7TcO9FNkjYbCmXKRSPO9lsquZXgsP458RQDyFEGOzv/lDU
hN3CpyvCogCeL2oWoHq9Q7i36XYHOrSUo8VafZ/cqN07+wQKVBJ++daM+5NInyq4eBXD84HX7xY4
jN/huRKr6JXb7l3n3GKF187w75xAn0ANYvLyJJADM4bPiyfimQjEVKwvAVE+E7bBSkvrmHrenSQR
60wuRVj6x2O/aZjDkHrFhTi78fgb+cy0hRs+3xEAAf1PSMYsTubsfQhzUA3wk75C1gaISjiSidle
oNEn+t6eM1tTGuRlAyWMgY9vdyTeuh+MziVYSgwOUY19A4+apCrvXKtrbN0nxyczjIBDWiv4FmEa
dU0FMzDju2k66RLk/zcs7WPXUZ7FR67uL9IsJ1W/EW7xq5iw8FwE+PYRtMBWuW/c/gngg17dEMTe
9+YPE0iofaqZ2ix+BcbosvYlmeK5in9m33d5Lrl5CMl4UtpfUmiYf2JlpCNNdjYT2ClkT81q3diz
NleZg5yV12JuzVd69DkpgtyKR4bXasP2orkhtr+4mt23yK+cQpkeh0OSWra31dPBFPwWZHnTl/bL
poX+ecqU5tIgfSnBknIAwo1rtqwP/FUSA7Y03x1VpBoM2s+Ymr5RHKxZKL0WmoH/dDbUNRBdhjUo
GDAFDxXgtJyvVQH0QnruHIkVM7fW1Hl5I+z5si43R/JU6XtrHzWZ7+ZHwPr5+pnfiKnqQ0v5877G
s2rxeggY3HcO3GJcY5HMLnJA8HhGj78DbvFe6zDzcNTu/mNgEWgmsgmK/paJF3pWfFX/7JPCsDRi
2L6unsG/p5XxkzAiP3pIcuhKoDV7DY5GKIgR+CA25Zr6BNxtn0Jv1U6QxKC5d3XHHxjs7IM0e8os
9uxA0XtzM6mLGlyYAzjDhVeg4jHjej4MYqB4J0upTBOFpfCTrhCdLu8+yj6xN6p4SX/F++plVvhH
4+SPV3RyVM6WOf6tUr4YhE75zaz9RRtXSdSTEeK2rXLYInsRAYUkEgALcdymW/JZmJP+4B/+iwac
la6kvKfCTHDXNaHIu+FSnWJuptThzB2qGJNanIoTUBeGGTeFKkA4VFb5WlhpyH/yaidRH6StYFJj
jE/6mzJdolxuvzvaY3IXZcPqf/GzYGjbHOiILu21+nAgN2KlSw1WVywtyv+vvxWibGcLcuTJMiw3
ZCZN6bwU/49yP4gH1Sr26aVa0l0sIw6FUhOqR3pFVTvoW6ZBKwghobFsBeukwU5bCoIH5aS+6xLB
pCIceLXHK595ikZ4yN/1c/X1IRV0HXV2jL4zVjlcs/szUjQdAQgoXLAXeeqXsKgDJoipfLKFpYFK
Aj5LVCKSyBGKqbO7v7ufaC8Atyfs2ikjsd870hS8X420gMp8OykDsinGbm2iC0suuAT1MAdvfgOs
o10h3+eTpdl8j7P31XytogdmkAybqjDb1HOSSngRe3CrW+4Bgxdoo1BAU1CCs8oJjsqZHCfC3Fk+
tvlpJGEZ6nULi9Nf5FByR3E3+aigd8pn8J3P+4C6kbid/aQzNwBrG6bfgIO5UbYyaKoRdXSgpWdp
rMNdYb+cI/0TIUMit+c/caDmQMdCPn0d4uyXJ1eP4ITtY9gCX7uT2jcZbjYi94P/CavczGI8cBk1
gmW+GkjUNMTLu4rRnika8xPl9lyKr4GAJSjecMksZYunPMcUp0LN2Nb0zVfUAeuPIXpMGhecI02d
wpkUNFqQnszttDIpkbCqkd32+0V3mPJ9HR8WfUWrsQT3s35kKbfJ2qezBWztJJgY7S4GAna6CNBo
E2FQP/kS5a5QA90xvaThw0HrDPTv7Hayeejkmwq35HW/c94TXaP+lwcCmg5izY6nGULqWigP1dsL
6JQ7fzbSQGG0K2SxCyJfLMwwGeX6bG0w/oSJIWhAkuwI8juo0+heN16tKdy3k0ZSCojqRNhgGuku
oFVwlrpa4R809W4Y1y7sUqSDiZSKHSb5UOWQ/tMYz2OgDaihKgCmFDnaFnFfgH7w6dsej/zweqLp
iyMVXXUGzgkMXfPF4NJjq7o5iQENjL6mRUsAnrYPuNMeA1KjBlFwCckGW3oPsjuWG0a8RUZhNvwB
fq3jxd19VoH5hJ0UBnobxyizMTEow+nSX2QTr4L47oeqyPT7p1Ge2jprPExMCeqqj8tel7rQw/fs
0dlc5vWv2lb9EcbDcvcoc8b/tC8iA6qbsri2GO/3DUz8zIGnpaNmhqQ4UuI5gzMEzQU/oAplOjeD
a25ZM5fGIQwlF7AwJh20A7Vi8fQKAmiMdPZAZD14yKJ4SZDThffKCps+Y28fTIAfFCkafEAGQoje
519+YqE3nGCuvwkXhGTZkz4O7Ui8mCG7Q5PoqtZrGwuR1Nw9i15MMcRVwL2fIz+HQgCB/+tbmDGA
aHF5bkLgxy++MvWDqOkSAwd7UcgZqCAv76FeP1HfNK0IFpzrP+kJUxqc9yBMAdIbgtn5DZqbB8j3
6XPLXaTXXrit4O0xFxR89TO2y4TjXFJCT8Eh65EFlzaD5OaDKeG8m/PL/0B8FTRXoPYBEZBnoDvD
7F+xu/oVTFeDMYcvYVVt4CdRwWmot6XmVweeToFB24OrIe/wINMDOv6kVW44evQFcTqigvgu6EA0
YYgnnfMjdyKUGlPhD8vNaI4yUEaKAqN8i7cfTez83H1LYIYViO6fM+ZcfsSdSv3N2r1tV4HdTF/M
RxNJ7VWRrYI3YnMfaqDe+du4iDADmQPGaAGHzLg6P84XmcntHewC05uRBvOMiW0HmLCMBQv0a+hk
PcXA6Ni84bsu/XWXumXopbQuefFlMN0Yx2TUg++cBppflEZMq6Nz3qh9K7yS27SUnkr0L0gz3KJA
ahj+Ufa7f13yn1atvLgXJZylmgAarluyp9li7UMDP2KgtPoaM6k4Q67JE1qfJMq1F36dRicAbVvd
NhAGIKZ94pgtilSN+wyD9+jPPNig6j8+aYRWyO4BNyW1N6SDuyU224g6976KYR0L6b3lteq8Q4RP
JILuxfKnb2dGbLKO4QJ08dEdIx+CFkD9uSs5DyKMGXIs2qgt2OxPevTesbf9JylXsdXaGSLpK6ST
vnqdoWRIcU5O7erYqesQq2Qc16+dGhHMxtz27rnKk21LL38i/LR+Pav4rHeOGmkNxULqJZEAcUPR
LCA35kVyWkuTtFVYOJU9klPfpgymHrAMz5WOlc2Bdoy4n4pXgitvBxjTwsyfgT71+ABL0PZQTfdd
jXgbQ3Kw7qMLQrsLLZtMVu0Cn/OA75dHleCZ7Ijqm27F4J5mImmCMKOgY4I+soBomDLVwbcyIavJ
eAlhUmNypfrq2zDtX29byCHVTdWsthtlHSRRHE0Ke2Ztodh38nCA1O8zxMyfOlSyMDtQzkODgkcW
wmAus2IhUn7XLWDeXVihCSZNWNos7Qa5Y2wJ23qpgdYIo1RE007/DZuYDLcvz1YlDOgdhCrperaO
axL2AHOwG5Z8YBIGs9on2fb2ncqx/XTYjyOi1bgcl4k/Ucx+MjwBi55dwJ9FB3jxRBt/vHDaB8Fp
3sALO+SUorOvVHYfdNme6eQ5qOTeWC3TAJb6rH80WKjWm4FaO3F2b/T1RrYyVHMA+d4kPENQQWmB
sSQ4JVSZr3Zme1Wk+Vs+G+LUiGjXs9X0hISG+lQ5OZYZEKzwBKmclVjFP/dbamUTlVseINbC6etq
yMTsiP32+06VoJ7Qht6XFDwi+brjMRzKKYwuSuEY53tqi+P5fI4gekLkQxqLkZyGwm+fuxIBECSe
5yBzKBuT3wtaGK+WA2vnsxbUbwplTfG8b/1zkj7LLM69tihTz5X4Yg41ybpgZUdujeuB99D9CdYi
eg+zvsHv6tY9L7oJJQ+7au004rfT2eHJziaveowiEeyapGFXKyivVnUqEwDtkC3uKgz+lyGGA5pH
Ki/ORpC3pl1OljukDdlnoxiu5yJXTTUmERf7Nc/L7x8eTlwMFBfrfHU4Ojax7vvw+VU6Xc2x2c5n
yC3Z0fdshjFLnNjRod9eu+BwTvnmrzsuLNbp7AQE+Qu+Q6ojQnK1n8POdoK3zbNTxSaKeH1L+UrU
KaRh4X0XH6VQg6qjBV4n/oOkO8bx3t9MVHWFdir4YrhbbJhMt39WRAu8ik03WIfrZAllVT23bBVH
Hs9mbYDA/jRdgPpCd8Mq8Z2PUIY10IEdmgjm3QpqGBEEXXlzFf8zLWWj0AOjl0+QMUQGhVFPDscz
JPEnXcqqa7VLth12eiP7GqK3ofM0n8/FfvkAhiipkbe6LNcAAnudEvOxyrsGntcO13Rz1yW+57WT
qTPNdIOhjUYJ7Ok1O43WDwLUlvaYGSzkphFjehjARb23uTyzjUaMUOcMqOp3pTUJQkRyNe650gAv
YYpI1yErRu4rnJq0dSO+6EbbUF6zDncE08fr7PeB2SBCP7KQRhTJQaPXMlGX31ae1q8L74SCrSnj
bvn1FW9KdLVbPr294IEpskBmFsbAie8LoQ6RAUPcsFxPAiUZlL85y4d/YNtEpxdJYtU2uxb1UexR
CqchYkTboCr0zMQFsWtoEhDA9aitrDNoZj+Z6vxm/lA/rfw/lJuWTDVxUWpa7q4/JwBMvMDx7yLb
jDgT5s35Erri21c9JRq/7g6sfRyLHlTCMY36xW/DKY42erzD5jkkCy1NfqS4GV9UuWZUr8A1Ylhu
WRtEkdGskalweaK09PEd1i0H3N7uyQthC4rek2y4Zd1sFejuAoPr0gMvitUHddDoY73V1MTsZFBP
pEbvIgtqVv2x9nNnSOjcckIg4eKcsyHXgH18dV8r6nSad68m6BG6VfB15eGVUBWuiivYKD/GRc0r
DsyACaHoXfmn1zjhX1RgGGYm0FhppXDGYKCSwxctE7Ssybs+nwvCLjEbIo8CjOPILpIOsZkuy6HQ
FoBn4gYNm+OxMQSvKnismpazohYbjLOCfegd4aFfCEZ7WsNOHHV83HC/3wa/qvZZmYgcl/3btXpS
jSRNKZyXRVhDJJXCIP1rS/glq0Jj/DwK13fHR+a4UALS+KaY3TVp3iOcHFX+mCDx/LpBwXfsI7sU
n4wlBP2pzQ9P1AdG0Xg7/80s+/ETBDNPS/WTS6KM22u1pD649cYacNMT8Pbmeb6WArUuTwvXBxz2
okMJDbAIY1aI0YT4wZlTVBvxqvpXQCb1KcddNI88/h7km4T5RQaOqOxRc5aW+QMdypWyqOmorGhA
UzOUHGetlPA88Y003VwTa0DGhxmSfBnaqFPvGrTvoCIUqDBpifb8fcOFvVUBhyhEZu59PTqC/t9A
lxxFrJHA6jLc5NYfXtCmSRSSeqz1n1JRjxBAOMFOMhOLTetn6gxwBNJJNlJ+qK2QCe8Yj1UgxNDe
7urGCdpVKHuq1539RedkAG+SI8q0+DUerVRkYL0umQAh7pQdJzwWAKo1Z6D3zwk7KSH3S8EvMrV5
MSAfBbjeM8YepHilQnnU5UpvR1ihuAlPd5gmSXZLebHpQ1948EGxH744CSwgDkI0ObH1RSMqsR48
NZonRKSTTbv611RzXtWCqK69C3fsmc6hlPLEm96tB1k5kizsgWsDBuKIJlK0XSj2qXOGN4ledYtc
8h0HqDOylgbZA6c5+HtjL5BAZNDxd8TjsD83qI4hwI/kn4YIJRmkKqP6Qp75dA1px+Ix5qT7gBap
wnwBJam9RZCDfcxHEx6chp6zIE76074fZC4BnUeCQOnhoeVUFjemZlKobfHNVOvbsrYyQ3pA+gZJ
5hsB/RVYocoJxHDead8JuoK5kmxPo5LYJp7MtMVgvhCbi1HzJbYk5toDyY02XwELknf6WeKmBMsa
PspY85fS8Xrtjw4M4CpXcY+81y7KUbRk8t4uQPloSffncmiLoYEFTYSDkZikwlAM9V7vsbwCJMag
5bNEFoCHsJydNJlMEFQFnwdTh9XpbsGYOWmq4AE1D30cv/6qtgkyjGsBHtzJ77wopOR1azgcWRns
GvTtz7GeioySwswxhg2wnkDabgu5BM1CaCDbFjScteGYu9rXUMBjitc1L1seyr8Z8vD1wfCENlWz
4lXXKXD8AFe9QiD0BIwWh53ZrIc+m5GpMlVc5vKF0T11SGMVwUUJpwifM0Su3uIYz8Pri/wT8sTT
ryVMuPcULgTp64pHIiPoRrgrYiCokvA60Pf8HKKYASlcaUIIMZ3Cwzf0hMz6Rg6rlhVF0xYzTyR7
zFaWBgyHVgd8Y4JGCc0dp+eSY0d7sCza3zuHF4J61dDpkvk/kv98tWUAXD1SNDKw3oEy+f0wk+Pr
6cx3XsjddW8yclNjjdgXyLM+DUKjfN5owOCZ4YkJ7Z2tlf5vH+v0jU2822IQiWS0puyDcOCPpGb9
Tx4pf3mjjxk/NP45t4wFsFdR/GnlBvw6YJhaD7I0lOrB9ReyNAwfQ+/bCEuFb1Pt225DvkcPenji
jf4rjh5x/jGGslf6RWSfD29OHBvMaRWcqMNwHAPwg+RZyRTR9q8AK59It1IQCVqOar0SEKZwWMKO
6YCKDCnJsDkLa2S9spKLajJ9yI3g3VBmbEBR7NgJBPPU2HTZOCp2XtjIJTqTQ0KLBKHYDJBrQ2zn
tE43lXQOZ8ZtdEWgCQuEHFDr7q1ceSc8O81k0Wb+AzSzMzCbUIVb+7dDmi3pEHNOj934koz/ReHK
dwMou0OilJnvmUwrBjxF+S+yLYsmCDwQOB/VtHl0jNuvmHOaJnUlbBxhCJrYYxN4FEjfczrEpTK3
/0YM/oqaomGTWX84SCF9Jlv+zLdn2el/oPfrbIb+e5KECV1oeIxH88svFhEeyhEdNBebZlDiHUjc
OkLKQeCArnGVC3AlG1cCevu9oGNbbufWk0QL59w45RZQvkdq+9WZIkmL+45uAoLYPYaKC+v52JW1
PL9ne4OT2EUSohVME5ixjQ5LIQ2UPivgfloHSAAjdWN5wJsbIdcV9IMBXznDXdIVcx3gJ+P+AFih
9bNoU+6sIdM6w3IrO/Ebps7c0ZpXzuc8mjQsdMup1Q7ckgSMJRGYRzEfj1YEF7BsWMk+v4NvYakc
TOsW+4ufhntpsqq/1di5g3hjoAEKaOOSSKU7GWKP9+k+T4usg0ICMFJBTuQzVkLu9u0ypo6tCJyL
tBgH3veZqz2Di0IGPfw2Mk3vMo1ZI0QGExDHmSF+PCkwUXTLPZQvDoE3KYAy3EspK7pbKpIrk0Xf
a7Hg/6FUeis9Q8bc2xBoWVsMBGOwYdTTbHr8/z98zs/oSicByvMSS9sqz8zwRTRgnM44Qv6vlyTY
eCZyw5bjMx/xGFzLYLp4p1VLGP26EBr9L0EHZNyyfZxy80AUxXv5FUmN0iLfkhZ8GCocoO6oyA+g
8JXYVQ5V67Q7vA+Fa818HucP1Q+AVdTMOKkonqC+8T6i27KEtwAZC5Cl1NcWnyAvXPbMxujkb2lw
1e5wM5lQE+PW7ci8tkk4dkveya805ceM3yYzz6fT4YSxVYOLWCn9g+Mb/E6IQ2PisGtHfWpIyoNa
Vt4LwzXBddX8IdKvqHa6I4dEaF68Tydqhj9bG1y3h96SI7HHgDXafhK/+n/q/bm2BBN9NP9Fxvxk
WNXsT1nT4MYcF8HH4i51zZYXo5yUZS/jMT0EhBrWWbHG0ZG0g+bdncZkChAa1vk4tzT7hhR8vxh4
g4ZMsfyjT9vCrq6MHrEz6psuRPCIxXKQDy3o4YxXZdLNW2xGELqgH7z5caNYQlzrgaOxbtFEdN/d
d4bIZcTSu4ZMlkR87svAyfZ7ff0Q7aeWRCSlCTNllVJA+a12Nne/bmNoQvrARaKfGSpTdocyLI4d
1aijFFu2ganMWjFWc9aF3M8XtkxGDXmbcFGlZVVFvMW8xwe5hF89KFF79M6ZsdS5uCGNEbEAOQkM
Mm+jgttGNgExkqUn0RS30bfr4hlUxcxgHMrGGr+MOIls8YDEft73NNH57xOEQyuJSA4I8o7LHIwl
NuTmlwbLSD8isnJG6X8ISGP7Of3rFugARZiXpc/rBwcjuCIjtBA51PU9tWmFeHg4b96167/5PJmW
3lu+8/I2MO3GeuW0RijSHlKMGhsZq5+i5vi28CQC3CbuoRiolo0BScOf8MqsbRTaqMaL/3jHl+KP
xA7Kv003kZ3tnXiVJ5aGOijo0zBPyma5WfjI9eWWosgdM/KdzBF7VH2VUO7YU9g8ckkXQeFyiKzf
RUwQ3wY9DtghCBPv5X1R5gWPgmHRxkiPwYxrJbL6+LxHQY0IRjQvgCvPCMxNf3pW8s254J79nJaV
P/NIS7qGczTY06g2y90CymcgVinCKf7IGbr26IcKTTs66R2LeZEyvMhNXiSBkfjKTFakpSgfdJfT
BgyWM0YxyWP4cpaTEA2eCKBPscIkL8cLtMNjiCsLrKumRFyQQ9RUDeC47v3WDOFxpFUH/uJwJJgn
ukf1QEjHnt+clSxedivu4eeSwXnnwyPQj5417+hCCtGLcpy40/PuH+nbFMc8M2JJLLznJIP2SJ9M
Xx5m4sSbhrDOSiCuNrh0IyHy2jmLtE7uy7BNMcZsqATvkxPnXlKPchtysNXavn9EpDgHysiSLqJr
uKJJo0IYiP1tYfWmxTejlCG55VinzE94TYm35a4fsqjdRvlj8xNOrQZyXth6XVBw2l65mnnxoi1K
n3InwiF9K8aW7d464P50xz28KGVg+HQcdVrwUuZl3x0j9c6UC0aMyFggQ95eHr97fBHf9tWfjcSs
ye1MLE2t8S6tDzYLdu2ENRfpzJOY7Kr1RfqyEbUUcb2QTyR6SwuQ5sUO0H3I++8bBmpAr++wYbvJ
YKRbb0pc6qg+4/LU/Duxf+bcokoNuPDRinv0Po0RkKrns7N6x00RrAfrGyslvmz0WdeZW9C0Hbl2
YdLxdo+H831URL/igTWJYaw1clLDNtUARFjSQb+yHWVqVJnkZZ5j74Sdk/RfGm54XqwNO9dkB4W+
buSM6EqC0mshjkphts8igDrbv9d9WwSR1aF5V10tkeHFlficHHzCb6ozI2A7Qwp3KKXvcBr1FTFR
3v10USUVx996Y5ZqDeMF/+l8J9Z8qkD9WbCECS6HnsBYI4EfYCM1G5rbvA15c/L6ApsqpOPshQ2m
FTo4hRnExhLM2awSjlKugUkXZYIwEinmWDz5R+i2zDy4YH438vQQnolO8Iokw2hg+LZRP9umT3ul
VBiaUTOKdYy4oC/pw5gKlHzFaB24RCO6ut6htbz0N5Cun+6vTzhEHhERt7X8LRfanIA26wJA2ANN
R/4SWpv+xWblMVxJWApI4yI8V5HNo9E1U0SzCjNrzKw05oEbVnK3qJ83mZfqfhxl3YGU0nWWuFhY
58F93lJb5Sk7EBuJmo6Wu4M/sXew/ktW9X1v6lWDFHaooy4mc6VGgFyV2fPsF02oc8TPasTBFFIq
tk8AU3RCMktoGtIArzVx5nVMWhFmq8qp8KeW61qe4yirfhvNQ+X++uB/A/XXdiNp1yFqwze8sPkn
bpMNtKRVRI3pMy1X3vRJjisnr4BK+oE3kBSdRSYHpSHb4paeTtjMScbJMAMcWgRledZKsLhpOEug
O4SF4BFGWt0bglrTOaMb2yN+VXCo0lWFM1qqoia+5/FKC7XM6k4WByn1S4v7QvFJJIbAKIqOIC2A
lML5h3NVpHq9E+bQcgE9smA1Xx7yJaE+y7EeXTNhlU77cG4wUcu3V+zmobvxjiEyzoupjInQss2k
mcYqRMdGEHzHTYeR5di+zgkVgOIqbzCkipzZ6IjNQffqezGiC4tqG1zaOMcL02eEhkS9hOo3hq7P
9t0xJiY2WHfhO91xvaf0xGLeBEH/CLGQ4n1aSLFf/nrAR7TSPGDTna+A/GzkXEy3sATOpt/qfuch
LS7Zr8uXHdEwQTx4t0df2REyjnhLfhMssdVqh0TP8vadFIqYs530pB9zhaE96jr3yLWCcR1ZV5zc
RK47MC6fS/uBuIpZZPiBgWugeiltiCN1wiyh69+bT4DE9CbLjDsJIMUqf93s91Pf/3lSWpu3FnCH
ejn17rT/XvWCNoMsAKuQjN+dDAk6cF36krxHCA2vsJZUBLbuuSAfrVavEgeNRZCsbTnYAokWfpT6
McvMiJwxGyNGdOplM39uvjOnI8mHRKvzU02CB4PV0DKFqQmeI+MDgex39aQTiGuJ/scMzdOb8Rat
vHWE5MHk3hp1943lN8muk4x1h3FkVdFXgfuEjffExD7xEDzcyfvXGNKUzaJYp0V4GRb1fLpH9B65
PCrYIB/Bi+kMS4a3CYz2M6S4Loipureon719Q/OMJdvpUgNaLDZoqgFBfYP4nt3S8pwE2sT8CYgk
HWcRvAOpJTHRL98ao5C7+JtF8+zd5JAxBy1qFWApVv8/yShI7GGhliIa6plpjSH3lYpEav47yIMO
KS3dqFOLZQbZN2tpjj09tybL5LrC0HmJ4i6178IiVUyBUGNlD3UshUHqT1UW+zj7TWDW/ZKJ0aAL
Wu9LBGdSeq9q9Hf+A7EetQEd7MqnSsjBNN+ZnLrvyTHee5Qm/k+BU6JlbtR4/jVykF9xh90xoBhY
FBANwQGoXbPcAEdxQYwvNgMCoqVGA7spt0U4C1lcoEI9W5IVAjEkvAlFsfa05KTQ2XDHw4wBEZ3i
+K79V5mneXxpj8gEXla7SB0qU6VXoXL4cBDuOfVpiQwRVbcwkcJP502X2TdB+q5KrsOl1uAaEgJi
TEsp8LepiJhNckedApekhhm/v5cdxaD0rld2DAqpsuRV59tJjc5WtFI5CzqZ5+DPrqJvMJ3mm6RL
u+VIcWrGxRfjBstS3SoGan5BybwSvUB3XaAXP6R5zQNYmQJZ0ouesYXdah7t40Myx5IhY2XnSvfy
yBu0xfMi5ouPQFtBRT1aOQZdG5FMDwADjuxQp6OWSZFHBAncaS5w1vc/ikABviQ+SCSpwgsv5QW0
7gp0ccb1LpsBAwd3jayoF0OD4S/qUcwTR/D7PfaGt4TbkSdWmPWMjXACESUlu+h1C3N0xyIrjn/q
i78n1LxnAJ/aoKMzTo/3Lm7w81/6oJu0EiuU5wKs1y5azqlLHEdjODn7i2R9wOG45sgbQYapBHmi
rpu54YhMQDI+6ksXy5eQZnL56i2Y2wCIM4Y8hpW+XuzrIp+fkXFoQAm1HQbZxowxxrunDOtzA0vB
Kc/6l+bHsE4R59rN+K9VYZ1Ig3PuEHHPTRpCFi40xZwjoR0djHs9zeoc5F5oW+cTB6HyPkRxRN0T
1l53iKokCGChjE9xH4NMfoYLYK1xC93uBg2poKRRPXSd7HnFwJ2aMQb/BRd8kYg+KeeAs0MAQ1ia
VLYspM6hu3PMeCVLd3N6wvlVbjyffjEL/NZpLY91he3HUoxUyPn9vrfCqZeOSDJdSAYK7SUP9FVW
y3yWEeclE5YGL+5M41DImJiLufPL/vFQJhQtXGGaVRCyZmlf/+5e2Ws12JIvQL92vqM9Fp09/yfr
t8xTVbM4O5KWF60QOAP3H7g7Mnskf6uHju5lo1OnBt71ozQaLu6KqlFNnFmwvrML5kt6J7pS3G0W
+ZrjbziEUpLTb5LtDgWcoS2iOpqoBjcIjxJN9Bp1/kHWGeiCxCWX912opd1SUMrU/lxsVouiYhwf
2koM4JlqsWFWI7FO6yvczjG3uzIgTzF4MXla7s3VBG1pO7jGHAwORile3vv9hHzGsAx7mPnsT4yf
Y2A/aUyeexylajizWlrG7rUAERu1VtgFgAWVqCX8JdqKDV+tVcreKDdCkxKU8eSvoWrYiEsI1h5b
9nm161pOUIessMj5wwXaBck53QJAOCrIRZBO0HC4kOlcN70uUoCQ8mKVqXlZ5VbvYU9Z0biEUKFb
Ijk+h+Qsu5N2C/0SmRCigwSPASaR1Es2BBSzcsBR8/UMJJN3JFfGvzdqBHVgD6MYhmddIhDxREsq
QwTtyOCI/zawlnj9E5DhIhny04S4KjpKYGgw6/36GjymCCDkOf2gYmaYYd0TehefeJHnaUm8e5rI
E1GSkxOZxHYmoY87lGfUHoLSIGOtUvlRaPb2G53J+L29BIBWHxg52OgRalOYtZstStIbZYq5+Vbb
+IR+yZSr6nTgEvOR0oODzayQ9MZjwnufzDmOykQDKJqoPLbXmrX3kJmaYH8EgK4R4LbpX0yeV9Ub
yJjVOIXYvqb4A9CTF05Gw00wcjamqDqw9vkt/fPiFBuGF8yuWyHxfVlU2DuOsFzbWTIU7ZVOfVED
ni/FGotmo+MkjqvsR9vId3OImOgnb5ruK6tx/hLhLFX1kh1IzyTd7fgCemBeYkM7HoHyGDkdi8Dc
3jvuViKOXZF3ZBsquUSR8UxPoGjLwvvdUXDS1rlSPbaWpZ48I8vrpy57e3WfaKbDcKOeRL0Rfac1
HTdDEHQyiZhE7/057d4eOdneOcGwrYcqsRCbk/79jZqgDiVBRp/owj90FJguZHBcz2OoSerCQ++N
dDjRn7k/Ub3MR+cl9RYJ4NPDjwXfFpXvQHUjR2s3oDEIcnQITEvU4iDt6Xi5EqTI4LC9XVHr0XYq
X/L0XB48nB+waEbMuISCsSm+S8wfaiYFDEILgqqTdhvXki2WMijTv9kjgctXl1e3rhaqYuqHpz9m
X7k8PQiLKMlyU9rjHkvRUnJXz8Qd9MFWy86qFBORXfdXh16zxgOxOx4L4t7XBTnMtxCcXhDlvI33
sTUbgr7sFKbxMJ1p9XCMS4WhJ/liocJB/9HFDgUbbp/vyYK72X4klg7oX79RnrK4/bbF6Z7yfagp
7tmsPRXQOgL+MmXvTTkvUIhf8Qyan4LGWooeFdc4NKEmuYUjyrKMtu/kmDgZEV7s9U3/4jjlYrYD
69QqXyaiNoAduil10sk0ACGgsx4oAxbAw5N1XQcy0LT5Tus6HmjDYLjpyozL+dIm+udREtby6gry
b13/7fFjvdW+3KARz+5zvmCTgo+pb83HH+X9/QdoMPJNuUsLPDKHxNzIJH8p2Oamx9n6XKnK1BwI
9c8bSbtjQ6cABMlxSSoYNN5WIaubH4P/kNFk7DJ1E1zP47zknI7OIZBx0LjSzdXrNpIgOHzQg9I1
GbbYUIw85sANP6BsBP6joJDdonl6cPt9GHH5np9hmo6/Tlq5STjbKgfgEWWlm+qUZm3QPSE4poJI
Krv60P9smQi8OKq+tha2lJ7KNjg3gJqCuatSoJgdTQgFKxYCi9U0/DsUBhfZyEnbrsGtsPwW+1ww
fHMmSsWCJNbpHe2R7uTe/MlV5OonC86rv0ukeY0wl5yHZ3eSoxsXp5ZxVdKLt9DiNaXQdln8xY/F
CDN2zbKHUvAo1FlatsTD+tcD5rhsUoFmjDwF+WhLsAPDY3Mg2RtbFllu96kI2qmNLQPU5DZ0dNDm
QSm2/p7CRrxwP5zUXk0DGT2Azei/AngoyafAQK5cR/QzcB4JYyLpKlVAJJ4aAGl3pf4Rr8JkNr23
bYS2mzfn4URaNQr1q7Zx18sh4Re5rgYToRmA0LMJC736VZgZOuHxusy5XcD8bsaye/ZlLAkcxt6Z
zDFtL6/qXW77DL1qnf2hqp2Rbr8N0yC25O8vxBtQbGZwzEV5BMMWIWpX8kXQPrzSqWEkYgZXSl8l
gr2hjTIaJumbNx/RYAZyMmkosFtdMaAG9D+0jALjotloyLFaSLb+FYRMfooYhjrEfEa/wnWQYtYF
5EQqWMQSlcAPesl91INE9gZgE/ob7WkTvNhVV7b8V4Gtxwha9sXxkxDpqIbohV1fKdDtOEwjMu2d
1LtZZQ06uvzuoNHXHouexCg/GeoyUrFIxNhN7gZovqXj4jLfv1LZ+9rvbRS3N3z0cTswFg1PO6VC
knyhvarorxDZ9WTQM3KOu+dDF1ZiO6p/DNMD5nwC+50AswPkBhFxSgBMd/5VvatPpI1kqmkuR6ZC
hVQ1iH8Lk+UB9zGg0t/VfG2uoMT5NnwghwLTTna5Y3e5AEuUiWImY4uO74Bik3mHs68vDWVgIbMO
pjlXo5cZzwnmpZT9QtURlRAx2D7oFutfeBSnSWXTqPE8Qhs1RPXDSabfY4hl+SLnR8qtTtyuFSeP
NIyejivov09RJ3gOTETVxVVgsMHx9/ElcBnQjmzrn02StS6YEwdCtGSs61pSURoDOm/g0c0OdX4h
EE6Xqy6VwAHzI6O9fx66E7+RXbc6DwdxYO31DGiFuqGLWmz6Ocm5ltZK0jOY/vViT4PbsjqQJ47V
XCU3gUTTE82k8LEPZIHqEhOzliibkQscdihg5h7lXfkK4e1EV4OPUCchlLRJ8dnUV4FxOheEwFkP
TwSLLvZVI9SyK9R3Xr9wUNy+Nd0R+edVJBnAR3C7ylScUoSmjSx9x9fdpmar3cpth7Plgd0YMzoF
B9nzc0lNGYEsf2BEuTQnpJyXvQgyslJmaa20NL/kbwdaxYM2YaEEx+EMW8y0k2xZECD9RMN7wR6w
rmwir1dqQqTJTFEh4pVJUKCXHDHbaMNHu5Z3C/uznm7aayCUzbig/U+qWRaHW6XLHzC9VaxF26S/
SGAWqzmxbzGyjeD7SvjxlPQFj0YgPUA+VY0OYLgpN5CsyVXPJ/0l89j/tuLNvnljrWuvnucOFYtl
9jJPsKLsrEg7NEVplaHYug16uzTki+E5EiglklSWvGXYSJV+IETdts/5Ul5bTIstKrqvKsvOknsN
kL6uP3+goSEGZXwPICYtZ7iTDK4izFtSN6O/KBJJGBEyx5ZUbsZuuZ5Rb25JP0g098cwffdxM+et
K1XjY70MqahU1vWPWFiWiZieTYQSq2jV1x+bSwiVy+g0Iy0lP1B24G8sIQreDAX8K93YU3GZJwos
kMLRSSzyQMIHBtuVVHylALOgOlu+HLyeib5FYGQuZ4FTwoV+BnOTcuWYiXkF+YDALMx6acx8JHCd
IaMWebuuBIrosgz/Z4Lg3gZ5ldJm5PdCapYNFW/CuuzTO5qibYRpkwLBnIds8i9l3IaiB6x4i1+x
mPXPvVkR6VptoXebL/815H6P0wYycDhlCcgUFSpH+OtBh8/SdBEsgDPNNKqN5jxJkLRT5tw5hMix
laCXdNjICpZ+9VTX0Cr/QKPaiP0g5seQNpwG5wP8x2NLyOHMKvNDYdE1Ughxogb+c4KwaLTbfUjI
JvIHNHEt0SDA/zxy0T+vfOoZnEgL7QQysrvwyZ9tpUSeHTHGelUGo2UHIgQC/+jSa7yZwXizfVrK
YjtdzN1kdUcJEtAo2EOl2n2Ttjnt6EmxE0LuvQy4syZa7dl3B30xiKZIMDYpM+RIfS5CFxnCZ9uC
V6EjkyKrMzclak3iy2yyYN4WTvwlUWMphzAYMqBfpM1ldkSWVR4JaVdIqTyELh8Z9pz4WRp381OQ
trAnuXPTsTTJZBzMW5d/Og2FandFzRf5qipYm6V1d1kCjAvchvwnexw/28Ik3VUqDP6HhGBEVKy9
3FVXuj2JkOU9lLk1XzzpjlsVdteywJsTiRpuXe2PUjS617mEVHK8SvWaqtiDTcH0voy8IGV3uuFC
fLtrQL3xPVK4RkkV4peTgIO9bKqVcHtQ0kWocwMStTiugtmRTuiMCE0vSp3U7+XmPOR2bnO/atu4
izDeV0xP3Zl1qoEUkRDoNycFd1k6FW9UiIU5noZAAcI8u6OT0fwPdLVPpU7+JGOHuBhewTlQvkFi
Ia9AFUHyv51MEfghiOfTgSjM/QFhnyI0Z7+/R7bTTSxEbrKJT4E0YszbokNbIGL734EOUlFuIhSQ
oybaHWXEy+8vjtXGKYc718tx5rCrs8U/DxnKBff+cPHaFl9TE+w9so+T+bNkbUQMCBMtXABL5Uwo
f3Jvwv0OwIaGxklpsYa/1uh0/D3vi3EB5qw3itP/JSlALFZJr8V7bRKYtR0wruOcrL3QoDNFTAY8
6Rf9DEmf4I/yGJoFC5iY4G583moB5aXiuv4On4jI0lipY/JJv8JHHY7A6MdoUuI3nA1gN+VSOFJ3
L5KAQQGw7krQmaDaz/xLCW0FYqHCEmtwho59uaZLU+2JlJXZHEZesjB0gWnQqqOisZ+8C0pldOl7
TimcPk6r8LBN7nKRKCztgQzKOb0mToZnbq9mexi352+kyO25+pbNOc1lu2LzvBUpxudnRxCocgWw
tFWdIxm7hbO5k4QIN1fdl+rYStx9SOs5SehF26f1xq1nj+aCu1oHuCB8rgqmHRrOzoiwV75OpbgE
ZkoTO5wc5iLk58wLrek1akVCpBwrbzalNPg2IcTmnNZH2WeBu28urC1WFhI1lF7gSXnraQ1a0sAs
n+HAuifoT39gFSD22ZlmCbQYvegMs9xk4NEduwTNYPxIy61MN6A721TBhzbz8w5qS/KwttNjwkFI
PelYZaCB0FIAxP4R+es6GARgyj4VLkkMAEUEetNh5eHOOqxuZBCicCZW0ueouSdCPPxQNpCMEcm1
qt0ZLMZ6qAYXStqoZ1RPPoYcW7/VUbnlM6mGX9n4yc7WJRUyx0McHVkht7CWZ6D+cgr1so/BxmDy
HEt1cTYKw+lY7hwQdPZomdSTtxM8BIEtlRm91MnK5dohCCQ9u/jfn3+ZBEBOVorGJyjZ6jl0EBt1
1OlETr2oqommnCzEPMeR0ASlU8j/Lu/Wy/Jz89VXiYKoDPc2V16G9CV6p1p+/pnJyn7tJRrjnyHa
vzAHz9cgqd+ELxqQuS0V6AABrQXyrYapdp1SPSUjGnpz7khBEhd8rzvYit9IWytc9mgfBSjvsNKA
yOWN6f249lEdU882jcRkJYfKxbNwvcUqgSWNetBpzE9FT4hN7TA7/V5rDrlrM5ZT0Yp7j3hohwUh
/oIVQZWa4ly8R2g0DqipDEH5ae0OyZuZ8UjQ7o6PHeLw0I/4Ahooj3jCVa2vCvoWqi5+JXpvKKcm
SFMKJQRm5NfpkrC9S9lJyhgW34NQxD6YLzKG6R1rYJ25zYXjJLy4owHJlMoaXeTcVFEdIy0Fr8rS
xgrJAAYRV79WI5Fdhj3apRB3Z4xEDQdvYZxAaEabeG4H3MkK+myfq0Hj5c93BLRs+ZiOFxK0vPVX
VWKIZrTxKtdqt9+aCL5/0EhJKwkrycflXB/J100/tUi4MDruL5WBYzJZmgVoBHBQjGRLYNDeJrH5
GnN2uKN8lj4XF7tNUvaWOoo5W37mdi5rv1vGVSIphI5tITioaeWNZTwqjjHmnh0L1tbGOruxtgVN
RdL2VjIirbGIK8TGhK7H0rvpcBbARjIV/t+Ru0tEU3fFs6EOk4VXXEzE0fMsoyE8qMyHqpbcL+jU
PQXk6/esBhBLvwVQ6YGb3CGZo3IuXz87nlOlL5MtqB04YdjlnO3r73KI/TvqZa59Y52HNCdwmCuq
LR2HU87n9nYblyxXm4lvxQIzLhSPhUuU2sVeV8QZqpjGbDd9f0bt3FuQeLNuGg2aPfycMRwQWKgU
gd67RHYEfDbaoZR5cuKsnOVRAKWgiP/8tw5m1YSpiQot9KmXDa4tXiOIjP+/3H9TpAsx2b8I9QCA
s4zP6RKu/QlL4dWZ1ifWiyyhVw39byLiyozrZxDDaMAeiOozA/Jo+2oYi8h3vM2cShNgZl9+PZ8V
Sdn/lQKrT5HEHxcSQfT0yVFNvNssxHGR436ILPFrEBN8VRH5U1WKyxY+I+pdvISdmx3124ocxgEU
jBfhqkewaUsWzFFqSwY2YgObkqwFmqU1UvyVzFDauiLRyE8abQe1OVZDDKysR1O80/xDJGqb4fig
Ypq3ea2VeWi2RezfQbE0LTWDrmd69ZMhfn1nUwN2bngOUv1nM31izeiDtPlSRwFucdQ5fXGvCkqJ
FusaTtY0+uCgwXvXSzF7n01tPOJD5Bk1Fy/20KPmStVxbnVdMATNbkOvIheo0J/KP0Xskq5COXL0
ZEvWgAc1g0EYeeHfonTw9w6tRN/x/WUs7cK1ndXSuOV7FCIkMgqPNzN0sSHNFqKZjEyi9EQKgQkg
yaloiiExbeOTb7JVIQaUxHxV2ww54xK1njd77+3stiQEvfLUB2VWO1X++zfAe2fWm4bn/FWt2KnM
aiQnWyD1UzSM8EAxpE+ZLYT1ixYbd8hX3m6VAP060IZsr8a1g61JtO0WaLuYVYV1PybFEY6NnH6B
DG/UQxl1x5qNpyLMswRxsdEZD73Xob/KxjwPW2Esv/NrYAcnqIg6EzCOZgKKiynyuAc/gfnhuqY1
RMWNn82tgD+iqPGgxyLMpX4r3iZ/OwsnlUDJLluRY1Qtr6PfIFoxc9samIuRs/xJQKruDH539vEe
V+WjvM+EOGi/UW5UQr8lHpfm1w1EftaqGR+whIFP1AtIIjXqRMqTqpg9XeJ2FnH3o5/7GmW1NEpQ
TGhdlSKoPxlogx6G+tV7mZLYMpJthKXr1HYhjjSsZfSuBq055cEqOwCHHJzgJcRl3F2tHPz2idrq
bohYa/Gj17jfh8/1Gpb4tjrPVLucZiuSDgqnOyq95/7NfenkbgomkgxukOMgZpGic/PCpErJskK0
gvQZwPDQdXy8+hdqYfBYYSpBCDaG5QR7uDUTirpd77Rv/+nr7H2tWqffOO5S8RGaNBIUoiMECOq0
kqQXg51MIM9JigEKdMBITCfvugeAcrKaxMSZOP5oz2DDxJ1j4I9/qfWOzXP83PUl2QdVL1rt2fHY
2UCn1YqdUVo65SJpBbEAYaaRBkBTgcBsBAaZPndMxy+NuTPZYOQtG5f+96+xGGxna0AnCuMUoDuu
bqc5uPWrsFLY8RBQpihE3VverAB3bq44vKG77fWMV9KzEpBBT2b9Xt0pm948TTof8CGaZjUi+XVA
MvWOKYWfgTlFdYzp4/6IWye/8mZvUXU836yxJ0oJp4dOtLoSPflhuFs+PQYId0N0AYhHQw4UhMpn
bzgzcQMQNBsEYwNpFro42cmPj+xkISQsG4uGDX5xdbJcs05u9e8VYhtRbpCpbSZMQzgasj6YDXvA
SA07m00F2Rs15QIAte83iqLydyIoydghCeeKHX31QiCQy/2ZBWTQokA9cJkYUvOARxXr6teNorTf
8ZbuKbY4wG4F9YvnTpVponRTGcrTWTRrgBzJ4sI0aSEjirWhpplW1vwcn4cYood9xL1HkUwL3P53
tDg2bxK3yGILVuOmMJEYKp+fVNFMtRYDvOZ/4EVcRJlPaipLS1WY9RZ4EcbB/W98aBKLjajv5X2F
rT4OLOXuGvqamP5oudOPOwBHYMZW3Evk3hL+uJnIpQxJsAjxch8c9ErePiYkwlggpNq0Au5cRaeU
07aDlc/thysnoV7HM0ZG41yHayLIiyekJ4Ee6vyY9pLuW6gsyNoz4u9ufFRE2KDhnRSskvdF0KSV
F57EFMgFoo2xCQjFEInKUQyb/YHqb4FiTLgEFRL4ja/El7/sh1nC+gOQ9iUCSQqUr6x+vz/P722R
myw6tMwRRLqtUxPrxwVwawMjjg4Xs17BMIntWB825empKEgBT5eq5Di5DK35w6/3W3/qEa6xDxDO
GYwA39mBaFdblcLnu1H6O3lU/1L04t348DmLW/nnAWRPZBxwvwolVuSyVlNfcWprRmGahqEaHW/6
G/nx69gOMHTnYREVAlTpZnv/pQcOT+ipOqrIEz49/WjG3FYcg0NnmLgt0nvWuDPKW8IABtFcfIIP
5nuRFt4G5uN0FBRH+xClouyOR5gGsBOYCE9knnEcfXia5nIQuX+l00ZcfQElzMkLgnhCeetZpRYM
cNe7E/5HsB1gUdiLKYrma4sgxP1KCvNo8O6d5drQYDlBLOAc30MkEO3F3A9NZ1XMQWhYRFPZteiz
SZh6ZkVPFUJscJjCZUBAArQVShQyd/lQLuIYIv09NcKgJ0ap9/oi6O5gPrNNWtZKWJVRJl1i9c0F
mAOA56iALXrcMQ1ZWzvIJghkZfKjzCnGvIYv1LE0/RXmSc36gQAo+a/R6djsG0Ue/MqwJYhZmLmu
CxIm0DNlRk3gtSCE2AWYjgAUDD42wOevWmmUSdJGjBUaDT2V3JU1eR8Vwp/DDmu96xh/FwFWutd4
PqdHpcVNK/rVdoarP8WgVs86JEpvTHg+QqS/6tTzm6Ns/xxuZbLmZGWXT3RcI5ougqHSm++CkXc8
OuoNH1kszPTl3AHw6UV7E75JYP1DnFjz9e5ThkIQk7SeJ/1eFiWdoFLc2ETpyCLhNLQvepZlB7as
DIL8lho54HmVRH0SQuisAAfN5NPyL/CN2vbi1TKW6nMyHoeGP4JBWlKxkRjhFeMIDx64sYE/+1l7
XZnjpInMLtxLrdhKujj2jYzAx7XDmdNZzmL8w/LmQ5kHqDNjJ4IT0TBH6jXnoz4nDveVr5Vp9r5G
AIajGKbHDl/0YLuEM0VH2yUczwROa7o8ZxYpdnXUrOyGXAiSjESpcnZZ4nMDWXIxTAaB144DBzwE
t4mZixG6ZxWBCZNk17LncYt2z6NY4klXH87PFBhKPFBwCIaSDnjNlXRLNAC/QgQpv7EyUfrbTRmV
2ZcgvQnf9H+XnratblhpuUZ1a9nMN27qB0h5ENshro1gB99//zWO78qSHEb16f0g4uw4MlaNPZgI
kXaYpL+rMGcTtIbKwY6nHsvtVQE6zcREJA1uDvTtwfjBfpyqJ/i4NfewsTqvhrU/Dlp8OULZrF/L
jMioC2jv7ZH9SFK7Rb0rqrGpPZqg62PvzLZ44ZDMavCEnw2qFKQvxIT+UiY57/MUozrICUXcg4Po
ju+xMjq60OjRH6AJ3NWrvqB6V8MMZLGzdLDalF1FZ++uizwLWJMzSU9imeHvVO7lyU2NSLs8Y4Mz
o15YOKhov5nN4mrl/xKSnqK4s5x5K1STMYPkURvMlBGSKXfNpdWCrRBJta58CPmnlfmQ3fXYJaIe
DSaVdUX8+apWeTLDRDPkF/DtnTT1lPP6hMg/YQnOMEvHPLibEm/DjIVndyDe0Wig7zbGtXY8VbIp
wCyGwi2O4gJGGDM1je2DGCnQaOnh4lCNPHVxMIAtXyUM0R+lskm1svEyiDrNGlvdDjaB0DvqrxiB
v8q7mOY1pTVX6fZPv3+uZLEGvVzN858EHprN9zPmaFR8biHg5Gg+Wh0fnJZFwioeYKP2dTqNiE6T
EZeB2DnybdrFPVkEZAh67Y2nFcjRDtHWjsZF81EM0Qon1F73t2SRWtGN7IlLfo6TDtcNjBtq3rsC
8GCORJNIEXiJiJ2UBo0bwJ7WaHtyoI05K+Bel23CzSX1CY+PHoCTe5r5s99Mcg2BCu18NfdxFZrB
+wSW16d7OD8e/mqpwiUjOL54xOsxqlbUFSv/fQKDVkujbhqWJTyhLvCbMjPrvRtlHZR2zRYGo4Ul
A1Kg9QtU3VEU3/wAzWZo1+Z+9bPAlPPbnnpzR66TK7WLu8oycjb4Am0iFcVGeKN8rwQctFAoGPu/
E5Flawk38r/ZzKB8Dw+TotS2uerkU+zbFbKXJ470IvWdcB6InWfTe+uAM6FednsivnneW6vcaT2A
IMOPui8oi8DIfUgI4VAgiIwh5h2Cw6HhxjKAqDch3O52AotkvmhDNnCzBdTbjydvh6TmfKsoLIKQ
wrAO779ZzjEStBqwuDK5g9mT/ovRGjbY5d7iFYsmye2mAq4Ih7ihPPEjRM9TvPOCjxB/CAxkhkX0
D5m9hWDxYylXObH3xgNAIrjODHQr502tvxIkRdiO4Sx+n2THg4WKDvxETZH9aAMVIxVWWcDryRDr
MEJnBT1yjbuNGl1SzVc8kU2NAhamzhfi54D3fUX5E5DiB0WGRkzsV+9WAewyJ5p2ZVwjFQqVYuZW
9YmSVKEmI1oMkXQUhIs+l19iTd5QRFCoReUUBVgFhPWNk9zGdEFJNB1gUGsx1CLSqTitK3NrUKUS
Au1nhg7M4sui7LRAsT6GyAk1WkbCH4qUU63GTa0BwAekaSKsqfrvVZsIM4PaE298utaNYAsyEp6p
Z++MhLNUNlo/LTqL+kWwC+x3dTjDsMnpyp0S0SkoS9mTl++MUq8IfIZOZ7kOAq5XzkIzmfzcV8M9
msurvjn3R/6VeS8/fZq7cVj20r7VeKhmx7xXI7zklxy6IC5DeU3HeCnnd9prklpvKL8COwgrn+vI
SXtM3MgMKSbp3AeDYE/m/BVUOhDwu3LiBG4MLjMKwUVvYrcLRtrZuleB1DEWa8mJI5Vhd8WkMWn0
4/TKygJ6BeVruXmHQ84cps7gJpReH0wAkSfh5DL9HUH0kf1e1ZBN8tgrTZ6MWHUMYGpbLw+cKEpg
9X6ryS0m74rVSTQmUXK3brTkz37MjNi7L/bcm5f5CzBd4U+wReCcDv+/bXKhkK/MDYHz7FkAg1Ak
IeB+Q9JoF111hMUUfjibVLk9eUeo/epHN2AA18rY7ERS46jQbB2mpsyIlgMO0fr9v77e981anXiE
tJSIjIungI9lP97jrEiL78FdLXNJg/qMulS5846J4kiweD1yQhK8nsxcXULs+kEBU79rgkgvbA52
8gS8/2RCO6fklsfIkxalGs467mlY9EoOwsiQf3B3dVj86TlQ3Zy5mgj/LSF7zgyI477c/TwCg68x
ABLeMhg+4szjxdklG/XqdyNKBc56FDFedzDq9jMp8ZhjZibDhb0uFv47kBxkKSJ1pUTdPDiGJ6UH
8I4sueHQQ+XYPqjy6XeE+/aG2PNda2VH+dCj5yBqfo2ATsHUc1Jz2NtCoN9jqx4Vb03iEffB5VQt
0qeStRiQVmbfMbeuWNURDvhEus8DK2+el+mtAWBjjqDrUFYB7ixRPTOFZKlfBVavckNqumJlhFAm
93FgyUSmW6c+x0Merk1b6rpuk29CWoElDI+5o7TbuJ8h0RvdzjXXvnS2HJrzqTrCbDcxYLRw0rPa
Ea7f+P7jSFsnvZBRZ8lV8+5zE6NZxfm8x5x7dEqL3zlsb5tY6Q6Ff10CCv7+xN4mibOZ7A0uNSMk
eXTr1stSqo0PPz9IhIAJ/ChkS3XrU/rZMNk7XeiIIy48sBwzYo+1vyQUAVLVvzifnEG0TfABBP/d
bKE1JmQS6a+N++cvRF6i8hqoBevV30V5NC2QECjg+gd02UypGOJjCtSDlehFsYRUmwaL0RvjkhuK
AU28+5W+a7PQDlGmMY/sRxHziqxAcaRw5arIburpY9KA/Xqzx7V/4ZNjKtFo8HY7zeKt5jV6xS1a
OB7+ppMAYVfDx8/GYLi4TdCPYQlh1/UEKQh5J/Pc9sH2cCBJNff5rn6BjIs63i0u7OXbfXYkol2A
dQLNhSh8reRurtdVhZjdkXTHP6JlJIi4Sua9+tNBIj1EJKlY/MQORWrOSe983vAOVFtT0gwbE52X
MXsCNr1ddfEIh4vjOFBXsQ3s63yyR6cnzYERlO/x+33x94/lAw5Sjs1oE7d2GfVHV0BaIw3bCLvp
jMSSBqUisNpTMlrZ9eK7/VufU6JCjxjQ8YY+SO86z8ZmTwzAfFHevKsc/UY0EuJTYrx+OBieaDh0
8Dn3yqlzhvgef2QhVzvaNTNJWo8dVmc7rSQ0upFnQcv8E2B1eaN0kYrPPsScBvP3WyXadP9vq5K0
+7ljj+YfBWmBxqJXQFAhLivPPovJtiZwY8KP3o7GRe3bsgr/rS0w3GgOIAEEuk/E/rAGYuFYgq5i
v9cRINEyt2MlnZ/GVrZD+XbakT9qhj6uWBSUOgucDPIImA5KN1xCv7dp25ZGJtwy34oJD/TzKWPt
kVCunmI3i8R1pDMJodpBGZjd7CtpnEaWKcZ2az369Er7wQqii7bHdBE+GZQDlLjWMU5ASyn43pnM
4LyQLAVP0vlQ5IGgm1f7cUqWNBaWIg4Ixb8ndMBPpEKOdj32OcS8CD65Y1IE30SOnsQt7nWCkBnm
79tM69QOtlJ+L/Ht7hQZ95cPCGfZDs0kzK4yRpex6ekorfb9VR1MMtertPK523IYGhpYPaPPilFs
JIwSMCqcVVt7gV9Wm2qSwoivj52vehzHPvQxKqSPg1kqnGY0Uw7zjTuBwiAQZ+7pMtWjx6w/4aLw
sdhqgD6hQZyh3q1Pl6nseUbP2WC23YtAwa5B7jh5qrLpjtdLS3Q2p8B5laxmJZRVpc6Su3mT2sGT
JFsGOGRq0bN6eNuK1g7vq50CCNv3KLvxY2hwaJMiMNqUU468QM3xv9SOhBIHwbhz81nL07WiR4tl
Fr5MClltt1P7/3bOT0O3tsO15tOqWSl7h4n7yz8TYs1B82JKEwLY4Odjsp5Bx9wxpj1BoQ31OZ2l
MXMkzT7PXYxZsDJpJSEokdgsWiuUBn3c7pJ88oiEbC+zNA8AOqNHwmKGEHDaQHwNoNCft4m3Bd0M
aDZvhW8eKn7JhhxP1YKyKz81DVbxJuUZ2PyvFHzw5Nyi5j8bB0thZmhDhcS62WgnA4HnKcQyd+0S
BdlcZvzwy/lODU/5eYepDz8w2j0w81wD+rjsvR29jOBmYPgijfCYZ6bO9ryQIgLsRrlqHx9W0R5g
O52AhHfF/vxQq1wGP3+YSsFAfadrap8tSAZVfY0VCSsRInYJdvgBvJjh/+epjTkqRbjTsLvlcbc5
fyLBbiQC4/bV0QdV1npzpn0gokY0ggvhlBoZp9MrJAx4hncwCntCQzC/KZwuGm3uVCQwa4dW8fGk
y/k3CTKhq0eWb3i1FDrgARnM5omfQxxgBtOgBOpADxS+Qu4TYLmx9/GQWt/PJ8BI/IynA02KB1yK
kCsAslYwJEPza2wIPVmfXFyGt5LyR7zKjVqzFGL20nc9SBPvGabBTdD+gZ8dbPaQTH9HXKj4ZuWn
ueXWCfHENYhlIhOEKngs6N9TTG8rhfRivq72cq3MX28FwOeVY1YLEvvoNhAbyqiAwB44LMCv8NPI
NDmIEzylbsNUuNa63TsKAsrhXndpuIVvQrNAeNC6wNSM1308px7Rgx3e/0cvlBTSg9SRgzRQInwh
gFD91UEHg+PZ3Zk5jpHh2T/UXEXlRRhic3iCfUGGmu73eSx34tgXEcptx8Ol6Hvcrz9szpqI8hBw
fBa/eRXtjKOZf8sOfx0+XVguzo25cJQugL1wkW2hxr/qW++aDeK40cUi4slR9DPGO2VHc4JJetcj
xcP2X+63dIrh/Tn+z9t4Beit1te1qJTp7huf5evrmBi2Iuba/73vL/wcyE5tD/5EuXTC+5jKrh47
8Mlavlnrd3TB1A0nDNYgP6fFzBuTEiNoAo6usc/Sdq5bPWzbTHINxPZuMCaSR+xXlhaTYQC06a53
RrcYqgz4MYXVR8ZMKmS/Wg4nvmJDgJ22sALAnHWXmlrKwRluyTdToe0jkgoKvP19UffwZ8ZNYKhe
gKn/Kz/s9pDuM24rlXTGTpBhGSEle7/yhH6voPIaNXTMaowTsD9UzqQFZhNczK4KXB0GI/MdnrgV
aIZfCJdh3wxl38OLibR2GmboiV2drQp5Hmi+CYogD1WqBeh/4T/Et5QEJ/9cXoz3/EWYdZW3ez7B
FxJiySaDy4oXhkuD+YhILAhDtkuYtjIR6pf4Q4PxzH5E13hF9A6RYxuRBR4wG6tTH3ixI6/e6y6H
g6wb/HPnT1fMztqAW2dfDx2pVSGwAZBIr2ajpzNshFqWIokuJd1YsYMRcYCRcme9lSRtGzl0AU8N
6E1QuxOhpXhNKDaGpMhDqpSWNzmgdCe+eessXf7piIxESuO2TACjH8XE6GaAs5E/VBDi2CzHXgTU
PqgTm/BT6oE0gVwRpp31PpfJ3oBd7UAsxJAS1+hXRjx0srJHWNd3amdUsRII/XPoEDQ+NpI/ZG35
tx3/qpDghErZKDOxQ2VqzJLeYz5g32a1wGI+TPm5DHPxRMj7guQ8aR2EULAg5fbNVui1BPBfKp1+
z8G0QxkgWPz6Bo3H6MHCBFNLTkl4iDvq9ue2NWFFbYzFhKfvbNP5TJcKSIfleEyD+78GB0VEIHrX
TqGEpO8AV2hu65DuEXae0ds5Z6BvXHGfyIHoC2NY2fwY+p+rFoHzU2a5L/7N2rEzx01sXAr/YHPr
XfUqBmp1ePGwZ2mOp3XXBlogULsiOlB3bNln1ADQ4mMgRlcoOK9Zei0qEV1DzVuXGzC0inUOO/lL
ffbj/VRUJzZXMVA5OYcKzyvXb/Ms1SY+iwWQ69qqEQTyf2WNV4WzXI0PWSiArRuaDF/g/k5ZN/ti
mcrdNPYRaP8aw3PiZGhgWK0nzLYalH84HBozp9cPr/Id16c8/JMeSw7OiEtbbLZ+9V7Ppq3/psm1
pKdwHx/UW4DazBuNcC/cA9S10ZytOrku3X1bH4R4S58VtJojshPD5FS4PccEMXFkX+CKKGd9cOWl
r48J1sgGxF0KCVxydCUeVdmPnoTnerE/32MlXIu1jpsGM4Va4C82ysWOf+9GUEuLgShf23NZ/Two
RG8RccVDN3O+yNAvI8nmafrw7D8Szb+U/Yg/zQYSNItOu+qVeSeSCBozAKqqZZgzStXsn/APxrDb
NiAMN5MK2cMW3f+ZS/4TgKENq5t3mp4IE0yp/QB27+tFtgJsIpjkI1lDgpqNRVFbq8HkaIKRuquP
Rc55VWj/xhmOC/03YuOOXg7699zR3ckLX2rAwoP0JZyeRSPBjfGd5BndTMbkWLicCI98Qxj4se0y
72ppLUQ+1P1AhgRaKu5wAhFyXzgZuuT27NNan8NsisVwbAGkbVrgGFiVEHYVdfI3T9sFtvna6/xb
sPRF7RemxTx06X5hZ09CK3iAuRux4A0aWAQ6X5bNoZ7pZXd6CfHbv2MmB7lyjFvdPAZyuEOP+mL/
UgCDc9Q0v5W4h2D6HU0keCuqE4h+DB1KH52lFaOk9kF+ASPrUi/qUjmF50b4byBQL7gBXeG46GSG
CWbyY3nnGENYlL3sio7IKNY/TQzRs4ejt94QdEedJVh+73FS08xVIfxQ/hBRZdgPijy1dhphHNam
RhJzzDIjryYDsrB+exm5r+8n94xat4vjfiiu5ENB5bI/pwAqN1np+YraoHE34clsHwBQKg+tqdnD
TjcwyMN18g628/YJSADW2Uz7H9XrdpMebpmlO4HPhM2Dfq/SaQIMxui3RyYcyzYiCyU/df7rY6pv
QcG8/vraL644c0Sx/JK04EcfLoXvwllAsM3Go2zMpok5AFg67Pt8dvCfINBP0R2cob8L3+WzIbyO
g67nywByWTgbiWjop5vIlLNwyBjyMlh8i5nEXDBDPr6ODYJXdF9NKj7Oc9El3hpAVn7E+WZ9MXgP
Mrz46LXvfxxdBQ9wlXEcdSXvn0Z0LDEV+4SWl+rs92e23oEPsOQWKtq5ejLqCpVlHWLs5aCoeW9o
3dWYhOoQy4ZGP3glP5adzq77RSA3rJE4UgGFWkFn1iJ4IrmycqvfK++9Nm3VU7NK/ewWbFdh2WUL
zK8/WYvwtY4ebcEC5Dhlw/bz+nZ8vLol/wLKsrjzvYuOVglH9YTDF7ym9BxbuUmZaZ1BKn//DYyf
MIm9De7xa+Yod3usXdEzS4e9ZGrhc9UgD1rNgV+ibhwZHrqSwzWmRPMJK8+Ckqw8LmvWO/E3OOgz
3onV08u4/qp5uJ4Md946qXSkP6MQc5HF5n5+rkxQuPDHAr382cQ5bIfRZ8CzuIrNejD/s3y9InbV
FJAeoxM5epRuoE7XnYQzQNHaz2jePAiz1RN69+HbUyP4Ji1+yMMvcykDxjWYEJSXQJqQqVDwQJo+
Y4nC2DGlpI8aP+4zqigLL+mawnuxv2x0So6z5UzG0TYHPHF7cggG6J8nMS7N6IpIrPHhptOCmX2B
j+mB6Wjayynik+cKCmhlaTDB2mO1YigYh1Kb59tA8h1+Es6rYWQ9967OKpWS1kB/fAf5dp5NMHHy
PEA6ARQEVFAgY9irzM34ExXBmgsjmVnRroUpcaNHUFJX03TfaDHQk4M9WsBbNUMXkbS9zcDWDe6/
hJngo4Dya+YbUWB8uVv16NjV06XpLBkSriqmQRd8kvoYDBfX6t5d2o81Ec6KaGzw63zhwapo+xVh
X7X6Qt/DikqWRvmlsSaU8/PcJp4DLDdY18b9tRayQu1AWvVR1tlOmll1aVSQcQCKo9uCoJj+4vbN
Z8VL1HVz866zCvAXaD3C9S2ufWIes5GoF0+k7IhRKlShvwArYDvRQKznWAfd9H6IkAvxmXUyi4Dz
AVU2Ei0FNxRrzjX7PnOjnnx1QuEo2Ua8SrjNw3g2kE6RFIc7otuioyvO7Q40UL562BV8t117cF6H
+iFm8aSW0tiFTRUvsIt8c2LPEzxVX6vIykJxC0CPJW8Q1h/bK6kECtgraqwc8sSLjd/RB371lH7p
7v/ujEMWksKHbj5WMwmjjJnM31miO2Xx+VBAAjtkzGwurY2+81NEbi9d8mqbBRp/F39S17ygjRlP
9mCbWYt4Zg/y+16E6eMk0iu12UGIsNspAJbevzpPacPvtEyndYsaWTz5JBvHOQYwJDiy3uWKkH6T
Sv73WkOVEtyP8WHUB+ILdGpBM4hhMv7vttg/Qtx/3UAQ07MOdyycZxT3nAhVrEBZGb8zUXTWAzGX
4pHXhyJYX9BSuDHlYl9LAnBiLXzZFEFLK0W7vfAlFv3/11vygSA9oLi4dwDhl/9WQnnAmtKGWFEE
HpZ6mnYGIO+flCBssz4BomsTc0MgZVVpdMfvoqMB5vylSwhH73oyR6w0o7uNimVBBykTlixYYu/9
jL3eibSAZfDqN6bthfWH8XgJ/ShNI+xDYcJo5WvzybCN1fwcUO5Zgx8nW9yNTe96QROwNEg/F/26
3huwUVf7DX358+mA29z3BiSnM2cjJjEQJOuFAj5qBIzWArmFbU/fIZ3OcRwQ0+ap5wA+ZevYo6iW
28gPjAFAMb11AKMYGeOMF1dkBEtMjYwhx6/6o7RE3GeWrv9C4PAKGlgncztxMRxhMHl4wt5y0mtR
5y/mG/AOLXyycUzapnx00px7753d0MSw8QbVggGI9NYgipkf3Ric9y4fhPNKA4vg+i37zd39p7JP
hX7gm07w5/r/G279lhmPRNuw63J7anF8ZpbfvfbCel5SF6Op6fs6gALA9rePNRfn9fNyOGOP+XL4
V58sadj7uwg+o0umu41OIAAxRsTvB1dDGh3D8rmt9Vvmk73PpuGoqwZYOkrugDpCBbIlqVNWaB4Y
swWoOHdHyWqqTDUS38Cwfprw4Q9TATkiaR6gFGJzKScUntfa+Onev0bUgNAk78EafALHsZzoLdER
oXD2xYaJR8NvL1NhqPvCCjBvscPB2ZlW+FkxzJaDUSBxBxtnbdBVw6leVlGoHeNGsItaYnCNk7tw
Y1HpspqmQEcIbKq9vqZXwJkO3W8zGbw8QUp2gDcmneEvBYCvBWGrRfGXWHWqxvomS4m/YNhFzfQH
PWFb7tYP2Ik/pg6EnSgn/zu5Q6q6fFPFhaIZIG/W9kl0Ar0Hc4k7sA7XKvYFIkeYLrVjbzIBvAQ+
V1Z+vDU9H29Xi50Ngp+aQYkzCEns4j2DB9U6GoAe2udPFV7TCkkQLe2KsLgw1EsMAbbFn5+S87oN
Wv+t6UAyMiiZAQP7gPIROHXXO8f9ej/zFp1wN1AoLlZ44ULKlL7SAbs1sPVnQrjqXWquB0MPZ/dY
mRPfOynxPVcGQ4AGEgsDOb4lNbzY7gXXo3FQ69uR5XwvIG6N34zXF2HcIhHwdXwWqs3+bdw1L4qd
oKo7k4jw0xegxAcByC0NyO1AymkrmigI5Tuu/rNxuSOURS/7CxWXNRnezJU2fmH1hBczjiCdIIJM
JLP8w6eehcuwdmS4lC3lE/IQObtIKjzvKg+fiEG/n5zpwTlT/qRzWkvW2ey+uJxjazf3mf6JqzIV
C/5iw9Nut9KyWZWRu1fNXbu3hwF4Zk+WEh2Bf2nhfhd8zdjjzPMcOvNKBySuoljZ5qjLqv6gA/Ya
NKnxNyylHWFRqR0zTBkSclSPRyF1A/6IfNff+cwnsXlud6Cn/S3RrhfNHW4dOlRQjO972akkiB26
lsQQ4NMFuxYQTPycLv9GMFLpbgmIx2JsnHXonwP4S84/9MYiezC8NDax0Rh87tMB2RySmZg0wPUg
H2z1DCdKgR4o4Lb3w57ZVVYNkCIMdWEy+l9DD7ksg/qg4OwlC/eM1ZigF7Og7grgjzOTniE+gAQ9
ijvFx1FcL7akfOex1JFOHlrpKRIph91Apf5Y7BprNbnPfyVXRNPA27PrQAsp0Q2eLSULeAejAq3k
/3ba9JQt9AX/LPbcWi9eSQAGZMy6pArOluJCQmUnPpD3/LXGmb3PHObX46KtUu6bi3TJqSjiq+eX
m1Qspg1v2wJvjfMCrKdhv1V8Gmzl48eRzHLGEFkeHXa/LCfgVb3NOS4w3kwrxRcTqUx1bGQEqMqX
kXMkmjQFRXZchTJdU8kt8Uzw5aNwofA81YsAA5qhJO5djryZ+2ahbaM1MUPRm2bGZyQkKCbh+iFf
WUXX6ODxMaWLS9UOoOexkOJ1Du0bh1ty5Ovum02mCnKgcPAnWpRjsKwrB+6G3Igd98StqFWrKxAN
R5hzWeEI9hHrWTjFCiIy+K6fZ28gvL9kI8rxQBiMUJ5Er6Qq1vK3jIMzRpfj1XOoVTkh4EW+joU7
uUDgghH8eZnP7ZpMniYaThDlxDfTuZ467yb1fZNZfqLPfN/dWnRh8z5L3Fy0CPdLOmSwiehDWPTI
MP/RDz31DntBQYmwuXLHsCYnMcthza5aE4n6KOvKZ5LYd9R3xbtj+utEFIvlxuE3KwxjCvP069XU
srAa+/Q5eUcm7PUQWbjEPUSBhS2sq2jxWidgOqjBd1MlLL0pmnvxhkWAFXbH1f66KTLEvkG91zCe
IaL0ZV38U96qw12OM6ACkeXr0Ys5jk2eOJeb7s8LXTywd492Wf1GMBakljxTOrk5howj+62oPsiN
IBVVjiXV9lxPM5Zjlm0dzOhAf2L0RCcgS22P0S/DXGlKvHDPASRaK14tfIYFFm/LHuC56wa1yMrg
hBAqcAtKlBrofAnoUrBbm2Ym3nya7whqSMZEJIvYP0qTvKmoXMv4sCH6FdSHH8qP0Atd7fM0wIjo
oqRScSgA2o0Ku7yJy/k8BsStiYpzJ2KfSSGBxFJFORqSLtxeYFsD+rByoHcBZhwASwrQMwGWYsmA
uwDkE9NXpfSurFGb+tqimlKRRZN0xWI5XYge9HawwRWatJtVd9fOT3u7tZUNCtI6y1BugL4xOqiy
im0R6AmAFpnqZlBJws0Q6Gvv4L3/Spy5KHzMtXcZqCgIcjlMhoreMFKLB7No0ZqfE1pow0R5NxK5
J71yv6DkQzr8RG0wQkaXoiMauOjSgjM/RCadSt1ufLscucMASYBhXiuUZXcqVMxkCBN4ANTu4wXi
g5RHWgBpX1xFmjY4sFBxHVRtulDoAgJrxQZvzwf+W1gieyax1m900jOBkegjiaE114XDMoDclaNU
zzpH55KcI2TGE4Dbcjk7ErSgXmyYYvq+6MGNH4h9lSABM/brrFD80cfAMiwAjVxBmcCPgda4Vkga
g9cKqzAj413V+EZ+8DJhu3zr62ziNT/BqYM4S1GNy0gypQeXFR5QJo7vV/AYMI8q56xBelJdGejI
G6KrUBRM1Eq02chF7yN4uUbyDfgXrSvRcycqRYXX3F2mzaxwjW4MuBxwnaVDXomIL/NfqzO6mJl+
sQnpUAmdz3f82wTn1EHHa/5jrdI0qkQ9wVdUWM4yYV9xmoir34GQ5ymyHCoq8fgOTg7R4+DanPQ1
9RoaVx5bjeY2Z+9SNmjCk28fY9abqoFykT938xx3mgKp4OediemIBQ/HUoTWIAhlHOMues1IiEnI
2qUSoNgeIkIVWKywUu8Tnb38yG+0iqKnTXMcFfqRtmIywA6RkkVuzouSfw8klpr6IFRMSyrhFarg
40q6miYsW409j6zdKB6lMiKeOiTC1TbC1MpmHupVmz+aKMzQ7Z3doMAkhLaBSOiP+GqSwbT3j4+6
zvW0vAQPcoYnk+80UKeEeGf+bJTGC8XWD2fSs0hRNCoif6KQ7pzm7IWxXjdXJdPHGUo+dd71sBfj
Y8oRChT9r4mAPEuFdIYpreK1ZGwyVi1uxhjI8LYs2DBdb/3aNw1SWwDmYEI3LunxkHDGoIn+WNSA
oXu5+CwmH7e2pFqgCClBdhzQnaUk9zOZfdvbqeiFxnpPOu+wbJ49nmFdWgtxK0RC8m2I/CmPcGNM
77eC3VOAzjO7zg27ljazFriRXwO9fXYzoWizVnf7vD7KpMmW9MXoHCzVxUvwIiPFbNf0fyvXpCuh
VP0gGndxZvbEr4gPrxlFJFoCCqlsIikWCEFcauMkPyxc/DY3kFQfVK2DhPUiPNfLOc2/fPfx4ajT
vHOa94uYsOLv9bcDcioqzQGP99kN6C6lrtKjpmY58+KBwd/F7a4XcRTytoDGdZPk0hLnCQl4lCcI
VnqKdMvAHc4sNNx8PgTH5w62oA8Eh+nKT40L2VmErKiC0A765FNQWpu3AhDwejLPGcpgPeAJrYp+
QWWlHVeiO0UvSTFIrxcW1eJuShrxWNS+4xRP3k3VkJDtWhzQ3uKXBfUpSs6bsg5UdBnXVqnp7KSo
f2LPhkrMAZhTcginPEdkW/A1PBmlTkHnnBFeD+0HjX7zSUnp1PATEx0B0QsbURJKx+lN3wm8v5OP
x3VxvQ9EBExxZlyrpfL4mNqnq06LlZs/rwv0PCgjSckx1nUt0BCwgAkVH0I06fib6M5cyRTlhAnr
gGT9JluQJ46r+1VzyRPe/BLbxmLxODjtFCQM20gjECFDXfVLde8J3KL32p2UGVsugPpiNRRFUffE
npccipLsHPgx8p51BVPA/fsCsmnOPd6nK6mv/Gr7gqVo7EWDDSE4XE8CxIBNRYanzAlQAf/BYZSY
WhZoexbHdZHw1a9glAJ+NMJcvsD/J3OUaiOgBT9pxibOt74pwFEs11LJ8JqoM/6acnmOvVkKqnCk
sK5RNPBzR9eBqupLRZYblbSrWGUeZQJki7nfxQpo59vFBrr2R6JvCGkvRY9FOvhVM4LqTlIkszEi
JRv9VSOWt+QqY793fBsqIBec4ZUtIU18fO6ThvDMrXY+Q/SiaOIpRIDXBYvP0LWvRZK+V6frSTYE
pQwR0GHrdl8sx0Rp62C/5l3b9o/2MXcaB8yuEfDP0rl2f7K3TAp0UGHMfwR+0vWSa/E6FYnopiLR
R/iALlhODc/StMS7MN8c/4zxTmWhmrYOXnsbkurClytVMyr+vlEYRJOYTuYUIy6U0gGU/wycn6+x
Marx64U6zcTt9vtm/UzAokmoKnAyNUFdiPDB8DYM4Sh6qu9KQJgPmp5egP14rJ+nIDReKVnT8WGU
3JeS2wRhlsS5+hHOK1uVg6VljI2Q3HJJs3IN9xpV8mOUvaUpXtPw+hg9CAjIS6Lt1z9ump/piHI8
ijj7kapyICGNGOxOXOBYxJ2VkrAQYrrWXnlUdh+CJ6J0dEvURiYOBDrLITyuFXDnX8vM61jttFiu
uZQLgP4PVi0bxmqfgPU0S4THWi2IzrNWrBR77Qz62wU/rZEgZ3nFGviU96RiurjWJstdsT2sBuuy
KVlyjYJOXeS/Y4XgF27sJzs3tEUTL+r2LkeVGNuBD5ABbC0VMecnZKT0TBvUS/lkCVcvQ4DxIGgO
xVhm9LfkDXfVvM4vyFsmeK7EcTCXOLvZLYpUfHoLDsq1SOZoV+iRITXTfDWku986hfUz0CaUdg72
Kf3PVN5mOMUGu/AT/0aD+q1FtfVpHtv2o4nfO1wkgST/NXuyTBQovZB2rcYLu2JwsdYTPwHDLbTk
+YKFEGeH/XkMsY1tDMyKBpxzKWtFtoSVVeXBkvpYz+SHJ/aen57esuzOvXmfRwv3QHZB+oTxkK5e
nJyN2MNoE6B/iFB0M+ubEVIBuQZLadIxl/iyOuyHJHV2tDYeJHqVGeQXP95d3ZRpjQWS3JZ0yK+U
DDGJH70mTymzKhVza84pJ9jyiyb3uVpr/gRwIBtZQ2k49bWohnEi0M5Pecp7La37yb26jQoNbFci
YfhvHLmjEElrvo5nAJq+Ifgdr3/Y8LBkXT+Lak/eIbJrvwfjYiYaes1BliyTP5NZk4fENrYD155D
nUQGPJqJ0M26VsnEos3dVw5Rw5FkTPacnQikMgdeOfBvLQToYHEW1DE6Te8y4BYlnbfNd6W06wSV
wkbIIBZ5DPaKQ+nPGyz9blsxXXttsXb7fldRVDp0rVwqO1I3IuQnUFvuQ9p/a5y7g7/negilLRAB
5RxYM7+Y8+E2EYUnEdUDet06qy+OF7Dtq8dITnY0YQ9Sz+m62ga+KcrFHWmyDaiRTXeUqtClIM1D
37yQTIt9XlkShIZGY5qsUPKgk6Ht3ORYUlWtGxsk1e2r6eoGs1LiYRZm7Ajo9CNncFNMK4Eiv5GA
DoGcPQLzbrDyLmrM2f5fBQcOCUvO64b7Zcx1KSE/S9gJmT3VcLZmO07D0N2kaJvdNMbjwCyvAk0+
5AS3OSF1oYEck50WMJrJho9UcDyADVYt5YZh2KGJDicYUba4ar554TlsHptAlEMUglZvfNTE+qeL
7SNX3ed3VtoAq5HndQgVpiE4aus/asyqHXCoYNlv9ufJU2JYBFYFk7oQk5h+zDSTOMPcHFFGWdPm
ifPY7f5kfUHgyC7OjYKf8AAPkkZIGa2gzODgj2IN9875bfepdnzp6OLDDRpnLEFyXpshqmBvTOyE
rAolAIbgZVusMvIfOrFXMdDuD16AfghFgEzVk0QVGVcimhp/u+lZRnR2HiZ6nhFqw9WKjeG0gSr0
eZOHA9njCFkXpgp/Fh/W83JQVxx6VONxS9JF2cIH4hdIp2u4IOPAYM6Drv6XzOlT4lXweV3VdlMS
NonyMHXIeFAhvkSD4eUBV+FR0/fry/hkb+QVaq7rOdvHvIT2OVE2v0noB06AXMxJlk9Qdudi/e+H
paECoKfETa2ylvyoJokesedynDyaErtooDuur7RTGoldZJ6vxsUyapeHnNy8Faj9XMYtzTZCkpBl
MZJeQpOESjnEeK/rxQyiSmk+lunU1s223jyoNN32PoKZCoHMVoe7WdAx2dYpC5K/nfA+Ad5nXW5x
TpLfKsBhxJIZECx/N/jHPi4ZfrpTNBZsl3E26HzldyVzaHqrBvKFFg0j6YQ7+JPxcKw0iDl7OUjn
+cfBY4ZuhZZBeibB3ikGFixVY3Zfm2+LdLrvvDTdReolLYDQ339aqofT+5r6wCtu4bZ9aYO5Nzuu
nitW43+74C9coK3Hu5HoAjyhxeaCltosjDizXP6rVbWp+4pv1cG5WTMc/P15ToHy5L5ip0en9apS
o8LIiXIHQLyt5fDwV3OURB69ZsyGPVnpt2Ve1tf8ENufX9AH1nB6hEr2xZuKhhKXaItoHF1vO0wG
1yfZMJovdz44zoANCYQjr+5FOeGeoaOW98IwH6b8B9WxfOTLDPvNrLl7t5AK+CKPJ9RETxJ7zvA6
aKsO71r1R2wubC1V22QI0h79UWhch51OF9B9DJ374Try9CJ5R32SpGF8zj5rAvz0v4o8hneAgR8B
sODakoVapUMAIABaDTg7nJjhZiF61MX0zTctRuLYAOqbJcnMbdRm+/+YXnTcYF+4NWJ1iiw7uqSK
ww3SpxRXMM8sl+fqK9cL0MHtmted5aWP8ymEIMB8WYMUHeek0ao6dU90ssdeSqpyZmjAY3vX/03H
KkVaHrTzgcw45N3QaSPBt5IqjAXopMk/pDhxb5/Bq+tIjoOCB8dVXE53xL/Kh675qxuMkrnn3rch
mXylt1Te4iHJ579QEq1288RTXw8KlaWo/sEustTOvLmkGl6P2Nmvu8XJHbJHqA5LVWalaoTGYy8h
DppbT60Mnx4Vy8Pgef7LKeFtlwE3oN+IXJZ6z/J8lZ+cpjXuxbLkePogIkLEDmi03fAyap0f25T1
Nm/xylMhQMXHfcNl0V/SpupS/M0kTSu0klzMIpHgbnSF24R/CPMEaldkka5vaAXLjjyqY50Tzk5a
71UOYo9ZHL1c3r1wSlTbw9X5oTUyq9dGP7C6f2IAQH47eHvIo6AaWWxTDlaJODf/XKEJLohqvy/v
/iF5Rfor7oExznH4DWZ0h52ItIGaiSOtH3kXnMViOvfXnKE5rWe4dv/XKClj2TlfadMr5TZwemTA
JNIwnkIwac6CeKsyo1QErvYz4pZuA2tWNNnHDk9dYZfMMMVWmRHvYQxj88fwHEVql6+v1DwAgbm0
RdYtslWL5Cp+97vqG7lg0V8qVO2pkE1xbRdEmwagTOgL9VU1O8uRORxdhmgXZr8lJSe5ifwdDIkV
FxwDjPQmYEJX0eC5rfDMzcS7/6I//ltH9LHTt8uO/0/KjbYEJl95BzPaV21OF5pviPtKW1hrJY4v
jHAhHBPFTpEK23V0XHggyKxq0NNQcX9riKebjH2JG4+ZiV0wOZaumC5Z2d8EctZ+vY3S5MRD/uKl
+LfkByP3uT8qW6y+P4M7JVoa3q0aXYaLEYaORR59xb+jW3wK+ZiS75n/Hwm8hQ5K6QHyBpVge6qc
NJKcXJLRRCu2pYGTYcAqrMUcTEo+8iA6KZQRPYE2XQQda2vvnJkGXKa7MkiMbPr4oXyiIIYoOP4Z
GnyTLyYRKUt73b5dBIpo82466l6FS5F/pTpUiD3xKNu8mvkrowWZbhL9LWaDzoNp4Ht8K0B8lSxW
9YSS7HP9jjikM4qy0bJAZGFVn3H3UjTkB9s7RnQHgDhJ+bUYWvvAPMs285HRd8IpckrqTtKmJvGg
dKO4thTHr8X4D7lsvk9PgLcDGuYUiebe7oeyA83UGj0qori6a7KU/hTyX0xZ9kK1BTGF/OCq2lik
pF7EPCGL8hlVW+sFwMtxniI7s58kQlErCLgoPmN6xII/RSBNSz2TGvznq0BWvqSIK2P0tv3pQ55d
I3iuuvhoq9hZKN53iTqpwvzFXaSWOguOXgAYRYcjPVk4jPAYpAta7R20QZd3vioTZ2yUXINm59cr
YdLktBqak1PSZwnUvICj1or34ccaVXWkLDk1YVwoLubzNiOibiacCi59h32S3t+RNmWbSu5aTrKm
eDNXnSeRNO/DnAdoRTuEV/MIr3JiDlyXD+EbB+KdXa7C+okvEDWCB6aNNrnrT69LVb/1ST1dApln
Iqa4zo6aKHhTRCucyFyuLNFsvGdoBfDD9t5ua7DKCLPJC53ZpP7AsvgZluEdfOM/xaLie/GmL0PC
IkLC4vCbSkzzY75k4NqgR1UPav3qWs8QvDDccdkhg7V1H9bv+KKMa7PJuHROOR44caGazRA6ZKRC
lAKQ1pGDgmEqyLCS4rE431q/nggT5katwzIBFBCa6wE8lr96u23CGmWni3uF0u/Ey/hiKn+WrjtE
OyBa4CSIMROzSwc2Rf5rZvE4BN1fmRI+W70S0/ryKqpN2nK1aF2xCq+Ch3D98m7zj8Qe+lTRB9av
7SrBvUDRrgF6CCBQuaYYt8uVnSoeGnO3R8ain/G7Df+gHPKtDseQ4/eAzUeQkPnDvwQDnMjLR8+L
bvxyBEp4kUVSK1/xXw17SEK0aTiWrVpTv9wws1LP43pORfaIeJl7dnTKFEwdGhTzUSdJojiNhzAw
j3dw8KA6TgKizqok3QihU91L7E7R3wigTb/kU5V/th87JmgWBuKUlL8X2EA3DVWppC3PJhzGJ+Oh
+u7xAsPPPguoP4aXppiAE2L8eloM9FBEVrNOkp7DcPqKLKNmaH9EB+qu2TRRBa9m6FhHjhImudcP
NUCM0HJUu28r+D2DO1o9oBpjJ9OLcb7SRtAh6DSPlLsHmgxSosCiSxm84IUBuM+WWUaukGsqpEsk
7w4gGW6wvlJtgVMlvfJkp16GiinBdHZQ491dY6Zu8yhoRQcvcvTQ/t1Bnzl/tjy3VrMrDAz5/uKN
RRnNoh/V9bTHczOu0oiotXo54JcisupN8c9qsMOJbGQZGYtF8HqvXMbjLtElv/QENd8dQ7oQ2VJ/
yp/iL0SiG579RrbOCwY10053+dsf3Ncwr0WgB6PEjI3sZJzGeNtRtH8sNboFwvHxVKhia+/I64gN
SpU5ns1MwW5rpuuaXVHRf+GPPI2+gZHZT1PGDS8ileN0TEBoKhnGoSlDDjmzk5Jj/d7wgYnNWkd0
jF55YBb2PYaqkuQ4Ob39uWi28Q2lMkEQa93NQNiaE6vIz0unYrNl1+i82nLGqkM/BfxOBzneHqAh
L78J7ElAGNcZs07bIH8+8XDFSzOxnoLynQnllHTv29WdxxzscHiwgxS6QVJgfc6FER4zpWTU1tkp
sLO02LMGzPDW9hPZLmT2/X4yZIFjVCKP3hZI+PiW2/DVzJBWm5DGJx/7eWQCp/BIW24G4hGyrmGC
ZiLnWwjPlkcWAd4C80tH2sjlwYszPXhzooxglpWVmU3BKEJVzthZh0uDRYHyKsCspZc0qkmxn8Wl
eg8BqlE557PXym3mjYN7BCqxyndswP6r+zZQnpipxzE9GvMlRYIw6Wr+ZvQi51QyECEKYfNkKfRt
B4+WQqi/d/0jIhAd6nCMo4r9ypYtESGV38y+M8LVrYpWoJ0KwnNwoIzKZC1Nrj05eQRt4qzTgFyY
vUDoXX4THB6KrCrd+DjxtUl8fSPesjXZkl1sF5zSoCGdYQ6JIyKfPMgbSXqAhsS47Re5/XiQpN5K
l+c8A3tIfCXfeDvJfNpY3sY8NOv1NBLwcuJVyKCenuMJNu0K18fOw+YCVFK+qsotL0vqeGB9e1Hq
eRfMktDg1RWUaXpA5r09sLwAZ0OfHYCagNkXwHAk8MJD4Qg/9wt5zKOjBJLP3KnP8d4RBSp7Y82X
UuzkkddCKkO4ccjKNlCUwqyZMazwreuYDuHFgLmfO/bN514okAP2yveXvjI0LVX4XymxsMUBaQsX
z95DegHw9bftVg2HmfRBojGEO9tgBpislntlrPG1U9MmwOL4Yf9T1XKosSXvkqH+Vg9fgI2p/WKN
wRz2Fr2n1/yvpIRcHC6icG5D1aChNQ14mn+xGn9I7U6RflbScwFbG87N7OtjYH7WQT63TfuxPEuJ
0l1HThP1sxaM9OJnTTTNr7JigWNPxuW45qj81PvPfdUAJXL6qoGC81G5GCra3RO2826VPjCxd9cj
JjwVlCz6MZglJuDnDw949/fxwQGmW7U/0RKJg7xeSgz1HQ7bSDB/DG8+RwN7c7pxwRANpj5K7pp8
3+Rzv4i0/2D4s7Byhr/dyvSOkH/Q8FI1Prv8A9JqxXGKwjlvkrQ9pY4AIxFLf3Rkra1blCVyk63J
yUp+aRggJFon/ocs4+XNCM8ZQOpYKn4t2DC9Q/Bp54TAskCQIAJRNvnXdltSaXU4BUEFN1wGsdrv
9JQhXFy67rSQBRaJn8avWblFHyCZQzA4K5iXGmMrP3sDC6tmwnv6cc0g2jmn7PamKjofBIGO19vA
w6f2BpeahLjDxAJER2RxoVS9zdYlrzmAjx6/gOoZsVrDHVRR8lR31ortm0uC1FmUQvFC1kCVityt
GpLV79dddoDG24SoL7+NUZ2BDkCj/aPUJWEI+LrYAADhLo9hwmRCBDvQETRR8+JJHj4tUkyfaY1C
/NrcurVCc6fgncT8R0sAYvVtaIa1Cgb4Srm5g+R4nMDzERrxnPJBHTCkEP0wFg1wP+abeCYRWerN
YNBsld12LFovEFMqlcUDroVdDV0Ke4E5ZSyITypb2T+DdxTtcthp9vPb8dYeiRz7sJUTWmMS+EMP
8u8PKWYwHoNj5BZ4rV46bW2VrvWgmS6oTXrfBvWHruVDTvQvjEwjb5IcUMGsf2sv0Q3idQqHYPrh
1DiZiERUI8BU4FI5fsCU7FnPN7wykIF7ScPB6Kua6d4CXQ656rUTeJz9fu5e1/3mEvFduBZ+XwJS
GfxGPGwYyVcJ+A1rk5qCaEwK/eD93K1YryMnqn4XCuGCh0d8bdRVM1wvXSOWI0v4GClKPAeD6aLo
t9v9BziaiWhSV/TiWkg9UUlpng5LvqoT4nW/1owcBZGwL/pfAOOaZv6xtUxWpke9XbbMu0q+Zak7
051DmfJqRCq8quMRMyv6tn08iU9ujcDX64Lo/rQ35IDndOs/S1pCFaAsVUHINX6HMUD0lh9DZAzX
LW/3pFvOyH4bZDtdYjB/OH4EnsZ9b3hnh+/uEwlySFezT1J24Rl2b47rok3R7JmmIe0o81Xp3CBM
0VyEftjq6xdpNU/hJs5wakIiIsvimo+aGB3r+3Y1nED2/pJzrtcXrpAUrIaNEHa1nqJyZMgbJpr+
V2jnXbXerW7vHWcr9XTPE7RCJ0GND4/kov5ZxiB5VnsiZjcdcIx1haZlF/IMt6I0hniZ6w4KPKkL
UOysQCd74Z45e9veouJIs8SpAc70YtCuu0tL1x7+ovTw37Wp68UGwascpKogwr/yzL0lLZsDyWoS
UfNXOnlEYhpdgTmuF7Pz3myWo3QiFwthZnOrH2VuejdahrpCEeUd4pvrw+RQVlf/L6Dee6Iy7cID
Q9SdRpmktyGvzN8FeLHK557y/zXkrhzd16ViOHWjDou3kX/aFrSI20pE6HPebu7bU2IjPd21UzGa
mvESKpYwZsCx1OBHpPiccbdGzkjjKkFxi1bkr1L26Jr3NPH4k/h02uuw98eiOVaIfnBst+hffF02
jNavxemQciwwWr3+V4s5ZOcvJUiI86H4VZBTrtl1+0juk6ufbbnjGOXRNDpl67S//9prsqx+5d7D
wQQqNPycCAtQwwPCajhsAzDm19xrBYIBahn3RowB0Y6r3rr8SWugTyfQJ6ruqDRa99wUmOEADvsG
KZDL7s99DtqDfmlDIwr07M5V/5o8ZRBpT7vXVkF8IjsZXeIiVuTt8m4oP5x3sPD5HHl/YVldIim4
/K9hm4f1RE3SVygSVUvwIrHwgw6IGU3C1Z/Npzyn5LqGPQZZt6D22VW6n7f9Pb0okpPnpxyqoGJu
HqF1zxeGyh+FC2YHFMHkpI/junBbcT1fVLNaDZN+t5tK/jCNGbGoH5w6r6wE3zWCbd72qLB+Sy9q
4aILb2UN3/DZ1djyzkOBbqIo8LS5qv6POeN2yB8+hIxJpRzHCRC8UpkJwU+TVcDSfYUz1ovgBpMf
7zg34F4lavvkpcTJCMq9BMvO+HcTLrFbVPXrdrPJZDcf6yndrq1mZVmc1KOT7wwt74TYhGlLc8FD
F0WysZMh8JfdG3e4NZTLtj01pv9gVC23+TtRBMQgDGseDT4FE5Vua7+5PnSgzB0xqRB6zexQYumz
ATCRGFmtofzxk8991xyqThqdlheN6MFWCCZHhbLhUIJE6xxQNbyDaaCuzlRGlFQgPF6Rr5639EVM
aUXfzmVX+q0seL2jyTDjLKCZOgvYNAJmMLU49cT4pQ+r5tGTux004IBUoER6dR41iQUQDaO+tMMw
QOmtg0QEmVu1DAlXBriKV4PKL5psR3J7/NSlA8XRTuKWXRhRuyxUTyHm1IATkiJC/Xe+naCyr+dF
NMLTtJC4FYRpp+4cRBSTz9X8jbwm7gFra0k7gwFx2+MlXlQtvL59UDKc44pyVeqzD3w+xS0smTte
ybrXnz03bFGPbXlNWOWaU98gG1ykCRvtiRlwfSctUFUhl+UvldS1w0no5xpQoyuQMlN+6mgcmNSu
fWBMMigF1h0cGPriMH8mclaLshxLXWQj3Rb2f59Wc3vYtqw9GfqkTkyUq4GS4Ar1duL5IEywZLe4
CVRMataQQe5ivjOYViUarDiHsZ2zsJK4QHqThk3IDKfdf6nZt88MJat2QIiE7fcOGenGV57o4Ajf
SoEH56SFMe+zlQn9O/tyqrYXoEwTT+y3JLExZTKYSsI1Njj3HVUi0qS+Sq3N1a6XJsExE5evY5Y9
yJF6TKn0FAGvJamQdH2YZG1ucckD4d9UDfPkvdJo/4uai0WAI4Lb3fWa9ieDgRgP1sv2l7PnUI8B
hwbbFqcDr7yVF4l+PItOisnoRHQpZlPIPrFCIMMzX9VLwvdsBZlJMOYRPfMS1/Zh6/xok7EzNHhd
BADPuSXWo6Jp4jNBHNB+j8SE1ry8EfPQrKyKn1rQFW3TkF65T6C6hMXtbKLSm3Qd3SaoF066DH/E
XKwXcOiGeO4b1vySwXWhdoARt22Mqv32fag4XUEk2uQKrCSIBVpDRPK+F7d+b3O8/hbzoxVK4js4
MwvIAiv9yiskpK1i33OUvd6FKp/TYIghir9dGm6WKMW8IIDWl90uerQnurkwNGt7pLpbfjmSGYZ7
S98i0KXwCnOos6/BxaNt0WBylFZw1V1zkQTe5FTcdRDElMwoBc2xmb37Z6ogOFfpxuCbwEz7Wr+K
3HSOBOuScBSm/yDXccEmGz5jINLQAmgZRN38/h4iF2CaARxvAgKXj1v6Ycz5A+ebbElR495/UM/i
cMTmbChAO0UIQdCa94BG6nhMiYaWgY/ySkyPVl5jzJn5puVZ8uIJilXOhiLS/ffyraC47WARfMUP
uIBjP5Z6DdfQg60fwYcon/NhV4pfx/xQrq6scstvUqD1arVSZRZR59cCTM+WHoFrNjdFZGi+r3RG
RjjH/frgjhhjjjR06SqsaP+xc8aDesPlqDw2SHkM8VnM+q7rvrcFFmixX/VN8c6OUxzuHz3koqEB
Z2kSnq6pl5B2ouGCH3YJ8pZwZAW9RhZS3nga73Tvg/mS8wo9f4pq5WYCVkhvCqfhQomagZ8l0LTZ
PUABrXG2mAuM0ESshnYOu/fufXc190iKCO/LfWb3uvMRrBI2lbNu3vWpf5D8oXKuty+USSV6YXsD
BMcYzMMehip6WjTFvt1oQCLKvPA9oZS/Je0wbN0OUo2uff//fb5Qq3KThCYtvn/c6veUC5pIrXdq
PxCr8HJEmbB9mvhpSavzV3bwt8pSEUGInwiLd08txIgADDNXa2R+WJ4qlD4oZZWgg3S0RKDWAEgx
GNMHpbNH5KL+EuIkKon7TTC1lTnVjxoElXdJhlyX5DsrTT6AwAT74JBtzTzXydzaKa7PCPSGJUd4
mXoMxGIdBNr1CNuN2FagpNmcjnR2xKEv+gc+qAo/OPMZx50Le8MiYqjv+dW65YCL9fT/IrHotrG3
SYSQdx3btGaiBSC1EL+oi1g0UUb9auTvontuESvqa5IoxyDiVgVmUrQVYLi1pDB6eGKr2h4+gPGh
3SDP4f5YAal45RDrqzb2SCqPKODoakzrPpVg/evhREHC2Q7Xv1eTlhoz6faliHTxfBrEVnuycmxQ
VdBluqOj0dcZ+1xE6GNzlJ2/lPAml+e38iF+jlf9VPaNZKnZLs2B0RQ5LHYp3BhTkgxBhiXQznlG
ySB7Q4jwxD6eVzlDqBQ/MLreNGpkTOlXlTjrScBOr5A152p2csJ/zcW9ZaWTi4dc4vRy7Lu9IcAG
5k43jTsm0498kHIVl+5ag44lxsDYSLZMuun3s2Bp9++CYX10nXbpAK/XBJiskNlrmqj07+c70M8F
IfHncXVwlZbldJvnxsW3XX5r7+3trVZ3rlsIEG9pZAXlTbFad4tpJFD4NI7z6A9azHxV0bt5K0UP
uu9HG7PRvM8neGmEJMa3KjdFkzNEThBSu2eG9hvEBOLqzPiZMPS+XZ5r+qmfIapJfBZTyZEgUCou
V/gOvSUQj3286M4InLSMmotwYc8bUTVN96RWcXS+zW6MMTlxr8dT6sfxBDFfrRaGMinb0qq5ovf/
owWF4oW1rrfT63sVgULD9gBoi9uvn2itJmhJxuA6ouZJSPykpf1GHOKfnqG1YzJhat/jGzBKvWhr
MW2kcXOjC7tX/KbwMYw03oSVX0axCJ+sHL5N2Qti1op6T0vn5rXdS9gKLHCABYjIonNxRf+8SefC
bBQUai4H758dXeAx3WLHZU3EptxULatOhpk61M43UIVa8HtuS3tUavU0tC+QLTqpdLLh/v2dWLsx
u6CPhAYW8gyErMEGxR3fTUjiWagyT0kqBjNa+5KQfdS5xWVP803UNyEysOyGwEW0n59HI7c0K+ka
LqXO42ltsEsl8S7IK4lX6oq/xw0KV4TQ7TibA4uPzHo9mN4HAZEB9nFtDIAESdTRdOJp1jaUCbQF
vzrBgtdsvgLICY/sxBJmd8TJ5qv7oUGqg+rLbTPgnwwHOT/iqHkrkSYHaPWNDFmwzrcc9LjNwjjW
hUCs9SC6C+IjYL1qtGtht1PLDIc2AQzaLnKQUk2sgJyMYeCJRhuzV91ZMA+cP4RIsRZr4SznJidq
9GRbE3i0jPsasuVPbQi6CA/BVyO3YqlmUDbbOpgJ4D5BGLXYluLHW01Lo9VOr4pYE29jen4DXG2n
aExkKmh87Q9tVUDw5Y3pXizV3/+Pwvz/LJl475WhOhLt00JHX0Y+FqgowuE3GqhxQ726Vc07fSic
OjkRwAPRocJHHr/+d2jduLc61LEFM8LIs+dw4g9PESlI5Sx39Mt30Qpo/NAd344Umz6Uca0yVQyT
LDUtsOM10wyP5QbhyoujmakdgLd/DW8IAKhXI5cvDkpwSNEIYndkNYMXL4c6kjcI5pFEd/8XE6r1
Im2dFH5w7mn9OFooZcN9kDsJ/109iGDnaq2+tICc4QT/CFNIaaoh3X2pRldf2S6cyLHnUwmOAHpG
TMt5LMuqyU1jKukq063DCJsYYe7Mi0SH0fokUw6UjYV+uRlTjZ3j11HhbcEmxOH8r8MntegYPADq
bdZs2T98MvTBKcwyEjpf0RJaou9vHYL17FXi57qs6frf2GfeOK2ibWeFcyObfLFPHko3q6+tu7z2
ztfzl3tyw1Mym0Lv5FhznzNxiG5jEjdWVImCTjmBQHOtH5E1Z7/PdHBb6VFKSw5hZPUnqpnsQB6z
4i8QoUwX3TLDmhqgoEjI+0IX8p+Rycd4QGkmGpkGlhHWJAiS6EGMLNR/6qaTQG/jgVjmdXL7CtBE
6dihZddTLss68y5ywMoQ7mGeXrryBQG7TQETeObfghjGj/skxfO28YUZZrpk9rag9REr+2Sffbie
BLiSn4s590Wg+UXaX0IdUJVE0EG3wdIbf5GjGqST7lNSuiHQ2doBxJMC85GBywdeRbj4BWr89mEA
Y5qrRa8CK8cIPuKj7Mjm2akIxXni/bf0xcbeJzL5u06TtnTQiu3FPtF1Xj0DzNLaQGGpCKWYOuma
u38iykV1EaNUGehYf9xGXFj5fgIPjBUfOK8NA1J7/fdCfSLf7IgP8HrnAttlwOE4u+/xC++dhqxt
pmk7o1monJpPdquvI2U77X/kJ+LnoGONEGk/DWqwB1DxCyGOvu9ooHVbZNkvgACbKvJDuakUWYD6
n+3PMUJXfAgyVCdPubsfWyNrLh98qEId44kdtFQFhIYDbzoswb3TSIPzRmglRFPiQsDw0Ir6tnc0
Bn3gouMcIsqWAaGhO2cWVDbSrJ8X4b7o1dg27IBdUXtgSNexhbQZhb9IqTKciaeToVYP4uEKbpg2
bO35bD9QmToGPG37Xuo/vYEemTe1iqIfeCyTNMyVt29jR/v4yYdlzpqaImRTTbvyRd+kVE78hHf+
R+1KlSJt8DqZc42U1AYGcr2CuiHbu+TsGD9ULixeuKEvbyYMi+Oa6/2pw3cwKlv3wmQDQgb/MF3O
gLnd600HiNDQ2Uuo7Wnj1jFEAPxhRk/lOhIBN89VkrO6kYAitLwRCQswPvxHkCZ/NqYFVyVstDjR
hePDK1YRahJNFvzhvvhH+e8HgQIoy9MV/JQFdgGjTKlKRNlO6XjN6UgUbKHI35H4gVfdSQf0Tvmo
sFb9NIJ0dgW6HXFctsEE9f83zZXBjlm/pj1Rj0sAwy+PVHMAEFD1HcDjFf/f7WfBTzqOn7rRaKCd
tz1vX90nsZGLescrE5pleQ6mOlVcfEn+Gy+p2IeEwdJTB3cyaZCLoXvTpWruSf+rwsMoBiq8HC2t
OFEiygDpvKbJbBw/ZaezCFr5/sJexH/UKpZZgaTXdbJDtYgxB5G+LSq/PAoZGcPqbYpyYTmVZt8b
tcNG7ykgvSq8JL4h3SB2QgMqTKHc9JYnl9oD6jG4AAG6ENPpZDMIhIptMLwgN0gfb2A0ucO2ql1V
OBJSyBs+fjinrLifzwyuTGipuQ6Vc1lY0osamzpEtDe2pvbvyhEtSFG38JIP2Ybyu2OjHyITXjej
MEw2tMsWL9cusI7Xlr58M14Krj76AD/eVNSZKI9ZCPWUw/nVCVtlYm1KFPSxhDznsV/84ilvujAS
cKH+qyujm2/kQbfRAa1GEYtBdaz9kYJ8o/olcmXCpyAw6NdKkvFk2W7NMYO1xdap3lYs67/Gj5J2
zvPF3KwJz4rCqp0Hg08ySbFg7mH1ESi3e4s+PYAeGgOmhVHq1fJOmlsrez8XLcBmFHr63uFkK+w3
BlDyTw9ZMiYEh9dIjyDi/wehPxevNk4ok7l8QFARn5cSm2qFeCNyFIzUW73nWkqSiAtTdbnApaeq
hc7B78C3Rt8Aj9995dk3APIj/6fR5DuFgfmazwP9E8X9+Sh73MrWuXGdvp1bA1ic+lg/fgerwzmv
qXqoaHsUoEwpKanLcjbY5HFF9BVfmNwyDWhsJGPrtDrRaHTX0BIAhOMFEojxSJ3uhFQkX8BJbpRo
AwR1o5Aq0a7MkSErVeNGl2PrmJQPapyEGai0j4qOrrch2b0gfTpIyyb4mDAktKbX5TsI9VIjMvdg
fwyXMHRtYL9f/0V6CWrGhN33uqRX1ONTX1bj6eJOQw8pEAgBFSw7EuFH5fuQoHMfNA7FYqBGDS4b
MHxgK/5ifB61Wc1W5r6qXLaJCX5tYgSzUvnCyzDIR1brjqZCECdmlmFv1gLwZ+p1P4v5rXA6MpLd
XVraQnJZdWRE5R7cIopRTdAsQWHmnk51HhzZJHIRMHDrJrBGX+DKoBfUg7C1bwZTcoOfAXCpeIBt
nv31aDkdFs0duzsRK60Fn30HmTHYyOZvKIO0sq4mssktyj/X9qrZSIaNKCuGcO5LFh205UhnVu0p
1FRN+NJApHsCrd9ykfDIQmgc/5ankmNduqgfkI0dbDMfRQxDz1bpvrIyEqL04XSYLXk9wUrWpOfR
w42rWjw462XPVPpLWRxiGevAa9OTo4tT5TicT5rFY1mGPk4ZNXVcfR85CoNp82mrrmfqbaZprKC7
X1ZYO6VztTgB906N8rmyJzFRUMIw8QCjHZIgpi90/R2M+18Z6vciT3f47wgpfDmnEBnT3YPdWesx
5/+ckQq6/TWut4h3bf9D+0rF6kUs6b3ym7hW4I/9tWiNYdCcZKxhhOmtorqrSapOuVgPmpdwkBlf
PDZ2u9uebo2qleYx0Ih/hHHgR3vHqS/KTn30VNbQDJeOqr5pKzydmTUNZympKseJINpoHBbh3245
5YL1Q+scN118/p6dkZFvW4XNoeVCsGQ3ArzHiisC235k5yC+x3E/l0b0jsA5qCKZTAi7pbCIo5/5
OelOYRhUCvDXxG8RobNRireuPWWLjKViFbQTEVd3yTabyoaxFtjt+FYDZ1ivRQ6qsr8jvK35HZFr
oDWC7r2dAZ3Xtw3mJ3ubwAKW3GMHCwdnS3gaq/kF+9slqyCwy+ZlTtAtsvNZMeHNphRUhtDkzjyI
0m51AZIrhxCSOa7lrCWdMeI7RI711yzDhHThh0uwS6i0OahX2ux8cUmynmCmC07HKbRbSVSCLRfR
HeKcS5PaO6imc9pF5kjd7FKIlmd8JGeZqWiNKpyYwVxBnfyPQgPvJHZPq2/3Y+h/c/05mSOmfZf5
PCqklMhEQv6k9Kg8YUjo/hFvWZOrMaqTDEz5fSuKh8NU9Rf0qL9sU9TpNP45v41LOtWt4X+T+FV+
MsYYiYaH9eQEScfQAln+u6LrHfeFt456Ntl0cLJUDXiMCQDAzzJdGFUqGt/D5YhbRtHNtjRthQbj
9G1MXDLWfezpPuiiNwKyByl6hrRBGqYRHlVzrXtRpS+i2gGGCP+Khb0z2dbTGO8DC9kDYRq2B/YS
MH86nTcaExIt7eLjnyyc35VRRR/Z9xDOcsroukYYCo7JHNOcZvT+F5QuRsKNYLXdjlp+CdsX7lEY
amW4Q/Xb+zQrRROQcgggqCGEhaocQuLEBadT3/w4MRT5JUN6b8Ng1te9bmv72Nek5QbkeSiQG2zn
vOXJvLgdMYfLZLsvoNiSILZdEWpDujpRuq83Sfk6IsrDbKRZhVWHJ03uQqsh847jPG+VqgtuJJdn
BbGJMx6M58JF78zSL9hcOg+mCMGrzAuRH0uYQWrmbwrQeKgi9DZErf+C/8DFXqWzFXAX+AiBR8hk
eH7aH2VYRtuXmmiALxtLRX3pzCSSOg/H83f6Qt4iOr7G8F6lhVBaVCKkED72GUSYdxJG0o2ws2qU
NflEgaQDRHeejUNJmTjr1pje62Z4Odj2+0QiXF6fp/K/2KpjDgTVl07f4ksfRAEjXgJ5dJdoFmBY
CmKcXCaOukBko8IBxKp/Df0V28TKKPNQQAusgdmnxP5ILS7kuRS5nXQELYB1eWWeGJ4hVnuEDBdI
xo7MMRZ9WCbx0K3DLf3Wya2lFWeyojvY0WCt6JWENbPMpbRnDx+NxmWiDZ2WNirGrP0O11S73DTS
CMMmTk1jUFsA4lkwY8tNC4PjmtxDpVroj5f7RBSlc0kpt3aAOcb/1M6uU2dnmBYfbTNhb/HPk+vO
gDlwdtNrS2evGcxqcd62X/zqDWttyj6196i3i5RhEleuGdeKpYKs8YUJj3U+S7T69Aglc1Z7qJ+u
P0MikOowuo7uSaquo9XEJgCvISaKOIU8C4uyUYB4BzRsyz2mhqtPJteKjn7+SgVDmiOH7si5qhLb
RINrhdzkuDDlVqQsSQZejNUzC9njrQmwppdTtRC02FZiSGBYrkmg8tzFwEvF4K9L+DKXJOl4Rn5u
2BFSHsQ7w2rluM3E0V90Nu6WmwSzzBr+Bdm09QXAOtt3LEAANcrYTcihZNm2TTkhyS/E1E9K9OK2
mL1sHwNYqkEifIpm2Sn/J24uI6SzzEeZG03OKPcQsiz3SwZ5VQw/gWDhwZL+vHWvJuRVOE2rPGRg
18yyzAGgQl48IJBToIOcLpqV3EwytC6l+R6ZzJzFXRoCQhqEzcYPEq2iVlT1dPrj833e8vr590j7
XaaPWIYGJioJjhUuGOeVl4oj9f0jNiJ1DoGmHm1x5iAGFpufdhz3d/aDHx8ohPgrwAaEjZfJZMgV
3fVaXsfjqqOIsHq34PuNZthyj1Y+k+uVCX09ANzUMtHTo3B7rxaLmfKCuzZYiNDEQ8Osbap8OTtg
kfHOKgo4OCMNfN4E/DsH/tsb7HSlNBc23+hhYE9kx5W+hnDPycZO+rFdJR0E4k4QvFENAn9ey4Ja
zdWp8RkVE9GGF1tznaXZDfJdiiLo+h+kGLw6VltCGjVnJpC2UgOIG+oYLse8c+Rr8h6p4gMHHZPD
9hAgbXXiJfg58CUQyhtM+qaSaLbYT+oL2XOC0WYt6fO/f9lUng5yTrRFn0uCpPqueneVRwO0YGJS
DKu55OMd9Eq3+ra3Le3Y2FSr2QnL2EMI7U/Xzj0MU/KM+WOIFyghMYwQDmNntOcyY86/5zzXxvPb
mz02Ge4KRnAxI4Vv4Cf+5spUnt4aU+tdGQgu34JgrGJEpifKB6J2GjDdlVMUUb+/0spnVAwtEPTD
abmI/ss4VUzFcWqzjnfb9jHbJ+AIGg0J68QOWyJ2Xd7oRu2K9DDtWPbstK+Urv3sED4bwK63cPA+
ghEvPHJDokBp3JOTMi4c7UHFhqp38oISjIcQXAUF6PxFfB8RTRbDrV8X0lCpgJw7YLbNwbN4vwg5
qECWD6MUATYoiIbinb4BxBlJVKkQLuFak6t8HcM/dOpJ74X9kbmTuBga9zkd/TczCxrfjvOZfBmx
/ao4TdlIZgIGSoHP76l0DxR3gfJI8vBxiL/HkyPwUMZ+qx+00WaiJnoA3j70KYnI139e3Q7++q39
n59u5/gyqd1dyTepHZgEqKgm+UbyJuocDrZHN+HCk1ZLDeoc3cP2yxEzdw7VW/zIO+AwOig8G9do
fAD/pSF3ZEQ5QNynNfqq2KRcASkKV6WSQeynObktKcjw8gwTDxmLJamv52cSjGEP+bWkWNt29h1A
pMdcVLE8rcaHKMaKECyFiTlRuyFuaZCeWzj4kqh6/RChcnwUm96pDPC3HQX54CGavQP4RJtkdM42
ja2pu5EMxn3uQr1zeFR+usQ4ZbSyQQoDGXdPqhPBjjMAubIKweivDDBD6pbYESZKEHZ7fIBiiaxW
hvxBeoOZwrHv22tLRHU3wp33e1J8yNvQRMuRwYV67E97gA0YVjIoxU1pkeGVn+TYv1a4Vz2xldka
9CcA4yM2X/aCl9SPmsUVdBKURbW44iuLHlB8+lijRUWNKuNnIrLyxZvvDpT6V7U2TggPBBpprrVW
23NC3aqCBO4jq50/tHWDCnpdpJHAFxyr+ZaucMfU4c1LE9fyZ8r+hz9ltZJohmuITZhy4BVD2Awj
+JY92KrwtCq4akrsGS2CF2IcX9eFIC7etIkPj6XLb4tJNMG/Qcs/FJPoAeLLjWxqVT3bMrx23lWH
6aN64KA5NW4PeWBm17E4VloC6KAOBN8ByVtBXbp/TxbMj/p0z0VHuaF+BDXiTh13hrNy9NER1fxi
LMHhPXvm+15xrHBdfulbWPXldRwjd9bYAsA0UOCsQu983T+6T9TtTgL0wvf6NfI2cjHZmHqt59VE
5A6ahdIBWeJWJ6c+RrGj1IJYR+vUlJFAxpcMBaCkUViY7jO5WpximxRKc4yzI4L78ige6EysuzGZ
wICWXDtTvDd4mZziuJMAYKgSJ1ou9dCwZSPXHw94Q351uNHOXIL1Ul7SmON8bZ7u6Rih2PaEAwoH
GBm+P3jaPIMtZzoYYItIumybij+m70/o+rocbs7DDY//jNz4zMIS5ljteBvXDdocdcxf8wueZz/x
Ua6eCrmRwN4LxpkpxOOASgkjv3ekr2/ywPyC4oM+BOU4g4UyfmL4rHMYP8S9Cshqx088CMi4SjBu
2Oh17lYAQUuGRlpeNzFiDkOnDzEeTFhKAqHfp7j1PFeZ9b+c/Xrf00Pjjt2rgChQf9DGVQdxdJaF
DwIlBxjNLRfNrX/YEMJcrKeNGWwqZfQsXoLmbYXM9Nxu5gxDGNAAU/RZEeMRJc7YZ9eZRzQyGVlM
t3gEm+nIh/wl8qKj0akUizcipoVbT0gv9nGa9Odtd3dyFvZZ+PZ+qtsrau3gBsrlJrOORMPMUXgh
xdlU1v8rJ/4o3q7TNoGmpkprXCAhdNkqMpUYHIfsAqs855vRrIp6uvhsgVCfSr8XLjs8KfjTXMuP
qk/DzTa5k4J7z/lzdDzZGAW1VTigCOo25VacpjDkLX/PtOtcbn3KKSUJq8sYQEQ83gh4yi5FStCk
C+hDCXyzC335Ux0l/UUGIrxYcGWKvPDTRxLAD6XeQpkBG3eeFG5D6/0yISZWs1LOTaD0Xwo5JFA6
jDPqN+P8dmnO89l8KCWJgkaUGafB3kEWC6kFAWzYSd3hxKX093V2BHau8LP6lmrGLlpJ84UDsuAi
0kS4vZ+J8vZkCiGskwtdacWK+AK0KSndtO7/eM8YaCA8p/V6JIS9l8OwcAAO0KDO/VzNgRGEEHWI
NMZdScxxFeSfs3RhF7uhFQ8nbaQ1aaX6wy6CNz6hoxcvZN3xr1JGHE3Vj+JZ87mI32DvdZQBNBxr
gcxYMsi7KO7ScYHywtqy1H+JrJaAAXjjZndMqoo+FNcMUqZ0yddrRp9BrB75N9eOqLqjlB5nZCjE
KEHiEt1HK1FqDPKdPuq1SREsDIhRDuoueFvA4R5x8IkIjtsY5vei0ildVGH7Tu7gi0TPuaDCMPLw
BKNV616HztlIZLhGjync4EDojZYGTBo1PL20DYNb6sa6FdGTjOPjruSRZL1j+OLkOdw2Su5IaBAt
Wd03i+0l8Vaf/NJMBfoUbG4d3tYjViFbkjObfg3uDOuStXBiZb8LGzVrrIa2Ptxz/R7gHr2P63wU
B1+ahOhHCS1SEICJJknzwnkXoAAi0IrljXxadsSKPgbi/4Cua0/jPay0CsvDmiBDQitHBV7Jqo1S
9Oa5hmVOnFsQp+6izj9aTnAJqho89VzXWS4xSbdTGoliAUQHRxk9vzUmhx5hSER80QfznHbyusS7
AkcTUqzMyHNelU6WiJ57pzesLpbCxt07vXi3Q+b4hgzSc+TqFyVXsOU8HWj/a0m6HNzx6Cwyh7vg
p7Fddsb4Uh33A3D7+epUHhaj0gmbmol69QnnWoAmVs3cHGrxZe7RN3PhJnERjEcMlxbPmYRDddZe
rrvl4SMX0/pu8dfWK5sgGBI4Yz6f67NxowlE8VqV3oc2mv5fAuqTqjTjJ4eBYqZHndDMPSTX1G9v
FWCLDsSireBmfSn9MQYHNFNIo44TNezKpcb+7raZuRCOYyVfQhPOy8BlXK1vGW78fIRq8T8YHlCv
zqVqRG9ryAI/StL2WLZjd7KGTRD3fyw+y0QUL6N6HUBlqgt9W7iWn1U9mijYWOAyrVe5XCyKazO2
ugI5Hyl4xDev594JTogdN7UVdQJIi1SC7xAyqg1W6aZ+k1dUgcbJyxrNThFBMuevr+QnCL9tVfR6
JXzGHPPPqDsCXnFOdk7qhzXzT08hCmjkKhBJjB6Ae7njVYeztjBkQLxzOEzUDOEjnPb8Kp1a2ePk
66YLcLJjOoP0dBWbbsDZg2WwmC2wVGQO7aoewYNGRqgOYc9/0Nfnd190W1KyfbqOOZ3LPGhI2Rcl
NqdSJGfzTPXgT8Vy5HgcZTZBXsT5wagnIq+yJoP42AyJKGyjkjTuEanwvU0Af5ZQBXwVx9r/hKCS
GwaPF4V+NSkdcfdvMYHpcsviCACSXF9LLCdM9xV2zTuptkFs8nDP4hGYWeZwFqQxxOT7rQ0RPg1n
ZBd8UnowMozGwBRWwv8JfTeukdPey//pRZXgs4de2EG9m4VxbxKOJf8GZgpNLzprZAmo9S/M7nhP
yR/Fqnq7LpboalhE7aDw7RQRH7TTyKMP5AV7VbwPkYFAdDC4ohBG46vCinNd0bFAbOdEjPUg1Ylz
tLtHQB7DPTqqnhlZUGYPNwTQ8AfC9WOQTl6VYOL43AIUKIuEWoPQfP/VsZ9oiyUE9FBDfeE/AYaW
3lKmxgYQa2xP/58PhiTH6EXEbQ4JhaAKeEkERh9lKONcfD1tQUtx4bN0awDzhUso3xdGtZS4kt8d
+4UrynDPeRMzENaRg9KclKvXbpm00uSvvXXUHnivMGpIalYx0uF1Mm9pbjTp68lWu8YaWIfmXztV
IIRpwFm+OGT+WofZvDx6EqKXxWzIshCUxlg0UziGz9Vk9i5N7eL/cOF1sARJ03aZtVmDy3je+87D
NULn1YaNek/hyb6GP+8U6i6OtxcLaQFO3fV3+8wbe0mu8r/4fNjNxH233U8N28pfctx5lXFSdq81
DrALNRgw2vztcppu0cnVyj/88qW59tf/X7/f0JJeu0/skbJTGCS0y+SZE1unomGZ70bBzAfWx9oU
oVj2yjRMTMZq/Q2inxZW23JvYfBkd9a/Xw+bRdN5zyj/5chP6JGyhEv62+9bnxfeyTQsQr0fuewe
jzCPbjcZ4cMI+YqZnKn3iE+SR+o3/lNtDxEumfHuySyNrpL2yg5lSRTvXVcLoU22tS5YBm5phPOV
kI/E/5HouONnHM/C+c/guASFlk0M1+OCl5G6sEpd7LHVrFHms7lQiFlOo5DwfnAUjBQm4ONvDN9G
YHva975Y8G86dNg5HNmS0yYXFkPr3bvasQrtk9y+/woyOzk2IQdjudz8ykn5uNPpjvq8bZfhWiko
U7bD8AJF58ArJ/jiFfLKRF8ic1sc/IOOofNCixHUyy/p02NU84QFIstCITdzL9Yk7SX+pJZlxFzq
pBbgXVoWPyktcO3PJ9ods5fOc1165maKK/cPuXozR/whwlwmsuKW9wekC40A2GOvxrVqxWlQol3E
eOxCU9tA3axrE5MCXcxDjsYMSySdB5G3N1XqxOXzatgoyUxjr5616Idkpr+BTYRy1+BH2aKnLJ95
/3Pl1WWg4ljAtAYlkVJfWgZVwPsZ5XI1t+npjBDcip0hq576fVM95HRuZzAQUJvKRZ0XXX5C8swP
Y091teiO2P8qIBrFY3YONf4n4f0Q7WJeVRo2PWWXJVPwhwq3MX+NsjOuA2NwRQ255Nw9kvEQMx+d
sDzCkmS/z1c7onxfd44TEtaSkINjFeYJTFXTG/yMcwILMUl19reR8ukR5H2PgOfq+DMzvA8Dcxdh
J4VSeEnnO/W4O4haH4xRSlD0AsOOCMKz1C6wBa4ly84I0Znk8e78u2QOV5t8KpLzZdBmwrT4GMqr
9R7zCivF6+hN4pgLe85JcYJVFa9IRCh7+Gz871lxZnLsWb9my/X2lD4kHc7V8M2Pt8oobbknjNvG
nI9UcFxiV4rM+XNoxBDs+wAv1J42Kx4OYIP2CvJ1/QuGWvdd0CcL5XJksztTURGgImaieeIg3dQZ
KsRhezD8IbxaeqLIXgjR0gscd83DNHQcMLU4HK0ZIiwG1J7kLJb/U/aCSemVTS5qYHMX2C4lhC8w
Lus9C0H4/S22WAzT2hndkg1WuAY3jgzAhSrDRP/Kvg8OWjw5ObYekKhjOGDQg7rEgUwmJOXWHvso
rrC4y5zAYmxpJNTKyXqoA4udk4jlgHOgfklJRgS8ikq+XIsjYOSu+U6P/oRLRbeG/mWKwCRtKVMN
+VPFgtOchsr2mOMExkvuj3c+bSe4viIo4ZPzUNahvBE0KTYibL2x6J9NSZIoxqGcZCqts5ShnpiI
sOGxy+DB7j7X1E224OQpBS2g2HQ6A104JqbUGYHpL8oICeD4lYuSn3W0wjwyValAHLXRF7E0gnL9
3+/TToLjn82N8Nk8bWyFWTF/z1yqjdVP+ZJBbe5VXcJv6DsTKjCXqT3XMt62VTjgrQY7YMVeEn8J
0R11eMO26X3VFQxIYKgMo5++Dvo3RfPXLfgGuOnZ7dXBDrclwk0rXeF7bt051MPvaKgDInn9wZ1L
7cOQ1rOA7ZttEkHnOKYnuqXwZSAQ+b12g6rW6LbX1BWnWhzIYkP66wrLo0EpbcKd6QbLQjDaFYWi
+A/lSMTjavl7XFMD0dKZ89HfvgnSRLIh/6ibxUczZv2SDOGVhl7tIGwqDTrk16f73RX/Gm+MtMEd
o4CvKs+bEnbjNQTybEwS5Hcva1tvGhftY/M5theIULVzMsWiOKlXvccg/JSvJIMSfWlA8yEfcTTz
XMy1+Z6s5P7+/TKlGZqf8gi6fJtj6niBAwBBF/OnbGZOWq0dpCJHWHDkVFy4/NhjuNqQ3POd++7M
q9hIwjhLcMfr1z9L6MNkPcczt2YrbexkIh0VRY0keKYMllYK1aBAQgv6r9OaldF+4EXVfXAfIiYu
mN+LNR7t1g/5JyoRkFbMeXp19zeeVz03mkVe46bXtQiZSt0KXz7AK3s6x3QvOKInmADc2gd/2eei
znI74LpIkuM0crhKBRZynmRMr0TPPz+EQcIr8x61/NJjGve/xDqMCUTaHSqqa0BzV3ppBkVKA0y0
EUV8H4plXzGcK2ZrKomc375J1AuXRbXn5JtAPHwmELmY2YumdkFvLpHk+OMfnNi92gM4kxNEOkDs
esu+0hHLICchCEfCw/uvZFusFyt2DFhCfZcmpeB2prRwLAb/1XriHciLRrQWotP7kpASRKIXDbPA
dYFhjKMtZSwNu3W3loISlwQrQL0ILZ17tKaEYJlneVnw/sd3DWQ6yYZy9xCeiG1XgH5rIwN6ZquL
mlww8t1jUHlg3LFoWckB6leW/GI3scjRsFZRgtSB/jBN4JcTNrzTgCTDlGOANKPTGEze41+nRRD2
4t5YRUaOzoSUVZLvYZ0GuYg5XqYB22VGFl274GF12OHNuUxEJvwwbSM9FKnC2ymeUSWIhNCgvcYK
JIrdreVXU1deVmGeODZzYKfD0ak2FqgQPjjBfYTVBv9Y9Ut+XjQfFf8fNWIjq5Cc4/3I0dlX3VWQ
aAgy7ZKqj2VhFCROaDE6X2Y7E0u9iU7n0i2B5BX8ViECPWOIJacIfkH7C3hUzUeTCD0A0db2NlZN
qO9xrKl0J0GkLXKSxOMmR71gIyuH4qOd8ahL0A2vDnU+KzlTxW7wavIKSv3S7UporMSkDxfJ/duZ
nGPJU/drEmhzKnVRA6WlVCigI2idTuHEVADY8RHehTJ4GuZ92efwiVW2LuCtOB5vFNlojT1/l5Yb
/cIWPCwAKO8rw53a2zNFegnOTwQAoNA5IuysL2AZDm7kvV8IxeYNgQutEhTTblBPl/hChYC0QgRt
x1+zvi1jY0SV4/vxfvgr2GdpUtQQdmiIItFf5dQ5YSXtcYw69LAVPh3uXxCePpG24+XDqWPWn9JX
o4M0hirHJ3CuDHv8LNSa3Z8/BTEBeQeN+8+q/GSRDp6/QX0c4dLtF61Pv6TBTJRv8/x/73VouqGF
NknmCeNdQoFIlz3G1nmpvRYdRcm/aEbnEaNAAioPIIKjTKfWSPoxaW/4gA1eqYeG94vpBx5sWFuQ
I5kKsnQGoOAxVt5my0I7Eyr+X3TFkp1xO2IRrrBQGWJR3KGASE4+59pztp/Iy8hjfrPeDTycG3CP
qJJoNZJBSOyckW0PpeHjZDhVDXTg+oe3D6pjvGcAV8AkhnPCna1DSTYbKyVLZLwQK9Q/N2IEhvsX
2LtdeZhFD355/sisegpdJuVrPJTKdMzDwoX+WQqGTf5hcieINstcl7567/a8AWKPWtL9Fk6c0vOb
keCoA1j7eOzrEHgeK2jDeucOQss8AxeRGxntRqsRdEI53dwNCmbOHuB8RzL8eXaUC8HQDr8TL3Ys
7/CyoCL5cgJP3ktwSwk0f4OkEsm1jzyOKRiqpbwVXO99g4NFkAGoLjH+nRgo5MbpE6Xu7wP6tbaV
sk7jHcWeusrYDUVJzdbQd9Rm6fa/GcR1mlFKh1PlZ90qu+HFVWXEzzB8hxFLoX4Vgo8gXQz/FMDt
4960I/N5Sfehnwe6Oh9wbQ4ikMPLKj9gGZAuYe9dycL1IDQ+a1dG0yFOIRxhAi59axeLyEKSMZBF
NJsgTE4MGVZdlhMwB4jJOACi66iuIv14M3dSJDYiCMuiA+JMNJNAW3XLxbczjwWxHsU6qywKy/a5
/LyrICHE25l0oQJ2zKmFvFwYFmCioe/kGG/FgAWccqt2iAvrqrnTfx/jS9NqbRobvT0OgbsQ19Pk
3/bbDDCshU8Zx28ALzlFfmbJ7857DWbJ1sjJfe6yh08gNgLvkaOULwOYuW/VWw7a6FQvvPPyZ7dl
DBmBAfCq4K1OQ4KCHOpXdtsa3kqglzzHnSZ3p/a0Oz3Zq53h57cbRZlxlBIug6536mJmGMGcs+FV
xdV686uWslVtMh40FqvcxDE2/XSE15v1T/StZJhqo2Tdypf3I0yrM80Pz2mulNF7lr5Q7Jc62t/k
P5y1Ieb7jEmVAO5lrw4I5+o4fZ5nZUq05ov4ngcdW7VjYUMHHysrCBQxBMWRkGErwjh310svBvyX
xn0rcKC6jp6Zt/qtuyzLyjHgGxhHuxdHJnKa4DkxiS8Bd4GkagyAu/K9ngPXSTgzQgkhvPShpQSo
2PtPIHOiGAGfepoNRup8rkmAw+wKkorXMN/b1zO54eRrUoDWZoIlkAuMRxn5VS1tw0pp7YKq4mGL
2APnpf4jAK/Z0TGxNqIUOmEmvf5spSF7yZ0BLXcsFkcAFKQelE0BU45TUUs41pPA44dzpaT/3iiu
anILAI7VvzVelxbn201eSpcCOP9vqFROXn9qZskGQ+j4TtKg6g1iIHUmU2WogsvypCLc2PbVW6tK
Gte80ADxBAp1pGsXnfS3MY2pijcq/1LohqMxtaLg4f2DsVItUCqJ1id0hirkaEjKWCk0+evFrc68
EPiAskGrREfbEGFpcdmPVXLwELcL6XMJ1d6Mpe2NOede0B6yi5w+BEhwsSZ4pQQZymIYLQWyUNy2
Tf4L8fTMTeKAhwdHFBxWGdsnMlu+XDWYhsAe/TaGEpdRz8Jj/hLgxy+5c/m3q0ddDThe16PCPlln
2pukveCxg330BldtHoVSvXWiqAqvkehNw+s4pa9hUWSSN0XL+406n5WQqaLdIvW5KntN6a6JU7ng
Xa/MVUJ2+TIbVQHvXxi+oCNbnzDTwMuJ2JR4ofNAh2w5yCsXKFnmR/HwBnoFVmgSbAagVW455/cx
TUiIWdloN/yTcetykqRmwnIr/GHdeXsqlwLYuDzbwHOEKwKsTW6xjzyMmG3uS7rX7gOfjmQyZSM7
A3JnGitSsnKZvy31bpY+aBDlzPqG3np2F1sUnDdwgvm2xOit11eU1gpiDyZMwBH7GZvG6IhVcpkh
JZsG96uuhyb8XMGRZdE2sZJ9hWTtzdH2WleeJfylWd8wg4u4ruV7hYsZzVsil9uz8XkwPZnw/r2h
NLI83lw4EjbIfiCRFwBhcVbs46PUGuh2DMVz015ZzKJdw2uNw3Ow0jF8FIVSiYz7vX0f+d8LNCrA
gXal7c9QA/l66mYscKSX/GBUCdyO2HCczjIOPkyHLA/JW6UjjNz8siGvjvCC/xXdKg6fK6IKVUvC
oNVkwsLUKaRm81Al2p9fpjBa70BUBgiaOSU1M4ineYDQaZi/XWJ8saexWZYMnMDS4+uigXuQCah1
kxl3zu16xgZekHc6ecGDy/JAFo3NGeH8Zam/e9Z4gxcA9LTviVUzYNI5gNwX3P/fUhiltr1nU71F
Fcpjg5SFnqa9zNMDYnsz94WqtjSS6L58o5iIeD5333gf8F5cOW1f6lueCyRb0gGw3kI2d9DOU+Xy
g0Z3UOW+ALy/BFNZ/XdP67IuiaxytzXajt+s+bRhjgdXMz/2FYXtUJUijDRnSQWN1PyvptpbzVL0
3rc/NvCd7pVG7fW50RS/+myoSZ8dB9klrn4tc9uJSaVFC3xExjSSRiS7AnqnTRn5wmYF6QNPdCLk
EkpzLnCtR8FvSIDYQcA3Ieic9ugLDOW+eocb24raJ18ap4RauBujbjeAn3qgMW2TKZG/aBw6Nuef
UxOGeEI/7TvwGwYSca3D+cR7ydgMOOWfZRKNp+f2dYEJP4Cu8X0GFKvoTpcQpFkK8FzsCvUG8654
OCTqZ7zo9J6U6JG+aEPg+n4wvMmV0hQ7xZYozVDo3h3oL9mv+ny76yP0NoYifSpCzp0pnLnU1lTs
dZddY0NB28c3/g+tzpxKgVzyepVVu9rxmnVgF/NYyS7uMSB0UhKNU50BJNdz6yrXZ22Fg8LEYa8U
vXgin6mhrb4FDY/B1Vrc9AkiKbiwdEEr3qKR/xJIZRUoZdAUf1nK3tI5jAhBuP1Cp7TQJdJrPgd4
VK/67aeqmdLSBp9TzLmyXuQfu13tWi04IAo42+0XNiHec78MRx7D/xr0d06H47fZZIxZBbx21frC
KrYne7B2jEqEQSt6vXaH5sjkc950vUmubcZUYb8UpXRKc4tB1vV2SVuIeyO2KsS3YZBjUuhkbA/W
F1OsCbKgPwGRH2UaJqTCJmiUXb//NH8mqJTg+eS5V+IMXCVU8rfAH7vR+EKF8g/S/4X1p17j6dAk
2hnA861sLFAHfwwR9ZoPG/WX5yLKsqnV2o0brbnZW7GZSSwJJn7MR6+iFdird4sCyouUgtUobjsD
uCQMq/rqgUY8dcTEMejWh+26wyzkilCGh4ax3HOEWx0hBkN7nlOBtkIFR7XiqsXiuTKws3FRpwSL
TCu3ce9Ejbr9tx5e66SUQkfDPzwrP3CY1e8PXIzzDgURzA+Z3ooUdMtbQ+jPUSwlzCi7fWROxpMB
TMYtOyD5q0aHVRQNKiKHz4Z/zZxQQtlvfnsdIt2+ueAmBIeLpGa1f8S9R/E2XEFP7Nth6oAP9aUt
6vIHTntGD7W6U7Ej9yRa/cveYeYEvM7zb/O2hbG5dF9ac7p/XRyy4nJsPetDl+JxgWdOrJrRNN4b
QD/G0wcSfLlr87k3lOszMgCUVDFe1fHPCuIRo/EnE4IKSKsrRbGWEzoP82yxP6wUBIB7NYOgmj0s
GbHD3WkfMB/aaJDNBzPN3NEtY5VE/42WVqbD7Qz6FBFG2bN5P68FsgqG65FYfL9OVkb+7dha35jM
znIPbLpdQGrCu+jJTARlWwSmEujrfQmubl0Q1hn9/RLM/XOGq0aiU1ZQKT/80idU9bTkapIHBwNz
6RMJnwQMzr3czbwA3vJmPf8tAjnmz9hMPzlF56MUIrLT2NZgy/FC32+dFGDZpgKxgoRZ7BNoK2l3
IsZMzDOEkt4MmHT+Zc9AkWwTB258EAcL4zUWZhnVU3QcUoWAvlGp/RwgkPgtrIclFE8hTAlJmuEr
KjK6Lb6cWoPx+ZvnoKj80gW3kmUBygvEkP4IkCtZ712hsbVUwCxGKxDe+Blaw/x8D3fb4Bb9PgAB
5jPRxsAfURINuvavXTtxUk8MKdNrQhJKu37nf7hX5AsKPyCODOjY3wGhtpB5GsFHm9labG9WQLE4
nooMFty4zYOU/GIub44drXVC0TztS4CN5Bhs6JBzxk5xdhxfi/EMzpPMvzgJMOCiyyqM0GfBFSva
iczOVe/AYFeKCjbKGOwPk/s0WK+/JUWGs2YWNqlz46Mkvtmu4H+DWWPEOmCUnZ9RQjoENQD1oxqf
owfhwIZHcj/WKGe0pqp8sk+BPOs+9JW0mgNEM095h14ZqIGrXMaBWncmEiPLpaNyvDZ6aOQfkyNJ
jVunUdAQyHoiigDkVGs9zoAQ47AbNc6p9e+d4/yieQby5VSmq5XxSQqX+ZePAGIAmwlzEijjHxVf
9keezEtPz2/Igtgp6CueoOc4KQnYfkmddp4zC9y3AwVA0+4PFcymUqYMxmDItJU8oGMxg1XBCm8Y
7g57N4xyqfrAiloOUkKP2b3FgsAQ9SLTitCgEj+ChYn/j8eIEWgzElMCGv03i5xYvjkgNCrCmWEH
BJDcJBxXqe+nmOILBsagPGeoWlGwxuIVOfuPLIEeVr0FTcMHgCqWM+l6bf6SkMzjU4boke2vDc6s
XNTWt+J96dN8ufjMPrOLBzXqe/39kayHIYfpDA41SdcuizyzooMuw1fog0lGeO8f6AKMTnHwQT25
QyfG7KLGNBOecrjYjpgLPndocERbwc9+tnzSspR0cvombbQj9wNqQv6yiITHuvo9PggwGcuWZidX
fQ3VFQLlpiGme1stLuImZ7sxropH7XPFmvd4H5YXqAINuHbKkb4cd6kHWxgI+NutdKcrQclZAgmM
4Qv05r2ajfTi+gw7wtAX+9ZSh4j2pYgeve7EioU3JGzcDOBxVhnv3GKwBWoNxOLvsiYzZRWe/tYj
dduhjq4FGz8ycctBxjon5Caq/zgd79GCdqWdqjI6f5BwIitizcO1zAeFplzlQ/KaJ7t8vhHnWEJC
kSzq5kJX8v0iWtK5N3uuMm/GO/Qx5ZgdXuLw7wYGCoxr02SvQbu/Df1HDE3AmI3GraOzK1tXk/VM
+Wb3ej91lA32eQ5slC5/EE0ZmBoiJdfZdPefJKcZtPeE3LVj+Y9TTnZqq7TE8KT0kbzGnudNYiXb
NEXpmY22cgvfEYpT3s6LYN/K2ojFj2+QxxbGDYqvoqM+yBA141PQR+eZvjpIG1N03w0Rey5HUizA
OzM+NREW/+ZqdDXVmkBm7f+Ehn5G3EmpFeYoe8xdEW/uIqT38NgcdHra/91otnjxDsU6vxKduFHR
Gl4HSljx+5pdK1zfXPNnIMmUP10tLGKAjca+3emXe4SCPUe1cv092Rg8d1JUZct4l4RAVwCQgjuM
6CIi/xXyXq5IQDRu0K9l2d1KYxH/aWqO55u77dxuYTnC8BzdD9ID3N2Yw9udZarm9uZM6rCctNys
Gxc/1v2n+m/bUC4qkQgGeON90qZmv9a7jxT+nNrHsSHq1oi/hu8B+w1N8nHURXBO+bGFnSs2zHNV
vwO7NpBwOA5zojq8m2k3NiW03PHWhKiqbLLsr4vnd0UYCAkdhXYkYVDBMXO7gFrLRZfZ2g4/sUgP
u8pZFxuoc35p18DNfW9+ld661DXj/Yn03AbtKFR/8Ulz1y1g97wt4jP0BXpiE494/lm36TCGHhhr
1d7xa0m2WEGSQvAOn3IEwHuSmGrUn2QouD3CYPyNlAawOlsypqHPFdz9WLguCqJzngGVe6eD08+w
KOQh1FLBQ0d7cFahqPLl7JhR7ySgfGSP5Y0Dq1B4mGrMdNIWMSZnX485+nu/dkCjBTbh9n7gk8uJ
YgVf/dqs1YmnoVI06e8MYwg7somwTvATxkq25+n+nYfZTs3TCAoskJMgGvhFOwmiQqdzb8OdQmKL
40TmouHiN05HNx0CYfOqdDO/FIvO7L2XMYhE2NHeGboVopNGJxaSZ1aLptXRa3L3CrA4XoTg8UmI
fKjFKnEPwY14Mo8J1MBj+J+/yCtVdr2XrkgEll2DPZSQHz9d/wxlu41qQP6LaD/HHX3iwCrc8yak
FkOwDTINGHNsfZtBrjLtmNeSyIcVtN67/CxvqT4zm5TS1ScQUK9kam2fGpL4g8TJdzC9OqNKTv+O
IywOJ4363UD3aE9bCD3CcecnjyZhQyEiLuSaup6yv02eI7prz3Gy98lQUTKcvWpGPnOsmkhEbwyB
Uc3VMaz642gx2CLKUElP1ZIjGsQT1qwnoX4rVPhenSlibosii5uEStHrGVkpEB+keDzmJvwR/DZm
IC7KNxRm/KecWVTgnlmp8XRhCKNUDDJ+dMy7E0XdoZ81hf8XDninsUczvN3yvx9U4Fe2DD9mgZ2k
X+ESYmy63N73m9rumXa9f0Ys8PQ3+NoKON5gcg5mVFdFJx39hm2LCVbr3ss3nNOAdfeOBNUN0Exq
2RwTG3r6bUXrLbOHa7zn/7DaCsanj9Kw6ptPiOoOScg0U7B672Y2tpSJtzQNUJxe9rrDg3aTyeEo
wKfsHap+y+2u4r0WWsRKHh9tD4YS1b0XHtNLyyqkEP8jtvGsQeMaIQNndEbom0H2ASrKdxxDWY9V
336WfYnc5rn2dfxceLjfbC1Wa9mAy2guXuLCPGNPYxYse1z58MALeeiWRCttEM3+lvkme3chdT4D
D2JYrdVtAwhXeVEboRhzQ5/mg5GdUawl/bpE1o6m0LMOjz1Fvd4ln+VJxXQaZBRY5TUgc/92Ns5e
LK1msePkNHOIlAI90LEeye0sQk9zTqg0oFMMpZX1bWIwjSWoR0kzc5hnelU5iJvT1G9NAg92ExnS
YF+TtWAAHfXDsr3B7GGQU+YN2pan/6m3ekJC4CF6ZGvikJ5VMwQ0tof/B1GGD3tTanm1Cnvt3jgM
55QdOOlJjxB5K/gdclIJA+FqGG6bity/uEsaXfqZPz9YhQdNubk4EG7GvaTcsCp72ZZKf7wf0Vqr
FK4bQqaJePmeCDqZ/DhJCQ4Hih3MauBfgEDRrVVN+vGmhx9dbkclLfcB4TPpyR6MLBaofSvxEwIb
O9JvAT/KMOrpQi9McTTVcFKHU9m0i/v9wIntjPbtfl04ZevJDZ4zk7CpdSsjyF4ARDBINvp53+H+
MJDbnVMZqa2Np3SfzdZzB+diFY+vvgpwH/DCVFCjlJZW3pAltxIMSIlNwgeI0//Ari4ZLfY+muGt
4vmZ/85oohfMuIs2/DhY8rWOT+OpeHfWWkf14Ac31AxObibE2npEFYp4fQkOHQ4xMxPGEjCpUJke
mXKkXzQyw4OSkRvaZBlYqUqYOPzMN61oVwAsh/ZeHZeBFryK582VFa+FMHanWDDYi2iVeEImFc2t
vnH6ZjwGi6+7LPUaHiMtUPvrjAspnVf44eLd5JTl0EUQu/TQPSOyoxWe0ovUy9qR74SDLAygGKTy
qDB2bMCPqIiHWWFHOe1Ou5MGIA91e+2fghjihu4bHNCxIkhr7YbNOXovvukkMPfKhvKGh4FDFtTQ
exs/MeZ/KZUN0TmUo2pyd2fbzWUGE4eJG8JnYb3Ax+rDu6nPEUQz0j8MxKTrNuBYn4zeQKjWpiiP
vGYl/BeechQMAffFmgM0ml3wXlH3DUay7/6/7ZSiAaEXoMPBphiMcThByQbnfFNsMMlgylG+jdyD
zRzjDeDfvM/2eT2+c1BJWk9tM8M53cMljTrfvZ83WtMgwUIL+tVa2SvySvYJQg/BWWC867z2iapT
dNlTu528Kb1gOVL2uLfV2Yh6BQfPEUFB7ffhwma03kQ+7sWoe5erBBbCnj32rO2dza96o5cfO5vr
dbSJp64kxrAT7JQrJGKs1WWsiKnmqVB4ZaLRtF3TKSDid8fv74DXdmE+DTzllNRe87LjTu4n6Mdm
19x2hQMomLEhEHHLDcAg1VDH/hk1MPx1IJXV9Tyb0+Zq2tizpgHCHfJXx/1IrIF0mzcs7xADwGqo
k/P4aH3H4iuz7cuqEQXSKEgy5I6jTZvBBnkRy6PwVv8Hs3JKeuOsFEhC9pgnUXq6by2Z7czIEiDU
RASg93iuZEKIQ+srPTP0HM54SRIncfzHOrEheSXpctRht0mbdPhfUPWn1bi7F7wBV+ijLoihpGg1
ri4caMmKDbvwuWiA840l7aemtERDTiS/xQcZL2U8LMIqZaeChSvfQ4+EtXfsjbo51tEcu269glut
PQYb7G5ysqIf8yEQmjbAzdTUCGzsgyCGHnF89iOtvK+kq0Beecm5+EN4SIDBYkWUwPOTBMng378y
u1jyKvPn+wqqk24m6PF1Rq1CRM/76iqmV81aVN8nCLawdObdTB3QfsaxCmm650oNSlxyPGhxh7MR
RJDcTRebk7vhNvcqkIptVlQlCMUeomBxif/jeyI73y6HcE/N8A4MKnDrcCmS88Zx6/gnrk8uDEc2
k+bJhuvMsA/J5asGwAkYgM0AvZ9mhMECptGCxQE4PZAfvqsTxz3VAeYrUkIN42rMC325IOyb1pVp
iWpvqn6OUx2Iqu/7Pn1eAiBEt38mpYFGo0N4eCYPa/cyjIDQah1NO2pLARa22JIE8cTXyLhJe4wQ
EfeRKHO5a8sc8uPUAedYUFUoJUqvakwRhQjhheckUgP2yp8L4BvCOs2RhVnSwV5gah+D7xKQhRUB
9ecNnIDItAp1VIb4ZlnNCxOdy2vml4scOYs80U965rMYNp75QpFHjNA74JYmlkBtpC/7rZOa1OOl
ijekpstxhw/A7+O8tTxm02ttXyyl9Rs4ORR2iAqSlxuJDWWljyXNKIAFR6C09xw+r8PXChy0TyQs
6nUYPeNvvT8qew9R0v/a9ZicAFlO6nQt52l1LPkmTDHXsPRq5wOXiCdxpWoe/iWz3s5G1c3whS/3
E4GdNjNXpAH//Nz0fWrMIyD5URN+enWAj+qI4gZHL95Y6+3gryyoNQEtVBei9KLRfDYPglXSGPkK
0w794qAfdoEnduh69S4Bgu2Aw0wpWNRdTUqlvtklpESxp8y6LHD+y83ZveqcHl5e2dZg3JxLqwgV
N/eWHrhXgqgHqCHgr0y4rv+oOCB3nZinoq+gtC2m5rbz4mUc2SZuTdp01z9SPi8QI0K6T9PdI/V+
5U+Rtu9zH9FXtV9+b1EM2It1h38FBukhl5NyFT2F1RiDBnB5L/hgRfdvNcx3lAs6flYERiubiBo+
AreblzE4DKa3m4WQd0vDaQ67rg1/qFqr50xXbuexn7U9qFHXFvNgi3sCp9jBfzswxKStqwcN2Avq
6dr4Y55owS86QmXyztb28HLkqiiTstxMdZP8JeQT/uJBQQrUBas35Ildqg1wIxR9CrFNPigjLZFG
gDgKQy35Z+KqCAqfX5Yrv2UaS3TVCk6yCnYAsYnEJ7/TsNyPI1a/ftaxPFH22MXWFVx7yeur3+4H
wJA7W4Oat06/GcQ+WLy4z4bYRKhAX6mL4vwTh90zc5rEBpmFVJcaZO8sUiuL9xda+MkYdQ/j6zMb
/yvBYXMJcGQDuQ3lFY/cHnLstZu6i/R1ovGAZoPOgeQUPoFwm+1dirZUJbJVELkMTFP2jlFKhRvt
IOTBscjbaqyHjdc6cOgM/e743rOw7mmVPf4RglUqbC6sA/f0jDWRT68BxJ9hHCf7xB4OvaXK7eeW
7ELGCB1MqqTfDChopqyAM6Gnlv4u1aPvDcaHtmIMv1GL6oE3gOEOr3OR8qslGLRdeWKOM9V/W47K
zAWW1EPfXRjQ1ip7wn11FGMOuTSinEBnhekAvLqumwVpwmgWnR4VTJtAokEuMSDfls6SaOgQrmaT
whYPrsCLEytim8llV3T/D67GwaIEygwAJNWcIQ+Mb+HL8vet+dIq8ETTVeVLSkAz8Mm+eRKnzEcI
5X1IJs+lhOCBYY8vXT6Jk3rXSoJE/jV+hQCYG0OiQ5Jwoh7DFaiE3nZw48bccOfbt8BZq626MaNh
94St4p6uyvmcwRRmhatG/Hp0YDS1s7veNPou2xaIJLmb7QaNZmOCMEUFIjQzm1ZXgpcw/U50DTNG
BxZXcJX9eJlcXrrxXH6GpG+PjhsVf6VQKYHn5wHipY/6+23uszRQAuq0rlieJmZdPLM8zPyMUXNE
2TKeQ5XT23/PUDjvk0Csq3UY1l76fTxfHu8rIdA4XJXYWOu+/5wnAoz/mX/hVewXkENRyJGiCB4m
y1oWSEdWQ8tnIVwd8yTjU8s2jYL1vnLwOEUW9BfBqAQj6sgjg1vZTwKy6iTbqPIG9Pxjxs7SKYlc
xlLj5+Anu2otFfd7TXK5nPfb/kH2LsVQ9zi02cXbxKVKDzZkk03LmkT8tLNFte1mvi2TXs23BBCM
2+LOe9vxbb0+41H7ijHLKEx6vXMfZWNg4lCdExbweINCyZFX11MdvuZ0gVdwDT6anvZLn29iDidf
z5D9nIYy9mISwe5rWILf7LYunzeBLTDZYViOtxK9OkPM5O22FoRMUaiFjtiKwOzgh2dwpuw+fTJ9
oOSVTlSuElI//k4P3nzte6wHnCJBdRFgUxE1ha9aORu5H3PNFiJeQEx5PTMwKxjV7UPnG7vE+jBZ
xyuFEKGm1qktrnhtiWtVl6vUH/eWil5Mlp0rv67piGE7c+AVIrxNzuXHcMFbt1qCVZzn1ucvBHn3
qBhf7YLdnL4IIlcLskljt7c8//ktbzKQlhZucLi9sQkSVzFV7nO40AyJd4tHzvAbzaXusHuOvP+c
MRYrluko6pBaSiOqKNq2uxSH065XwGTQfsZyh5SsDWPotQbZFMVZ8Ogg5FD+yHi0/C9pZGNSgDM2
Sf1n/xB5eCQmo9PuBVciLRN0NSjhchvAgvS4YVoNaOhxwBjygtr7JHqGc3c7kZgSODNsGEHQSszV
sVRVy9oe/hxz6tCs2M1JiSXIoDBF+roctYCaA0IVscf/qFOkTn9FkEC2f98mCdKXLVNT+b96/L4B
hZSTKgHqwSEz13bJv8MchCtlnDYL391VWVLQBksoJjqh19U63VI2IUWJKacZ0V3TW43VocMgNANK
Yz/pDiQ5z02b00oISZC5niq8Eto1dw3c+kE0Xsjwxom0HQ0Fudh3tv0t1kea9qaFednSiPIScxVv
bq8qxBoBh4OnNBe06UgNSp5E0Zr1RADDvjDPRMnQF5ZeHllZk1VtX9DLpFSelXEPP6Ist6sbG01L
34VqKOx7kxCuqPF0PNcaQbUvryj+K4eLrDxeLKimg8LFEzfxBedAp67dEsCwH5WDn8sYfTn7wObE
ViYX5z9IOsGWoVTXd1h7NhIs9pu65dT51c3A+rDNGZHEuTF7QuqAAPz2JRZKmKmpPJitH7De7SKg
RorqMTX5/MU4phrJMdB8TPwn9m3SJ/c4zEt99wbiup8tFoHCk7b+IIzr1bpJZo+hVBoeIM2eEJgw
fv/xxCwuR4bHDgH462yqfFF3Z8RWp06uRpisHnTfCSz5Pg+QYIUsn/er9YHkh5fbhopr4lVxM9nS
y40Sk21GcnJGHyHGsMXDbc3Ik3HTm9Rl/oybavEle/Hm+YcEnbzMyQhWSTJ3hcqyAXwAOBbmGb8Z
N7gDzvaP1Oh6QVfwMtH7QPSSiNlTrHuFCpYkXSp4nwNG0DWV2eU5TXQgnaSqGqwbFzkahTYyGlSo
ZmTh4quoQqPlWqKSII5gMl020HK8wS7mhV4eny/a0AIAEkq/D5PVeULqVTGwB0WVkusDMB8W/Qif
Er4L0xuFpG2DPfOx8geArzXnP9BhMmWIgKQNMSaGgu9t5qFj9/KyNpyyU4N8jV5at8uhP//BYHHQ
mkRCAPrEXhIG0PzZd3LjMcNHXkgCGT27NYHGp7Z8gjnAAwPxzSCEA0V0lPLxCKJxCcqPb0x8shj9
VrU3l6Xl/nyXOryHPomiAaQMuJrGGtmtJxHlx75kZeyWlFMWfhIoSjoSDz4JBRMH8IuKQVlRtt9f
wBM+Ter9vW271ZYy9dmtxrWQiXLxb2qbe9MEhS2NwJHiS2yrFC8T4XBjzMmSXcvoFV9NOb4rxyFg
O6cZvekg1JenHIwt2NMEGJWz9AREI8MSdjx9NsR/1Tf/AIW5LQ/hK4nhTVyrWr+x9rvdKxBvduFB
KHl4wUPJf8gsane5PTUzfEx7d0wT64wunqGEnFKaEiI4pLLkXWjxjL7tRNg1BijT0o1olDKqUBWd
zDFWfa8+3QXN2+I23IDfehsqExs9hColJmHN/XDQd0iG8HGedBskKp/JI7DksqBNf6IwR2TK7kXQ
ZqgrJsgPbVXHlI+YeQcxz+RIHgg1SCx3tjaVz7ZndTGYdokEUVAAOe8W7Hxd7NrcxBaJsrGZLAHG
xb7C+CgUUtH8VZ5gfUKHaUgBM/jepj3/qL4NTtflPhPUa8cbUMI53bwyqbr1iCzPp0Oh9JMKHcGQ
+TqrGwsl3pmGMcLdxcL3ptUn4gKzHB5IrN/oGGqIl0ih92jW/45N+uevRjHtC1rfe6i9YgrNrx5W
RyKB2/HnmY9g5tuXbpxDvAGDie10+sTQChYCBI8eDERJmPn8IeHPtWIN7QWyyqx206dvvmtOOE0i
M/uxKscVd1bxHMuMp39FGJXljEUcje/8i62wKozwSJq+cjILC5uG1O2cDAKLEnW0K3pCsJj/uyPP
aVXWMn1j/qLFehIcIVFDPFsNHv34pgBr67wjD7YHpcuMU/hUGF/ibHsvSexSK667HZsEES4jDglN
2iiEmBHpV8ZfFg1oWZar5KA8476PO8nfnqAbqDQxnlbx/AY9OT7/T39za37UMuVc6zGYdl+05yUD
nVXUqYTPDTpuO0D1PSNKEicKkDdWKM4cbsumSS8UbEwwFDgkAnM8alIu76A4pPhyCMFBTF87/a72
fqLkL+SemBgfmMAwy8sQRET6mNa3SJhVI0HZwKIs5z/cPJwqy3H1l9eWdkevZ09tJqkEpz/vS2jg
7nWU1sJtduw2ESb3pvZnZyOrl0DxmGLykI+jZ22F2giGJGTP0/gru25qbkZkk5GX9GYAhaa07ykE
UZbFv+FLAGxqTdDVdrTtvEAHwH6pzDoeHsNMErmnmmdx9pjU9wmXCwbxTyq1xkSJ3OyYac8+jDnU
mLnXkXJVT9nwujPrZcCaqfyGZLbxJy9ibDKjXNREnsnbvzM/1rlnxLGNTCRzmdmBIGl5FNg+8m3I
JqC7mlw+RWP4M2DqbC5qEovPN78G6i2alLqYVRPIM0zt7GrnJS25HlzXCZ7gPdTex8/9E4Mb8h+r
X1sTP51+yehCVKMVioKlwcVnpEQFNd9O52djh64OGVWuvPzSbCHGGXtTofZYBXBTejrCrcJutkAP
lDXom8aPv5iJ2eHCEiNjz8+ApNS8jFZUzNFFqfSDFrSiF61Fqrusm198SUum9J0RwMez0sMG1Vkx
3ONa6u949EIEXiyh5Q4EOE4+z1ciDyEl6qas7cG0XA9hIj5DGt5ryccwzb862B1lrZEYwVApF7/d
ajp0VY2X7UOlaVOZo/4pnvk1yot/TKyjNe3ByS7NtYad9236ahwDQfYoZM3AW8pEiIZXzU7IWao4
x5qT8WmcQVIcsT1oah/JYQEbNyqv9FIU55ybQo9X5hPFrnEevXax7UyjnkxNhwq/ZNbo91Z18p5v
grRngqw/ZIa2J/9bS48s7iRjbjDUiqgB7o5KV+b67Tf61CAIq2umHCxuacmBqdaWoCnQ3ASSjYJk
J7+XN47D7widSgbVYxi6O70DRJE24ewHeFZc0e9eF5wqaAgqR7pMWBYogNSB9L2KvruIXs/8Gmsg
P4Kqcx+U2cb6U/8XbDdHCWDLtaQzIJ+9a0xRa6b1BYhJyaIaTlmRcke2HcnPpg0gtdvAz4cauMtG
YeJE60EJLvek8pl8WTRGaurjfhSBT50HxdfZV8gTmb34NFY6mTpf3a7pRKIsJ+1bfPQ+3a+T/J8O
fScUl6BGiyA7b9xs7W6giJKdxjEDJCggf30ddwdArPMW1iKtlfaB+3pWp3boBmbHPXutLZx13c5Q
x9NpSbdsIYCatj8etryJn89w4Nu3vvifQQJJ7TBLtKXgzMWnvprs1CFSJoypTFiRtUBo5UPwyUNV
WMSrDmd/cr7tUvz4b9g0TVMBGqf1cxhimznKcI4atOERWdnyaGZpp3VWwlH8U326gNDWVogsrRyg
qFGbogCwe5mHmRi16aJR2Ar/Mm+r0LYocYbU1J2QFZ9apK31HIWNGexVpQKIcUy6/eqGMKr0EMmt
F4gwYRrufO5N+2TvGu3Uj4LGzOByywBu1jxyAgF1JgW8eaUqgcjXCxwJ4AVdghJjUiCK5FoYq8ij
zAVLwlLkNxZlp98CRZys0mWVLBB+LXlgc197+cJNuuduOPgXyQMXtaHmedQMI2ldV5s0H53nH9kN
wbvrsIIz9v0qpsSva8qBO2zEbDdFsbcIUPEz4gYhGAY5fLZ4DgaUOfX2rLv2HYy1tCCtNrN0t9ni
uf5LZW8eNfr1H7q2/1UtCerM5RxHjYYE8w40P6lEt1L08Xk7Zgb3MkCkVPIgLndn3U5iCPc3wva+
mUW7OLN++NYbgCaTqXnsfhQjeOINviAeMV5K0h1UzXhjxrEEWDUVtkQd0U3W2xwVAOEazCH3UwAS
yzezkyCJCbKRnx9lW5oNmzlCPPpWduH+M/tD4kAOH3OgHcnqzxJ1I72GI8cMZ0+v5bwS0cco/mS4
5bN4zNpS4WVh4D88dcQyJDnrXCi3RM1DL6qwHNw6F+ruP9ZNXuobOIVuFc4FTxNrzv58kLxKjjVU
BuataGCxVdZ7NeTGTF+YTiCAuN8/YE2JENbp+rwR2qJd+t03D9E5H8OitYFK1B5vM0D88jeOR0AX
vGAA6XGhAHMaH3FwOTDxnxnVY15RItznjTyBIJnDVYNz9GMMA2DEnlN0r44A1hQDQtoDB4u7x9e8
nAr/MJe6GcSkBvLD0H4Ky+nMj303CDfScUMpHG2f6xplQ1T5E6H2q0MrIreW4WyZcBtL4M2QAJOn
vim3Cl3kxY1SB3f+MgeV9NddLJY+4zBnxn/nhvKWJ/X4vi85DHdikifCLon+M3g1kL3Xv16zBz1j
TJp8a9jjIHDG2sdH98PbIco7hUJSUstn1yEM218ldUI9ff+Kl7VQRuzwwbktVaS5L2OdnQ5/76ZJ
AbMNgZhZTfrmmpcTWuAabbtoBcUY8FUbVSsp2lpbTAZm0O9Ut7fjqHIJ37dNMSB8aTViKumuxKuG
53xf7aR+8ZB/+tAZ0z3cwzkvDs3GRFeqnqiwckOQrfuHH1KysOh7brN9e3C4MiEinopE9wm+kehb
5SdcXpvTgLk/nVHBA0jy8gm7oOnEYwccywx+d3EY3NUzg7iHRRtGtQnnhc2p/Zk5DqZwKpHdOAJi
ZzXTXMX2ywss2gGB6DvGOxTgFwDVbJ9R/HtKOfGP7njSMdkXPz0BCrR40CEDr2MC0oCuF5CHWCen
x9IkfZ15JPScmZ4q8mO7Ul7B1roNUqJme8QQZk/lKG/ukySfumXKPo9G3j3lx8DNzbLrml9Zif6J
2KIQQNrY6Mrjkv1uogn+l+6EwdbVAKNU8feZCJdZgeE0nts9j70YfnsAsIOR26RM+8Vkf1rTDA65
UR9MRUbR2UNI7d4YaVY5t/EIza8/AevHDRtvdPJNCjOyEDo7WQ7Sn153r2lXBk8qWFGP62eu57aD
cEvOvgFX7EqL6c7VXCY3CRZwkANcc1ihrtQhGGq58pdboEgZoCuCaVbrxMqiByHqtw+uyvGHGEmd
KPE4/AhoESbvFCmUqqDHfzcDLnbFxzHryxF8MbqzriQ0qXwhXa6IRrzPt3ReU0CzmEzPuJsNY+0h
0forrRJqEGKhqFOf4DmfrXjn6lPGz6pndMOfGf0m4YuHy3UmxAOG1jg3dkEBTY71RabNAbrVeqrV
wxu37ojv7S6M5D4HXZwZJZb2pHMYWV1Hb+pec5iqlKMDKsYpPCY9WvgEPtjEUMOMxCbK7U4D/6XY
ZugWADZX+3yAJgI303WyvdK4hFqDgI3xOAmjz3Mk5LY26fQkctl1OEJEUd+YbwaQRQ9ULUcjRrug
N3lgDptY/wFWSTFel85x6qQCarYDQ/Oe6jvmeeuJJJIdv+PcJ9qjwIVMm3IZsc0ioO1h4a+v4MTU
jfgLtxWTld+UeEyfwCjAPfc04PVZuQczXuIMvhO8vmKXEd0/Ch03UvXGc7Kfv0DfxXfTWh1tXuMR
iujmN3pbnirxfGCDp46PRLSTzad9f0P9eEF71O9NZbQ+JNgoJV7afLy2EA0a2BXWK2G+spnTQgZZ
gKOm2AowFjhYbqS5p/rtZA4RZddEyFNimVYare2i9nVIL/bhHPVQ4byAsgXUotjhzOzlvK1mKMpG
lpsq57izbEu+1tJ9A9ZpqUxwMCN99+zvQGiAVWLbVJOwxofofqjnN0FACn49DKaSrUuVTetiKlIT
ifuKKx25qzZreNuCcXNybptc7HSmoZQD2uxPY41DnHo17W8fyMIgN0FUTBua0XHmoae6/LtNY5LC
oxuaV97y5EHpPdG/Av4je53ghNhY4b8Z6SpaVEzMiBXEDXda+SyqA/jTSRrGzUzll9H2RwFMPW4w
mX6opZ6IBvJ7o0Ip/2FpCA5BZqQaezz7ijCSmH6JhTgY/BY2fNDqgG3Wod3JVzcyxD6onSAZyiJx
jgttEOrJ2PWfMEARBbZYB5u8x0foDhlYL07J8klV03ds60/BR53ONKg/g4bbnVqEq/ae1v7u5qlf
AAiJkF0K7967w38giy8V5MCwzoEcZfxNEc36a13bd4jeeG/xOUWv/OAx6uPwakX+eHWT2GWi9JJ2
ke5RUlICsna1JNQv2fo29ZLEDMd/yu0HSb5tlcsmDwi2jFvuKj9m4zn2gbRkjGaIzZqXkdaF+50d
gCkIKkd9tXkPzYZefS2kgxuD0/asYUcUKB0PwpK3wENVAx39AFDDDz/nqpNISvZRGUBQmUCNWcQW
f8xGrEbo3ckq18DRzuSHNdqaVlYrwKEdON44/QJkuv+w5FUcF4Hyz1BDQyPOnep+VEF6rKCcsmwV
BaC4yuLV4ggXsRv1/mGNIJ/XwBd48lMfPfekvoQ1M9zoZkg4mQqrU4d/1lepEolqM81BtgTIEMzT
BKFpkIE5Vyh3z0xF1dfx2/FAn6HImiQi7PmStgJYmDgf+cgsWih5Hj7mmkygD0x6jRfTj7JFNyP1
IMrIig6FH1AYHar1NlLBRfJPg32Q9bVe/Zf8QadIRc9/JkMjIj/k1oz1MEAychtw/psTJ+oGBzLY
UynvscBgbn24zJCYII7eKt84cIqRv+uxJH6gC/qy4hY6/zxg5yKu9WJ4+WvkVkGxDkthF5LHSpXi
l294kjji+JBhBKTZvtq7Rzjqj4sw6HP7Tf6cenC/36PhJWbOhcL4GE4dxynji9CxYyzbanXbArf+
6Bn1/NrorOhTfoLX2VXg8ioJeddJC4skv79e9TxneJsHMFKI36oSYNfDEbUxjhdC28c9Xt0xcfSL
OIXqZFsnLqFuDYT4kEjP4cFbCKFpimJHsqV2LMLRbXy6x0bAtu/cBYrIutpVeFwNxStAXSZWNg/n
G9yoiasrSlpr27Q5/cGS+PGN4PD6KPXLSCCavZmSykuZ2qRCJ1orSPpUCHbbDTGo0F/NJ4g4L0ah
3Zcs9+DnhRNv0I1B5jqEgaF9i4JPG8TbjjS1kEELXGhZq72MSbj+I0Kn6z1c2j9yYz+7yN/dkJ0g
IJr7kkUYYjjdk9wb/RVUlJEgICO2rrxmQcuGTi+JmYcqH6jiCHg3fkjYJ7UigizeQ5VYSivYJAzw
Ra8VBilF5xcX+xNpGvh4QKJw1ENY0KiVqQqUTD+N/b92Ia1+/55l4qI+tH00uHmikmW7m/PDhS2T
qY/qZeSr8a6K4vhJJG2Wn82R/1FskprXI0u3JY/nn+4pX957WlXaxzz8MQ0uNJVUIU9ldlSGhokf
4CVjWyZ9dtWxYwOumzOeOxbBOHaSCb3Rph3vSgkdQr6YazNS1GuE8TjAGGrfP3Vy0w+3wvFnesMQ
loEGm+n8/dMc7k2s5KS7O1lsrTDj4nIlWLlt6S9ujN4uu2GJs0XNuWr67hq1GQfNsCxLNtXrUUhV
pbjNLRHmtHmYvfznZizEQ6swJ3Ae2u6UQpmvenaGBAzM676XgJn5bWuIXijovu/HNIHVbNDZp2mu
1iZEuyedMUAhbTdyVPliDldnDd7rHkAfYUB43lYAYmCMrW4DBlCC706wuMNAohbaWfIQyfWrIP3+
NYDfpZeVYhe0QDa8sJvCMxfadwaRE/X9E+srZNjHEQNzOW4RsVFbyIxUZ3HcBTJ/lwXWzvO5/TLu
LUAkhLi96/PSKv1uAO+MCyXugCpSEgrvcDlESJIXvrEzfHIbE6KIBIIbGT73orCzOq+ZTHtcMfhd
gwSC5ZMzE5RToYmRz49oTQIwFYx0rCHuPD1mIACs8yZo7soSPEtUM5669YlCIcg1f3B+7y4W+/9H
HtqvjoQF4OBbaQd0NEJRUIlB6us6GQfQfVvYu2mb1pZF4N3178QZvhBx2Env9zzQwdaGC69yTfBE
3JwO3y0rkWZE9Tf9Tr+xbEh5xCrYYC4xtFN6or4rJ+OD7pqID8qQtx8S4pmAQ2QU809pcyfUma0L
uOBjdFRthfpYOPRveiqG0pB87UFX4zHFeECqPHqWGX1UWOiTBsu7uYrFFp4ky8OTYg/255mOPaSG
kQvaQJ+E2I9y5psYwKC4zPXIBX2zTjoSrQlDRPI0MjWwwwkOOmCtUb6QcEOzMr1i0ZTcIva7R67c
GYdW7lNTQK2ay990oels+uQN92aYewDzbnr7p3HYugGX0RLrH9/Rsffr0umJYFLxufWHXLBXU8r0
q4BuCTCH7GYT4iRGYsNkaNhNBtQibkqPcSZ0homgDdWs5bGLMgJ901C7a7i7SaQKyUjOfSBhbHxk
KwfhgdI2JE9Gh+s2E5s3I9bH3vOVzXY/mduoaAbX4oNYFfG1FOT8lXf5/EzCxRHH0mvjL37sL3WM
c5x0iCSHv96WPrTHIgRLM/BUTzPbdVRgXX3fQrskb9in2Pwvv7DqT11jCU7uOxpDrUIidx6nFLBb
LbiuK3+lkyljZwgWxMOU/Qg04EDaUMd3898FFu4rNt4ZnFpHFMaOOvOwEdVq7fDtvXFIVNEAh3Sq
xdPfHF1wKRIoErP5SFuYMBsKXm2acSG1nuxwSmTRPd1As9d+LS8DTSodN0NaE+P5LHJNz63SSAN1
MR6qPWuj7FZyRe/8ZIuKMeleP2N9Yt7KHFWr+wNj6KUqi71WS8tEGPw5PFnri0C44o9+fX1EjI/O
oYugunBlXmOoHDnGy3XBCHJzBoDTceGKYO+Mc51xbdAIqvS8ZvMgguK+nhIxSuGsiqUPgZHSt/xE
WZmLzVh6/QgIFfPqdqSQYJLA5AbBT+qUo13gSW2Aogc2zVeVAi5esdIvvvty2tzAaVFp4VROFr9y
jnq1QpyewwkxShAl7qpUcIM1KAAXf3MfEdQx4arvPwKrztx432c7MD30MjV2ahr6HXR0qYE6ky87
+ou8ivhaZD7iOpZ62DZ6rBwom5lCAXVgLoZroq0bJ6CF/3xVOB5aGQnAMPBki3IaIfsjB3hdfPIC
qOmKGKu8D3VPrwWk0sU9TEoliDDwV5y2wYdHlwMlaNkemmsxCfoTqeU0Kr1p5DNDVFwJrHGCC96u
FvQZZ1GKrD69S672wnjRf40iQ+kQYF84ZX9XXaFs4MM88bHlEXUYc862hbxEvUYK46e3QwhjdgMr
vjhw9ZtgaQkEbvSG7M2pOgYA9DD+mgTlZ+ZHPZ1hlnfbh+6PpD1hXsZA+HoLo+Bk6wDB4tXExkaV
bBntNzsCso/LkyGjantXHxJACdT9F59M09Tdc87ox+iaVpR7AdbXB6iB2hj+mMEyX2mDUhkILPeV
c1ys762V0Mh5E1xzLFxZW6a22rfmNXkeRt3QurnlHh4zsAWYNCr7tC4PoNMg4RPN6DmWbiISC6LG
BlVt8nKxEWxeCkNyEp7asTydQ7ZQdYDnm6H2EAWyhZa4Pu0Ss2qFDZNq6/vo5ayvsGNy8C4g27AH
fkEBkLvwMGHHhxqUOvYNRsWyD702Biw1E4z9BsoDY4bDQAeCqHcva5UCXGEbvWnNNx1F/CYWXYaK
PjXLLl85yihWHr/Rw1xyltnTXazrgy4V7MJ36UJX4y/58q4wH92ERa12Gnxpi4HuKuyKygH2kxtH
cJstSi3jaC+ClOVRni0MzjP7gvmupySwJrhu/cgkF5HBEmT4XGOZa0ONNbn2sSlR0GNwnmkPRV0/
triCNgsQehJOLv4ZQNOEA2H3HhAqcntbUGwlgtOcgHt6I9RLFr9PmavL6LdJtnNajm4TtezL9D7b
/obt3UdUhivFflJB1uOO+aGUgxjLjS0ZerNhqrtEQo2i0NO+9sP2td4zr6Q7pdKPTdx/5a+TmhnT
bUJ70NOItAt/DCRIZtIcK3ibYFOoIhJUiWAgGhezBioGzhk7mSc/grH/oSCCJYkDqSlsEaHNV69D
V8PFRoSgNek7aK18NGoj76qJjIouzFkUdgDJ+6n/eUMTo7Vz5Jot8fcnnft0F5tvKFV7R9Xbpqh+
F+IEbIO6pcJ/UsAOT7mtCeRU+xX7MxcPvdQfNbbnmpSI+m4vAfkDbGIS0rpzSrpgUXMLwrGUWRsk
zZYS7dKil+PbH7IMZoGU6xIUvN/s7s5hwDPp5Z+P8Si1UPP/RpG6HvDRurRfudAfGezXqoRbbWLW
+d363fA3rDmjQg2iSVrW/O+FRPT28q9zoySsp/Jogisxtu5fp4BjnthIkvTV08gyRK6yySLMGsoF
TIoJfMteGqY2+UKFo7VbIa4DXJ1OmiOIscYDv9dFGqo6A8pLdRte+dTjS6xljeWZLZT9ZWyWVdsg
SUeTra7QTzceZjPuc8+xgCEutK2ZLR/3LLcXk27B4wrmq3GK6FvV/FyEb9y5TsyfAVA9Tw2/RL+T
LcXIat4WEWHt1NjPEZablnpIlHWHZQtLUyW+6j/1WXBtlHsjWyxW38Owo0dv9X2O6MwPTWVYS+9P
H1PyNufM/7/AZyBzRem9zelMAHXX60P/nu2u1KbeW+53fmsXh9zhdIXA0pzzEPXqPpzL/S79ZqXb
pqgAKfaD0GM+LcHBzzkY4zPJrGhOWZ6exO25ICicTlSdzKT6lO08dTbJU5h/2Gq5INwhWYMRvQZc
BRw/zTJNoXlS83lgoU1KuU+Iroo1hIa3KpBrO+siUTKmk3g3KbzT7vP8ZPWPtIi6P5UMQHZuUM6n
vIsn4o79WOXn46eSzXDX2jiGWvzSiuZkXobfAcLVLyxUmsnRilIZ0yeP7LVYDPqSsZBoN1kGsFBg
cLGQ+ffAmO9YoyMzy2cPAe4GS/qIFrgT8weBtYBH5IFeZmITsOOXRXohYMvoNkaUFMOhm5muCOy2
4+EfGdWcWZ9WcNqZl05C6V8bjcpjjos3P/3IrtbQy2mDRnJNl94rgpSQ10sQFBjYzDv2rYctsbwG
S/lB3WOgEWkb9kLR5i4zpnIaaRvGG7KXqhBxIt2UM8vId251C5fgf3emfPDGHTINxJ7ozfWGS+x/
QEKl0AjW2izh/6dCfemWih/RvFR5FHCZmpMQHt6ninZy+3CSAMtpVfNbo2u02Cd1nMbHPVP1BrUe
L/MNiVNOVyrkCEI8G0WtXbQ3RHDMPLCByIDr+QTeP9PFnoENZnj+0rr4HnztC01TKSt+G4sfY1Yw
EifwMI+uW7LGRizfukwDMCXbKVu32CmRTh9dpEtEyWSooSQY4v6IoJRqux74wCfmNvHCLxMIBibM
Y/sxIII+E7P6oTuC8ceqVxG/CKdbOh3bIXItosyGTi54/7dt0hxEnTOblTQaadYhj0i3GK5Gee50
7N+nbLW2Rz9ZMLP9OvyaWLNWoovCDTTjSXYetlb94c01+cTtEYrhcLyaQ3LgkZAG6IYEOBk3DDHF
cC2BBm9YnbLCHtONhPV8Jc2rNUJe6evBJ5mnGhM7wL/K2Vj5xWK4VOeiUZWspGzkkLRGAWkIGFSC
B4CVsGXowe0wDvt0S/NzWpgjF1i0kgEG+mWr7FargohWueyjowRDYcw6+y/e8/PSerwbu9FPu3Qe
pQl6265vgZpCsqa0Cpjm2rwD0gsTkRAKc4YEJ6hPMO6l+z2ftZSHdZKOXkbM7H3AqvL4Dt2orRxz
SNLZ1V51uVMkh6st+6VryXmg2ZTwtPERjEB7NIEyOmYu099BDm64vDpcoGSiZmDDvPV08VYbV5GF
4Vif1ESigDOE4wANp4NYaCJ5btqPYcDHoxBDdSFklJydbsf8VH81GR4zOWDJxwUSJUNYI/0EjAeS
cMrY5r9bdCH8W0IRyRxg0pzgqI7KIBGJCb2Qlju7V8F3Y4aGnATbWNAW8qpTGjyRYLSMQStFsy90
04ugnn1+zSlXQFtypJK/YiyOkdgAwDJywJqbOx9VcF/5yn3dkkOFcd2qeWhauSi1fJKtebKY0dbt
d3LvYv/ls1nYGfj/Uqp5HLVWC1fruca0EH0Zqe2r6OLeh4bkaRUZ1HR+VYz0B0jdSP2KX7w2lJnu
6k73o1vTGxoBfRRWyGQMSAUHlYcZST9pWuAxudxJJpeccQrBTgKU0HhUagCT3fsK3vWv63a+xaaW
ioyrrYVPPW9U9sF9mpcM7xiCpzkqumIflhXq1YeKDDso8Kn3es/VXwqoDJRUr+IjQvJUyG49gQhL
tDwZd4LKWpf96XARSrUGXXZE9Fb9SaRmhV1aQ3TDatvrHCJnm/62ds6RG/cCp3PQz4OXgzR8SZcB
K3d8uBzp979r4U5sXP73uBoAl9M5YjZGpYNS7w0h4CUXATwWm4GvfUKMcvv303bsDQvy+o38wFfv
fij5m5yy+JPfYmOwXveWH8FYCu3PApU8wiLepWgIsf7j9W5zO7YjLFU+9k8d0tBiw6bnlGxuJ8AE
4A0ubGZqIl6ClzpB6+aDJXxQuu34LqZ5qA1jRdH+RnJeT4hQAerTbKpYn7SQPrk0xK/g9xf+jffU
ZlZTofvTm1vCmzeY16L2sT5u6MJVOEx1Ty5qqu263uaSzHoDVWAURJB4vsDYU/y5xRGnWNyE6Nt/
OxSPu2kahjLjFwfC4XjmD5fVsgB9vDP2XF01NiPAawVA/S1SxS98k14qZ0dAhiGJD/p0w/yIMPMv
O/8+rq8Z2aVY8hVaQM4qUq0YaT0dXfIT21IqLAiYEU7R+zCh9bb2d6MFRcLPYHUtn4CTZkgWSkQG
+JtE6naqLLdhzbAxP4EQD+zC+1/p6Nsy9Fc9JhWILqylwU+ixS8DC/0WsbiJzEjntMR5mR7/bcSx
Y28N8LjcQ1YKi2j3Jur5zaIpKQLGM4DeJgfIv8u8jqT8uS3nE1VHp5TtspEN9brE+CtQqiBM0vpd
ZLMJ7BlR7clEivjXwfUrOCwiSbIGz98tpjWEwrw7l4AK/31T0Gz7my8Kcp3UB6cqn0yar7FIR2B0
xmBMp0hWEXqH31T42PSMBZ7b2EStVr10qVEJd5h3DmseEojA2psk5NC4eWOKl4XCGSoJlWIc2K3o
irYggsnRzAnaHGGoibj1RPxuIBMw6OuHTl9Hk28w5ZTyfbONa6sYf9hl/3n96vSPgpbO7W+6XhZ5
hdK+oZh92Md9wmuKSpfy+FhBxpIPNb+iLKatTddH+WCAtp4nokPA5e6aEcv4ofHuC7X685E+sgkQ
BnQKOFigmVXvLVETyw9KvQxg/lEV2FUCKoMGtxky4KB6Rwpkn7+vHMyLWsWVbLN/ZMoM1RUUrKIf
+pHXllT4VSaYgTr7/4YHX3uHnQHA+3Uw9hpNKO9z3CNUhgOwCIGixbwYWqjdhS4s5v3Efivnx59M
XbVg/6uNYoK4gJ9pOJaS1WawMS6ueVgK6Dt3ySGmYkJ6C9OWqxETu2L5dVWdTTBoIEmD+W+PIVRH
CAGr4UAFJUraeY2XVFWUjQXznLai8/cr3KlCu/VqSx3pLaIiCYqf14DEHt8FqbTv8hzO4fnqraG3
FnyLaUn5gXNp/lbfQqO9dxxmXl4PcsKu0xEFG8u5l6i+DXx2auyQ/focEkYSOcvy5AVm3mJDPnBY
xo+sYXuZUx1PW4QhK7Sdfoau9tTon56D0kOCDjzkFKHmuDel6ig+GeUlxUZauD9XixzUULrwjs2w
k8KzR4AkvzL9f/DP47Tec3TV+bpZaJYmre6p1C0aTCbwjOv+erWPbRtB8NDuIzRW1z4pEjkuiVxP
1PSWuZwfFh2Wip2kW3a1t19oJ5kSyT04XsOqu6j9eeQ82OxoQGsz+kgABgp7cxywEFs4i/D0aBlI
mOGhnTJPUYXvtASMs9RtBfAwJOl0tdYV7f519vHTk1Q8huvcpaCUNw22OEUcTrZ/IGl9Cfx/OCzT
kPWm6qK5cmD1ug7GwQqK2pmC9eWLw4tv0czwQMm260qLfeWeunvNwdAH6jP3FvfSWRUvtrldt9MS
1SwMx8XIK1LmxXE2TlpoewgRn3KkuEEHnMYLf9N7WSnvLXYzsoGsic0JFqsYuWabl5S0kcb+2tLn
3X01EZTdkMGJgyNZSsLU7O0lR+PbOQ6C6BcwUdat0dVyGs+6cTrXlXvI9PYp3QcHe04uw9C7otvM
NROUQTEjcxApYQz6/4uZ5SrtZEk9fM+lur8KjrBcKgsTv5fkhrTaap18lHy4LqMugXvuPVrAOl7Q
YVofo2ViSRj38+hpuQ3+R66KTc2UII6nQvF/m3TYhqvkOoQegxhQZEzAIx8hTw2CH0quPrt0eN5f
6PU9S+9nkUnGIVUSNvlGXEx3AsdlfOY2agNDg03IUGS8xBOyR19F8X+yGnmtzJ3p2H4bNxmn1N+5
WfauLCvCCgxusqXmTM9N8//sbLuXtuSxuuaqsq5N176zw0iRa7GyzOhcqyk48ti1wS2pEXUd0xDC
RtZoTp1J+xU2XRCd6PB86csQrcIHXlZomS6WlLUgmOVP42pP2fMQaMY3r6CbLMsMMTEmPCOeWEVo
b1M5JwIWz0QFhyJC3Lm3u033X2TzMg5XdKrAN4+ZeFEEWSW2VJ6B23dQ+SrFj4f2Cg3yo8UEIiSU
aoXH/1XUd7xYPQC3IGDyjg8pVRlhThGIm7UoFPAwoVFCgfRnI2Ag/vRoNPVOH2MBL2Y0qlr5keya
mLsuAEzNP0D1wQA1C39yjfm5mZvnq3vDv8G5qA2oycRdP6eCCrq4drI95TgILPZLKXPyq4c9vKPk
/u0jPaQme8/z6//onyGyuA1x3tKFB0f0H1FQlQbd+jacNI8iOlYpexMe+DS0PcQp5JgBF+yUNn1Q
wQ3sc+2LAHVzTQ4bu3CEhXkYJ4dE6+8UbcTcnJIUHhPCnQ3EXjyAlk4GS8Sk8+0z4sfgiE7wt6fb
e5HPbexnLpLdZxia66URWm38ztycK6sQ9EYLriBtJaXUFi8RCG7Zg6aR3mtGh5MTHqXQGAJuBgf9
LScNR2YOAK1MIrVFLZEqFH6Vdgv51egipYcUcLas7Y1NW0N5DBW98+T86hXmSaIzlVfasWQel8Kq
7YFdejJ36KM51BuCpNkv6mCPcCcDEZMffUoOBpT6dHXpfJAbKRH05bwE12QZUjQXkxN4d1UIJl6b
wpPe7pvHTZ1IPa48CsShQcBQRCionA9yVBAneEv+6du0UGY679jjrhOcxxNf9phvhgpm712VZ3t7
GiuLw8Z4a8WuzEuJ6ktAAjlJtuk1VJ2HV2mhfJR5DfneL7oozCAeJwahi2C+p8yDX8Wvoq+XpDUF
Od2iiIKdJJLC+EmvJYh04xEcUHuvakPyVH591FRwf+yGLWCnXfGCGFaRz0Yam13dwvPqOZXBSAob
hcyX6YCGkyHnGQUIuwDYXZuRDZ8WnpMX7qRRNLfTQj56FZz6nkwb+Ea+J5DVqOEcOO3/sjS/JsTT
qQQqg03ygfvfFSTnYlEyd5sxFgI88KPCoatjcHze1celYG3Y2TLxp2WB6T+IJIvGU3+8URT6+Qqg
55QkgreDjOEJ+f+YKW0w+Ihv9511fTro0pH/Gua+dtmnjibwqL/N8sNR3ay4eHhJ1jneTxmmbg6O
zslJomWzZky3Cgkoy5UH7vrpfHb9yvzx8tNxFEg54ohbMa2YkuF0Hb4mbHAFSEv8qM+Y2EB+MANl
C0JbJlSclfT1aow9A4aza3aew3IhbecDkpNQ3KLgUxjyzu8PZX2gwFlEwtBSD8df3AD8dSpE99KP
pK2wtKGUYzqgr9OKrlqpFrkk+TNJZXJ9Wcu458jXLHu36bUp3qiNYbGeddx/VJRQHsikrvAVHror
sxRclNtoJix2EyEHbL7+kTd3ozzah5j1f/UXf4jiO+xGsRPZQUHA5zqzMJdgwZ/jDAZctqrORCbm
4sIGqpWK39IVhgvCK+pcChFuBHu/BOadoRo0ZmzcQ3x+92eyjlGrGdvGdG8+Vs5Mtx5FH2l3c4AR
0117NiEgzjxTezJAkNpUP7SiUVbBSqQ0YQySE+h/fvdxo415q8UIe5R56vUJ1mcp9CGfJRGvUdPx
7M7F3KkIRAierPs/pTCL4WLyZxfD3Lv3u+n0sFaHoJmblS5yjMBQBH5Fs85GqscZ+J8pPLuNy1+C
VOw75UYOVR/8EHlGEu7e5oWL72SPtIGETv5cttplDQeGz62PLkKNQ3EJOJUcqYLv9pF9E/GWVmUp
Cvv8SrnssWND7vgBYZ79CQFuq8ygCRB94BTBlXExu1eY7t1A89WG8zYieq20sRx3jMFl5/BAOyZS
KGvgnZoepzxAazHRZEm5sMgyCKoxTcmcbtHvkEvW2ZoWmjyTbFnGK5wOxklyJ5nocbzmaqecA56C
GhgnJhAbaT6CpcFjiCsYRAAU62B/B74+Sk+vpQftbkkjKRBmJ1vLZzYPKouZXzaKWdkSMPWi6s+i
3IlwrRnnahG8y9JDlulWDAtmuUsqIIos8m12ag6XSnCnfXdgactqpa13zikFelP9SN7wg+9Rlgk2
Ue0BPT0bNZtqdbadI9ZJ5OdFW8vKPFJ5O5hXB0QovFwrfAYnhuFXvHcDC4/ZRLynqgYGKRC3fxeF
0pDB6/XXo+W57U6J9zXgl4ToO9mjTUMm11AIBhykixQwAkXHkIr9Hps8OgYZVauLdptt8lKTA4h1
NqN2sH0QfF0JzWWbDgy5X2v4dr+Un2ra2w8+0kKKslpw8UMAGEpRt8LqTG/a72KlKUb9S7W1V+h8
n2/1l32fnEUPu8nsKrvx5pbNw6l6km4zfTPoX7YStvcM0LNJH6PJjhqSbdqu49OsVBQjoJMTCIRX
w3bAIDn6F1mutaNRKYUtNd8NH4ut+4V6VLg/+dHvcl0i6D9iyohscfxvbwDgsEy/LaPytXxpn5Z6
/SCISwx5ftGGzJ9T+9bn8KYYEfnBMLbUNailny0H11J7Wsh+wiBySr1detoaUC9Hp0RvDjwIDjNy
N/c87tOMXPdhYOioFRM/EVdIpmHVigmh7IHChJy/NA/BXexBAZw48JipwAhWsEhCixvq6edYzZ+o
+k7RVHgj4UnuCOdT2vp552KFbz61kZshumhy9mKYzSVdbRpvfo1hE+Q9keAcbxAj8qBUXwXxvk9s
o621Egfspd7eyLDbpH03Ebtw9dGUu9J8jT/7PLm8PnbnCQLSEK0CkjpZoVTJPGUB9+Py9XW61/sX
/e7wjJ3KHqX1APHi8iCKrMsc7mM9Y0m9KkDi4POTy5kNazlgyFW2OjEPVq3QFWYmhfQ3xvoawEhd
iGViNWxdcL9F0FMknTZFgwEZRLaE8DaUAPMhmsgrYjqlyKrTKZnSIt8npdydiADLXaqh2hI9Nzmz
dWwM4HkAbWCGd+Yzpl9IxZLqTMULXqCR66mFn7/sxSECMsmh2on4tbKb63Gf+6RR1SnKeVIlzmgo
ez3zzpJZ/JFX3hwQUzSCuAXAtz41u+iZTJgBmMW8b4/uyAXWFOaOjSouXF7vaFznjzqdKGhFa9bc
zSiqWuDEayW/X67qU2iwn2mHQDsLRG3W6c5vfuANciXcN79g6U4DvnVHihJlBBOEvk/pYMPcz00e
MrFFtgD8niw6PvUoolzGm5GCJTaT+P3e/avdXmIiJPc+kn7TlQnFqug00mSxpn03cG5dOCgko5UW
FhO5YwOppizHaq8hY8lcvmoMLzIyZpgnyyadg1rOP+xO65NXl5V3+Y59TM6BCgH13KmU0U8ByzX/
R+fubjEeHw98YP5eXsVQ7D5vnsfLiTm1vE8Ry4pH6e9mCv3pOZWEFqVes65HjArHdS4hLOyWlSf5
v1HSvdHr/LIe86UzN0pMTjJR+cvjX5hfatdRGcwVYo/NegJoQNN6U1Xbdw0EPrL3YWV2mnI7FfXI
/Skb9cG91JgLhkWexiVqIEyCyjYQk9zbdCn+Q7UwpSlZtP/WGK1LZEww0bKze11wwrSHZe+sqi/a
rTvSkjgtDIGJbXJYRAhloovrjP3udBUb/3uwVkmZIKwrvIPOvO34XTLoiaKIsKnl9pzgXbbQRQqV
ntz84eUHsjd7Ur/dscLAhQ3dXxiMHG9bMjFIYeFiM05v6juFEkJH8xPA+8fvo3MnGX6qdP+bTj1j
p0HNQebBTUhjBGLNu+406Uko5w4TXOF8LTdnt1yMlO/U76m6JWHtduwKoaKisXwzwr97UUkcrrPj
aDO4sOb1VGH/D7QrgyVhToasZjxOERHX+wdutZrsJSv1KTtdBViXitGZOi9oNn1ypKuDGrrvpr89
7sDmO7zjuZbOQQCuJbAB5RP3dkqMYtRY4oTAJFC1HNNvSiVWro7vh4P3nJQCB7rUZ56A8L8yFRsn
PAuVBtJhXrJk4sjbbPIV4CuTmeht7WB9tlJ49/sDAxy8FpkGl8YQFJ7OIYEZMCI86rxJquIlIYdw
K9aPvvqcc1IiAQnIy/UkiYuJbK8VMg8a7BOjQrSUifVEsrcdZjsU1LJS8UTeclfotoVwUebCeO6e
aPyCA7rm9VelXEM6Gvee+zSBGhf5pfaJteKBIGuO296UkP+X3QqC7Qck/cheAbOcQrUCPjidYiRt
9dDHbRZsQn8YLPbRI080IMlCGmzQzdbH2EJOklSpLWNUHU6JoStUTpLDFrJNoIWQ2qgjSxSSxz5y
yM5R65D5uPj6y76jKj0kchKNIfI/H1f50U61/IWUj7VPXFCPtrYhvZK22D6BTwn7sq0zQXopLUeu
cwa2Rz5B+n0+8grWRB7qUV2eBqKSB5yoNi0SYha4lJ4nDFD5PWHqL6UO/WJ5I0/dk+yxPIojsI0y
V67Tpc9kWhTSD6PEJbwTaZeLtk2s2tWRvhvEUnH9D7cScFSofpyWXWryxJMT2yeDw3gTzzpgBNho
ddpF385y1VfNW4VsiSLz6ZMYl+/JsMTFtiuZBo904Ks2xONAhJ/fjCQuyCOQePhIVG2o8FuRp50z
YmugKvumA6RqPPMIk88/lruG66vjihvTbZ2JcOwCnqEVmJJ7sG7rDTY9bHLzc8XRBTqZGAkAT6Ef
/dKuoI8MROPQK1Ux+R8FNthKZebHmSN7PGrQwNC186QNO/jOkeiNfMHhUryPi/f8AH/w+1bxLPDF
7ONcQZm8XpsLx4h/SEr77RAl41lCD4Bwhq5772D1UXcMyEyV35vQd22lV35zTgzYcqw8MpwNsETM
tVDGOV2qka1hyWMxQ5WywtnD68mT8Zw3Q8iBSqSYiB1AKINgP+86D89mYy4jO1uLptOHjVsjSRy+
0c1YgSfEbT/H/Kb85Umxfdj0/Oy18neYc66oMZcXz9geqiE55ixEnjfiFuUI+qwiizB+EfMO4xUm
jTfcP+sWRfCttFNWwdmrZixMRi7El/1YccsnMV6+szuVl6OUWRhpwKVFz77e6QbLQEzDQIwhcEL3
K04RH/lOXeu8y8c5FoWQdXQmBiZCX2tmSG+StPXkLGKDxPWpUhgf4Wa7rPJhDRJbocIE+37q8aps
3dzg3GcT22+C3hGl/8B5o0NYuRtMmbvkdWdBdm1+gdeU8fi0GTn3CLN2E1bItFpGZ8bbP6zKyTBk
zUBB8tMEYm1CplX29HyIlnT1nAeQZT+D+NgQswwX24XCuhEvTQBJ24uuDDIwkNZnSDZrQSNWT0E8
K+ekmHKmL9MCMGZJN/3seNLH0wxYIQN9PNxYz5uuAYt9MugbqZvZ3BqP/pk3FyFeODqKDMUqN7Vj
zGIwFaN9o0uENdag/wz85rDlOxyVzw2IfKKf1nSitRyxyg01Lc7dQrIC/RaM+8jB/NiFmwBBz4zq
os9Gp4U32Cf7AX0Aph4ziPwg31QWF1hAqyaUlQrbKOeOJJqc5axReBjwrvna1kfuE9Fk6RTgtV98
KibdUrKkAkJDJ/9uprhAXyRgbC1DJL9m1PZgyobuCUr3x8K75+/sYuLrVih9JzQFszntpZ8Pqk2y
zZDHTtGK8qEDml76L6ez36Pp5lvQLP5P86KGEeItcys7pwq77fAz8qdNLG4tT1mSM96IKA1SVHwl
T7+KyszTXogLG9EV3q/VsSVBha8rXtLj0qntuA2EI0w5dZWH0/2e+3cNOoaDst4CMib2Jo5eVkKN
prsfyL6eKOMztA4XdOA60kJBtaU4csbtppIaoWQvhW/eCmLIRR/+bn4NzBKV80yDPBjxHWaEewdQ
401lWM435mrNGGm8C0MDocxNdvQJv3ZMBSGbvBOBJnNF4sKGpCf9mkfgZDL1X+YFVsalIJnWeyG9
t/tjjge5OonopjAIOcCyMuFMyzAiW+mmacchMt+ueJBJWPSXO2mLbHGLSSQu97BA1sVuA8ZU1T6A
WuAuF3X//KjdvXHfwZypEKSMKhyvIUKvIwQHTGv5Pr9BlcuSVndTyqoRvnHp2nBhiKmOE9knTTlH
XSuxyTmz4TDeRse0bZexe53Aw3fJDftltB29IOMHH1P5LPnpKCJpm8pdhj4/AC948zz7vr2TYAjK
iM3+wOHXo0yxQJTj07zTAWWbLo2wuEK31JVUt5XHFvX4AQ6avTBR2eYiim63sxuzVDK0UJIsB1/J
EMZERZ3GeMFmFzDojV00DrLXL6/xC6/7lcOJFUIUSLpnQTqjqGPq/tquFvrPmtAC3mK6UuoO3j6j
kz6suBFuqYF9vhARSdWR8kA/mL0OHV4Z2Y45/2WQEsR/7gX55vhJI+SstJr8PcOHd6xOLW28ewjQ
h6QVOCxSDeq8VhPE0SlZXQsn4O5mV+vWy+YPAj3AVPLgqR26qD44OQmNi7rM0+YQC0PI+y5ud+f/
tu2E186njbxggxWtoLDRXgKlS7jrXaKjDk1vwiy+Wz9DrIoV0cG2/e50w6ed18rmm0MXRFs20nu1
mWPcQ7lCKjUPP65Um9P9pO6a17clQ5ksvWn5yRX6xmW/Kj1umol1+eAVZa2SdySaaJeSO+9dpMZj
IQiOoogWT6mop2jcBkaRlRKHle6kULPUa6JzHvn+TPrEFYZOZmx1MhqbR5oaveEngdygQDERcCYS
EUvTN4YWMXYetBHZm1tQnLBcYfSbJyk1FEAcSjFTo3X8FRcEyQRVEB30BG1mDtt/IO345k+tUzUu
1D4PBrY5rpY+VxwDeI8VFWj5rayIFZZz+MZOXgYHqwv+7OILsZ25ZKHkUSzKjkXEqYfbr7zLjT8s
Z2MD4zKG9tlfKpelAKDbd9aDfc+O0rmI6kXm9bkY6KfuEYUrst+K9EZ4Ssa0yTNE1SJMsB5ytH9Z
ovdFhcDzJe03TNUipn4X7qhaw3bXLNR2PmOd9iHkhGKW0L4lHkeTNDPiQaqHNLqT6WhVvU66dILD
rmC1v8aB2m21OjCQU6rn5sWhLzsZTj+kmyZR+6tgm1BeeVQhz8kONoILtbFZybkzAdpC3krkuODm
4Fq0kk8B34lSrJPRO/LvFm7DglRHNhmQ3OBWT80Lg3gzN8PwnhXQlhP+J0OrEBMM20FlPgaqmKG9
HYxPbTsqTNldq+9s93AoEt6n/DNmK3f+wXUi2kdRWdZ/ZO4XCnwmxU3kDZAVl6IkQjIM0nJOPt/8
S8WvdiOOrbz3Gxp6hv3/fGBR8l3mBwE1eK94PnL35Fn9hCYL7e6ONAFKkpXJOXW5eYmo90xwoHdB
WhyYVflLLiVD0gtr9mHBwZReixCukKlnh1tQ0XPUcyjmtMJoAZ6VCg21mcfLwScw2be/Bwsm7iDf
oyz38cnJUAt/W8/chs3nbMJZizVRGo+wkOQLOqY5/NNcwmCBb2Nr3SSOinylOjndurQcwG2VeNgL
L0OCwhluFqpNo/8ciuXV1VjnRww1NOS2vQPaHPrTEuUj/vxxUMaaJ01r3BQYlSpaKLd3PDIcygj4
KE4NV2hZChGo0ele1MQl2XbB3sbebIDUQTkhWlbe3E8MuuTu05CMTcJyZcx40i1tK9i/kPMqeywB
m7nTB1AbYRoZu2M8IClZh6TT+n3keOYt4U7y/y0aVhRX8cVP+fCijmHrA2GEyeYAsASWrmXI+wK2
jDxY5vkLFmyVCLyFYkgWOFriM23rBwW5gwjGkNkod8JhKllsyFozUJ9OgY8aULoYjUqGYLZq4HJG
OTZsJkfpbREA6iZLvlGtY1rd2d+18/6JBy/mfoJn+XjZnwdYAdRMuPLExnVfgb5zqt8o8za+djC9
wE1+74t/RemznYvw5Mmtl9b3b4GC9zuhBX7AAZoIBb0ldej+h9PhdhQKfhibZg8hoNwyPPgG1N4S
FGS0txv/9CyjkQVgHri4f4kTWj3ZYlelOQDxIT8z0Pwkh02TLgjdHXLVresm8VNJ/Fi+medo8/91
NAVdDYwTKZO6rSVgH4gquZjFDHcYnrBwS+sY8mylJUTnWHG5T1pc32qD3ZWqdFB7reVSlbGbbpqe
DldfQwklNfcQtPPgK+X/piOZYgx7FZE1sFdE+T5obKC4U3hV3wbOJX0qLajssqaOeznYmsWUW/XG
QSe4B1GBiXuf1IxHyaR+NpM57E7kO2m/AdTpQ0tn2GXKGSWXYUFEKNuOrSOt4gZ9LTnFRxe2tVOT
HnvDDjJ1qPGIo6MpATH2czmnqkVZIgMJt6/1ZeevzDon/BuXX0tv0kjruqym5PLkrEI1/Bk2bB0P
N2zSRTby6wsw0EKYRd6gpKkyJf7VuAa7kXVk7gJT8S3/lohI7U1bbZh69uFI7WbOzPU/JtxPREdz
VmkvtOP0LJF6THnkrWDLtdJQeRjzptX301H7co048mbywlm6cX4qjatAJlu3bNss7eTM87x7jrQG
Q0cDsczR9zTeV2O7z7WC1CvI6K/FDZ/Jqzq1XbsKhVXXaSxh0WzypXvZMT0dg6BTCqfBBWdvOryH
/tWCB1HivnjRkT45sc6B/emf7XA2Z+0W8tPGE0xRXOcs11zOjXvhyrWd+rShhc+8cKOUStadKwet
KxIrCG9WWLeMdpO50136zGVu05y12AdLo7Z5fPvuK29DztqExZ9p1EJCWDSqWJX3xY+NmiIHIMFa
bEYsUdJsPbxTuijx8XUmrpBJCw9l8ydahUBJ6IevrIjYd19rrJV5+QsZyvrn5rNLxuedFzWuoOMM
BnuS6BTpfUglGeaLw88hNGMaT6jT3bBvSNqM6f/R50NYSoyBIG12U/JmMU2PQrg4K0abAbL2I4Iv
GOqUCBa35SOifKsRL8yhI503/mICYbebML/uguGz7MTgK2hDPodVbU9BPV6sLR5dQfRlWxmVczAM
K/tozvAaxcuuh5HNxui0w20U9mZHRAK79GVUVg6kUOgJj5YBToNTPuHD4BJXZ55TO7QmF30cHlkp
RkIrkLVDNzNgO7tryapwxALf5L5a1tnEWRWJfSe6sPQw6Rhe6koz6ideq0Z3SjbnkZbCvEObS31F
Vm/YVc5gzDEnATJLJ0wAwPfxcIpoyhWHIKd39+vIEeh/I9/K6nYdH+kDOZBB6AR2Zw3bt8n+sQ9o
hYzuukzcM6vxFKeyaLpLErrQIsyxSs7W5RLo6aBDR2mmPICBW7Ztb9uhy3APYQaZCuZ8+yW/USAX
1DMniEQ02TjEf+Q35fjVY+ZI70TtyAVt12IutemToelzHiqeoUPBpgZCT4zb90W4fxnGOHjNxt9R
PBAC8h/UmWbrMDC7MLoF8ATaBrpjolY6uCXLkbyH6pcAjNkjjJE8i1EqdVOWr+SBu1asp231boUG
2FpYNyjqkvma2YkjQa00QZAN8hZaZvAtoSG1JMCHz9z3zYdYQby8Bm1+850gj9Ivkt7QLQIOTg+5
aJvbb/4uEORCWGI3bd2GpyFqPDPqRGTYNBGMQW/uZ4dfz01vPdVLQfW0YmyVdT0jfQQ9SAkDKIhO
nKCwL1T5t1H1bMgscwEAE8UWwT0q5Dk4vfBCdZtRTFXesO8nIUsiExVh8KPvrmy9PM1NrZTnrr8x
AQzMvCD7RVwWKSp87pu5zIklm8MjoPBMNjeWk0KHCUtRr6pPzrTPm9jq44AbAoll6RmgpIeCrSC8
aSG70wU7tQDvs/w224HDSNNtj1z51PWL29oqzMnlyWii6MnF+Uem9dUpa0j+1+UapCUhlPf4teK6
RXlAoEMiRhNGhyaX30qzQzANPv6U3oIcP845brJ8jOQ08Bwnnp37fu6g5hOkLGLfgv39051lCzxE
R4gchVm8mpjBFKeHQCSXCkwIbTh2TR1COH0hu9KMSSZeYjQv9UlHSpr7bIehvpfOuRiABz6gfbjO
h9WtF+62VlVJf7XpBuv6E3m7cPiXh4Z83h+YmR17PVghghfwpi0zqk1fWVxdhTOdNsjhjNWeEULx
lLv7pLpX6vxT6hwfvOfERU7hiVLcmX8UnDBj7SZl9BFCpv3+IbIxao/YyXH0p7EloiS0wuY0YMt/
vNsTIYzKTiDjFn+FGhNiXjNPSEacoif053i+mo8kH3UXumE6hNUo/TU73qAE0ioQP1w2pi1Lhm7b
qDqLDJdsrwI6c/pBGZu1EfFeIiVVz4RmajOMiZk0j6roXVuas2l3E/noRcQdniBuHZPZ+4ZlUeUN
IW8jr7bk/PP100svCdacKLFI12Mybb/7lF+amixV4e+A31zzPB8cUkd6f8pgCM/+VbiEng6GZcj+
uQg0oRr9Y6zge2v5EXVMM4Wl/HlbyKi3jtgLO2v/6g+nfkljxrpn9uU/QnGlkahhU4uYT2XfflSC
VrC0KUSHvRol6fKTrkjv4eW1fYFSGWX7B72VZUCsz7OzmGY4PK7F5ljwBRhGie0Sop5w3cstiYKx
tpHE19Js5JnwE03LRrsQLvtQ9ta/e+ZcHgzaTVrMknxsvZqPwEIzl86OqoHio5ea3BTLUjeT/18/
Hh8oQuxUBYaU92aXtiryV9i5hMkHhRm/VHYVrPoKrc4a7I+WjXlDfLbHANCh1ocxJhypLNe0tCZ9
GCvcB75f8STZzgc6iNYe0sZ5YIIFM61tsLyCCI3oRAClIqoxVbK9lhZdQZsYlTc1n7qS75QmsBHd
1mEZnBtH3cFJrAtV/Ki16pV5uUQ9LFJ3T5pcVf0XxtxBlJ+gAWkCrDneZNCbUr48sWaDa16mshLb
DKNRsq+pi2RzEBbmET2TrgvZbmUM23W3pArwmnrtL1kIzg5hecPMcug4jgHsMaz4ce5A44lhplIm
vlwd8vnmhRi3K8Wc3Oa3IFOjQfQ1kEjPc2gXd34YF2XcDE9t77eoL9w9sugopFhZe1vSx9a+GbP6
jQIcurTdtlRhGCftNe49bAx7ogQTZWZTwxnsYT5OhhwUA8pbfQ79Uwq0ThztOkP+RlA+GJfsIQrn
+jKuHAm4DNdz2clG+5Wx8zfNWGEOGicWBDrGfCpF43CeL8MQbnBRjAvupuIYaH0cv/H5zBKldzBi
YY0hcGld8Ctbpbs0TLc+ckVGfF5mTW+f1x4KsjWlGD/pEN1TpeHRdcGLNvdvkR00carr6WuKSYLd
R7SW/jint6rwJzItJkl+nl6dj4q43mNE/eMt8q8NCpbJAMUzd/wG6g4VEafbcvAZrTtM+bz16ihK
vYJxbYdTnqBGDPcKnIJ266nKFnC04XJfd6f5QaUwN+DK1qVFVmo1ydoUFdm0OsiAp8I5OxEWKVpN
A7Y4H0R7fJC2f8r3Ez8fNDFJaBVLLoUM9uiyJuv+60Uv5XeBf2I3y4gGGTP40bVzvD3qX+b5iW7T
txhF+4+ZzgP+gMh1Hp/bWKrTshe7RsuhU5FUUzp/N1/SM6K89CXN05bbX3rg1zugl4g6TLV1vNXr
voTHOfObcs7DBS7sBg6S/GDz/vUe56+m8Bgt386Nf4Hx6VfhyN+uvJ+fJHbV2eEdjsEGpkzJPY6g
apIaNjmRx07j6uhJ3JqyLeYgVcjhMe8MtvhluiX8S/LJjQofQ5ne1GvYg1bNLwMRHkwBQcb93/5X
o4XBVq2Os8z/Au6bkMDQF1IHw7/dbk8otoE1YVjm1fqoX/x5OY1EJmr3HuL9EJcrltjG1yeKkFXh
RuB66tyqf0DEWVaHd9CBxSqTnB9vt1Ycs8MAclrq5I0hp9fZ7KDsqR5bxMEJoOyRb3/LLbAqxHxt
Rpd9mH35c3A5XjDGCCBONRQud4HNxrPSn6Nq0cnaAtBCuoZUUMiq67B5C0MGtLP5RM2uVU/1TkVB
G4maaHkOBMiF/Db0zLVu9uASvt88bUuFzXQAXwiYGUXb8dSmpODhCRuRuhBPgh9ML7vwByfshueS
jHT8b/vLREhjdriTP3MhbhptIj+btGD/dXfhWsKEfk52S/vuzvFDjcXc+67bv1hJSZg5r5t+APLp
0QbykyRK5o19bvSUqAoLqQd9t2JWloYL7Mzyl1y6CIhsCTWl714JXWiWfbs1ZCjyhQJ3ElXNLXgL
X2VhVzs32r4ToIqxv0bOj6zrGu84mDHFr9hjwBMN9sbt+q8MrQB6wPG81eqx6d0WUvIKBGxhrey2
iZuNVxjB06rMNijWuyGZjfKxVwXZA/fOjVMlYygOvJK57lGOeu52mk5bYBpZJmOBoGwu4MNaQCL3
FHWrtd+Uxc6aFh6d/5XViTIULatCR1Cq8/rz7pBLB/ygIyrXkB9g9YNwNuSDf3saWyZXe2G8kbqV
fBAcLxhDnyaZNN7kZe2hE/2BWop2NE5kPaSGHX05Cvwopd9BaLV0oIYCxajTwFydt2YyaeTYcaTv
vnSs7f2XNvvSBbWWZGpSEfqVn/fak5MjVeTLF1fJyFV4ug3B/aRitcXpI4ESVTpJmse058HDxRcK
GJ0gPFcDtfud6yLkGZaFpcE0R9TDJAKOfSfmBKecRSeXarBlCshqDKSOVvMlrrGseDQpEolIvwk2
PkrocuvjpBupAW+sPG2BV7gL5015LE+bqE8DuYbofjkFfb876B38n0x3cAYPr4nYtCz+lc1jveZV
gXH4Ko/i+gpZLH5axovfYnoOTYb70PKSs6BsMkPzemqVhxIygFCQWfvCw1Cka9+u3TdG0uTHSOrK
EVfBCPq3+ZtnzEfyTdwmOMIUDse9Ga4qUuJ/wpij9cp9JFW6oszz0CZJMZhyFwtkFtNPVc56Hn+3
ma25DdIEAACTmhW9F3tew8rl7sJVidaz4Qfj8k9HJ8sxHQ0OIfy1fZ/iJqCWpuDZ/wvrLLbaaWI6
Bglcm94yUyiWfJLvfjZf6XeXWFhZbsS4hnt6jKnI415YlnQ81/i6EriwkaKI40jXUshuIFMhrjF3
leFQp095TSCSu0Ag2zIUnKEX86NXEx4vlgmlkpDc1UMYHafKhuLsxa9SmLe4YBEl/14n2YuUQ8Ka
6XTkD0Vb0O1bSYQYc1Sh1P1oKA+oLYPBWRnIjhIikeAN7h9qzxzGMcrnKKs4l3PPvd1CtU1kTZYM
FDBZtsJyA5eo3caycZKtLx00Zn0/QTwmWYwFAHBMhPw+CGwqfz25Qneq2AXLrzUgn7VoO35uiqRn
57wHtJIZn95yoUa0Iz/m/UkoyPg8rMDu6JH4ObaoUn3N3odMWq14M+LYOzq3D2MYf0YcQ+kDlYHd
moB31nVnaQLizBvsSA5ERzXDp7oemEZyMP6wd8FwVlNWgy461loFyWEwjgrpdLOdywde65rTYTqN
JARF5YrjlZ6lorrmUdAA71fjCXXr1679iDHbrACJJjyN/dkbfQ7ZP1hgJ8geryRp+VT6K9HbnJwm
m5wxzU7tr6RJcsOFHL1vxNsSJaJfqYmXrLmArPY4tIbdVQplGe2YJifn4siWZHBU2ehhFV8d7wd+
h+OYtRnzvgcm49qzlqYfvKpPdtAeqUtVhTAJEq1/JS/46KRjA/fTJZ+Lh/ImM6vZ6T6sFJNuNHLn
yZU7Sy6QUCf5ztg/4ydXp6yr7lbAgFOyY11/zo2QW/1P6CT9fi1ItIv5re7dpp7VCx75YEbOhei5
pFEW9l2ICvUgKMGPmw2/KqQRf1VT0xcezeDHfmzOUow5lwh0q6EKxW3iKibuDU9e4KWTzB/G+Qxt
ZVZ2KN+gPYtok7d06j8Jfc7glpxErdu8IHFSNsQ2+v2DW/6duukUcXI3GU3IZYkFfCQZoGydRSTT
WHZyaOxVi9ygUVkZCAXxYzJnCXn5iHdQmB7Ukjc79wQALtbr72kli4LFs4VBMyBW6ccQmnEL+t26
t+o7mP1cMjQwL3NworuMVSkcZv1kgUhSdT2SQEZBMYFwocREyDau70C8506w1dXHAUTfXgxQROeT
5Y6waRR7nxTpmKZ1MeisARPSa+HHd/2/OsxWXwlISaJkEKL5WzO5U/+ul3weyg8lImtt7dRW88jp
kN/vCoGkon827Jg8wern9D5lH7+kw1l0qBZ/yvR6kc7JdoFjM82wD/2E61jJ7Fc+ZqQMw2xfaCJb
XR9M3cjQdrRRB5zIqz+A4jrkMJirj1EasGk2OtM1yG56jMc8cWNLwTLLb78ZfvO4CNmqsmHCU5+j
8gCwSQucyEYkwk/9YCm/he2SYU4l+latZrN69sUmO7JwCZYgF4hn2CRubDC3Kv2swmDUUoki5FjL
0yufACbmFqeyxbWMWqp02z5h2ppUIL+JoMNpPfzVkOe6MNaQdqe2sCBNwYeqS7KvWKBxT1C5lQ49
7gdNdboysXggRMH2z66UbR4lW6JaGkk2z/iw89NpezLzXyJDh0vuCF4q/562wpdAGIhXit3Bj63X
d4if1WK1wTbi+QNPr0dQkLvBwUKP1kxeF9Kkbi+VMdG8FLZfh62K0wHVtVwuSRDHYOeIMSp1X8cW
ApJnTPjbO9arp4brtCy0nAcXT07Tc1trD206g1xSsKxS6P9xuYOUqoqTtSzSQSGMvvKEYRKE0BX2
v8ZMYgoDpN9AdnH2JrtqEZftFAjgc1LgjwHUKcdSBQW9ib8k8V3jZ6ps+EUoWC4mBX+9ftG5zDEC
DEYcOOtp1Y+lAqGlMBo19yeW4xaiFCr4wasEHzwuKHyiiL/QqJbdoSxLcDXcjVH8cLpB+vgiZimK
bsSUfCi7tlKWpzbHnd2OMwtGM7gUAvNI6gBla2d64dYw5ULzT7brQ+m9A6GL+0/sVzKiBwe94zbz
2oz4vI8PRDYj2e+TuG4x36Mlc7HAB0NpMAUDnxLHu2iMLPyblaCj6Xy4h5AHSyCyTZ0ydVNIrN/Q
ebg3FHXWgtewITYgkjfLGQYA2Qb0JnK8Cnhn6geLWftuPcX0hg7uZyDb71fii6EhORuiUqKkrHhA
PYr/uWLw37B0SuLgDyThHMU+KA5cBUI4BoTwg3361Jlhyk0agOQU8lrcNBIPJ9c3l75UVBQrLq6F
kZI+BdowutDbCxyRKFjnopwz9ZGvKGJZ4eq0sgZaI89pt7diJeYUhU3yEvRshRCp3khWY+S38w1h
FbDB+Un5Mkydt+d81hmtFlg4JC7oAozfaBqe/gn3z2fN+wdngaz8oF+/9z2tQEJyw2JwaKiRYNm8
6issSitGtUoCHs6rvt0paVGzU8Jo68FxXIMH9lGss5QXT7M/USInGPs79arXYroYY40Z1HYsE919
v1xHzH5ZuGEZJx2+qDONH2JhIHgei3t+CzsZyD1yIf8jLDG3ASsQyIt5eIYgubGrYpHjdAAQjpWP
4FbuGHdmZCAnSOPciOIqD0x9q/Nm8qgQOw+OQaAcWX5GSChCt9Py6+5oEag6/QfD2eWFL3SqybcR
HJkgRviJfkHbgQEX+oC2DUNfnk22rnWxS4ozKgGqaOHL1gsoD7ggrjWZnoGMXLUiHKI4IKUGvQBx
4yqp7NZAPbIHP1VbXvi6m3wehcFBN8OHkumEc27R26pnbMPovQ3qUc+QQj8qHqn+CFRFX5MbNg1q
NcYo8L9T7pm3tvCxZsn7moHNWHopEZ318VzOcSYr+h9lkv4/X/zWQbIUJHFGQSlk8GUxL7tmwbZV
wwx3xNb2UjCGc23KVqLmqOigvM4+gaRWkiZTW31aLeOuDxClZAT1hskE7om2U8sWBtpOFNFmZSYG
Mn5PjFVWHwuHXnJtq3VH4jg1w2LST663oG/Ez2skoexnYG1tQSDCzJ8lhvQfyW5GBC9Gti6oDnyX
scTpfatsEKtGyqFUQBMxBKyd/3zNTbwe0w983Ltu0lh6Ba86dORA449Iui2qzaFLFBczrZ/ca8T0
+tXZDUoqadYjnTi9FeOKLbpOSh5mIql0OJvAdGhRij7y/5Rb051FAS+uOVZDU4g4zA6NuRGCjRcj
inD62B7I7VAufTQNgQjR6KUdCKCMT55ciiopPP/toji6sWyrOdFR3zZQxO4Q8bu2WAwF1NUnlznS
dngaL6C29DhCBwMe1tr5wfN/Z+VdgOgwMdi/fOb6ZfgXnb1xJwQozcRbxDs+RehKVgbVxX2MPe56
JnoQlh7YsjzxuMABPqLe7IdK4W6LHZgl1S/XpQJ8t3bboI7bMcWQYIn4nA/TOC98elYp2kmW81rl
NlCoEESQuUaS3Tp+5cU4CSlbb6RNVRo31MxeeUfTHIbJv7BMmkYZRT8kLx41hGl+xv27USJMpf1u
XiKgCaZ5AVhSRY6nOgiIzjuzJHdLg3ICeu+1GsRr5+meAjlmFx5lFbW1GactoI9p73aM5u8K5rpa
EYjsG6l/FsdDoT198J6I0IVGiIXNDQpxH21fvUvwCEXAQKoZgrinXxXrsMkVYUcUVrq6oUeqwF2D
byw3uPsQeIsny40xjRaNIoMEL0BmDZr82Y7gP/c8pLzCDLlA43YXfe8f8IfdU/Z7OD+8H1VRR7oV
22mLGsQrVnIuLLWbLNg/WtX9mkaez+buM3CShDeso44l6P3YfA1ZncMyks5eXM/HTSbBoKnTenWm
jTxYbIA1nXfqMgk5PscMslqrIWZD1V6Jb1Zk4HA6Oy80c7MgcfT4IxT7ItD+zyKL+W3S7IWiRPed
+0/9fwOzdHbn/AaQC0VjnLA1WI+55RR9CmJrWf2e/8UzV49sHIfno8J9v8wDeRYT/V6M5bClu1Ia
j4p1Xa64HMwxNwPBLElJkWtHG8pmbvKMbc9x9Gg6B3ZrAtI17Am6sHMZiV9+muoNUF73zNgIXQTr
L20ARV9r7etXg1UPbk8x7hEax/LerHHcu5eCbo4uNX0jmLw85AiaWXHttk5PzRv6i6U+AQ9S5cbG
Te6amo5480LT9Qr2qIz+d+LrhiyqkDW5psIGS4d/sZAqohSUT4F7A8hI7lEjAaEv3WJmIYnzn7DQ
skwp/rvxWy5HsuuxZeh2yU6Me4bt6jgfyOZQk9S2nvCuD8J+mAuySttaE3Vb9K90BkniHPDQyTqA
BG/qinKpgehVq6JSNgoQ9LzVyN6fm4lXRTM7DvvxABcArjN5WIJ5UDRddVKH7VwmXFObQte/r9fs
Xeji+1sxYNkMZBd4WGC0Q0aUZiZKdNnz5bPIgUFLclludB7odAVLD7sdvIgk2NFgtORf2gjDn1a8
M2V0gJgqfhl9meiVPnEpxk//t9f4CL1MFVDBgYGVosoLNeswzjhcprfWynprRcYoPJ6DWTp9QKdA
mKzD+bwuQaDtvKO79e/+7vX76kT+SEt5PfEy4VWiFLUIN5beVwRIWO4PWy8KHBfNGUOpDD+hQ5Jy
gj0YBX0jCfShmqB13t5Z4aIlQ+ThcLH4hHM8fBwtkq5ssy+XNbzQRs5EoNb18xVTjsrb0xlcUAHI
lHI0gwxe909C5/X6VTmKg5z7KrMUJy7c6n300G1bcxM5Rh1imnFNibMIBTrvYANMXJAntTsXDIAs
R1ON8FOm+LxREw7ceNLBlZ1sYzNMeBHRITWUUe+i887zJSOVwQKl+anrYMLe8pS6jvBS9A9B+hXE
pPBEbxi1HHW2hi1+/1yorafvACaimfCDfZYptojajcTY9mNni5ZSq7MZmwuNRRPUtrTTYwA07UmU
bEPQJf2WqBFRbhCMz82ozl5PyvV6eK0QL+6kHwtNVs0VOYwlKVjRBU/FgRNIlRXuW77qqmtk3GR8
LNc4fSBmybajTHzFGxKDR3TKNHnm+ooqGhCyx+zFcrr6Uy+EjeZncS3Xm7haQRiDbS+iDGyYHL0f
FvPnnajn7x6s297p4hysBhIZyP0ee0YAR1E31wk5qFbeMPCsSWUoaf2zwTGx9psGjzuXA+YW/C2z
K/sJMZZKjZG2Fv/xD3rVsr54uogE9yog74tHqT2Kab+Hjq+OHsvMRZiJhfiMu+YsDN387OFiQdDA
Qczb4jgTnvdCYUEf/o4Xr9OWaGZ9qMLIV/z81yO1waAl8czBHTs59N8T6/94ANr/+SHu+o7fASWC
6ji1r3p1Aw1kzjegDAE3ZcZ7XCXMEPtpvc8keUHRFzJvZ/slHv1A0MAvNCvT6nO1M7afS6PLczyG
XOultKpI3HHGhWCignOY4779HDRabacJSYpX+4TeuAyOBioGd5yLRim1pqJRP8kX5eHFV5wDm/18
j8Br0aSrQXpFH5nAtEd0LrfPJSXOlxeiYtCAnKtjA6NCtcIxtCjsgNvkKsoGJi80nen52k5xrQbv
PlXXf4h2nf2/tJVgOHOx/X5qS7snJ8HwCgsFPSnjMVaSubijEq4NCfL/m2ilmhFNSOyf0pOfzIk4
zI1raD8Dgf/XZO9MyIrQ2q5qiqZefoZSp78j2583T8UyaVt7i7zFy5QnHJZ+mlFep4HgBr1yO8Dy
pRbMdCEGGetOmeOdQoDP1nJXIiKPrz0dYQXuzu7osdnpvUHCVgUsfAFeHQbjUSe7WKBpNHd2z+71
uRoIxz5CmebdM4MXgHgP3+SKpqxQztNBvdEeSmVOxy0kDkFaUT5q1MyxdW9QHaNYGVqVz6anwS2W
ZVkWQXOA7x/T2YS6dAba8Ha24csZfsIaYybLj1V1Iwr7GrlBwYEGC5yuhIf6v15jWUKFvG1b0TES
TeF5620x+t65NquQFWYDfPSkvBY27BqNKRaybt36D4C6CxXB9xKo+TlmKZrA8WaamnZ7OmU9/OCu
102F4v8oRSGPE4gNX17KqGuEHAjmwoGPXIIpDO+axE2Mw3BrgBEz5GmIxjxAFYr190NUFY3vv5/4
rMn/f49191p6rTcKezzppo8sertcW/maQKnaGkh3pvOfCL4+uQ2ATkt3yORZ5ed4TOjaW3dIdiYO
AFCl/kiYPm0KrPoDl8OyS4nggMUrNV6o65HxeBHUBs4uSfgQYvkY4sLwxUwwTT3wsCMMXORgP8Bn
NQBzZZASd3RpsighxgNS7KVHm7gFD7PTlyCl3uOgFBDxcX8WiLNHl9CABv//6fhU0xzUYzi/vLPC
J32CVUi0fpihVoLqVn7EGVjRA56ajeH75+HAunCzSlSSiMvsJRnh3W7yCh9GXAghUuYS8M2/oVAz
NGuaZI9RxoaHYNAbUHXEr6XLal1/W7e5zT/Y405evEdwiujjHe74RuMP5DkQgm6fB9p2PlIB/kFP
NMAFu0gry5HsReXHLa2gFm7iltZ7CVP1mePFJtAyrmz1LfSZpJoByVB5Z7jDb0xSzOW/U/TzEzjb
Vg16X9cN36qq+qR45yYECyEtfHr3rb5cLbi51QbJCRAeUxt0FVZmtm7241LoZ8uLUaePZ5YaaCrV
NCFk4IzI23cpM1iJvPh2r/bfG3RU2zFpfl2RhzJdPVufhb/OPl88l/eaPQRW+mtvI36X3Z1WJVMF
vpnu7ws459kyACgzOB6IxyaOssHyNUHL8LXc6Zr9lkn6Q9FSI1PvW8RfBPbTh83Jd09X1ly4ETMP
EreJ9C3n3g1sv2aJFMBszeKWIZLFmFTGIQudGepEYSdrXDsBzGFcUHyxcRdYYWzFJAJ5JLhA/Rxw
ecFkNjvCdp0yOqa0DELLnBQ/4Rt9pvpBaOCrM/+nMZQ9QGGXtGa/uSzUOEKT4fMbIih8Klw0EI/2
sp5aM+n8bRMrWyc4WxRKUWJk7uY4Qxa+QsVjS0Wa9RF9FtRF158buI9kEgjfVtJ0hq2CT558ZIA0
OGlalubvOyyuuyUvGaY1GOdNrs/AqPITAC+2EaZZHaGowflND+DWZ6/DThn9SlxrNa8klaOTNVyT
6qXKUtefo86ahHGd1b0B0WB2QA+zU9z28n3xj7aBsYF3LURJGGHenE2Z3xv+iP9oJQr6moAZHJc3
k4FpJmMs4taxRtmYma4SBDIrZq7O8h4Ql2TG6yVih6sRvvF6+UYerG/L5UxIIMlkOAZezxINJpLo
lG4KaBbcxAkqP6Mom4G3gKkBjTiOnkfn4dcGv8mwOx6HxQjPInZ+X9miQ3AHtL2NigOIBHq8rLL9
fZ0dv8BGqLEQydRf50gPJ6c4AMjPH/sSE8a/x2g3fJP95HCMfIadHVJ6BSWest6SDw1fwipt9XdY
ekiSCFgiJoDAuv5e5lDSx86NIR0uXIhpWZt+VQoTqBk+XqONjc7olX1Xxfrcd/LnSlCn3TydLqWe
UGnJEdA2e1rgSL62NQNW7jKbD9hxG6HU/xtcQOYL3u8U5CIaaK5W5OuwuQp4j4XWJaCzdDOPnOJf
QxiQbAydlJX7GY50x3QQMoWkpXrF9bJYEKM6GP2f9lmWld/lDlv4VLaO62bBD2h/T+2yfSZWOtu+
XgQo6et6z5pkIsHi2hatlZ+YAIzDQ1d7X8+0ev63f+07lglYeiVGkV33Ki+oWEHECwICSpCbap01
E/kmk7nLbiqFjOn6vzB/mYriIpieYJgzUhkdw41byFN3OnK1JFZxNlO5UT5mKot1GoCNFncSskEX
+NLVP5qtqtP98YZRfvVs/drkNcsyxEFMWHHMBhieiaQUOMPWMZhKNiLZxeLxdhG7tVyJ/PNIAmNq
xbeNy/ZEbX6TTK7WN+4rfNs3ux+ogggTks66HzFzDJ8FuYeayhV7VR/DX95DsPeUv+WzbqqmtQn2
8X+MIQsvqL1qDYM04U06mt9u9WRY7059reGBJXy/84NH03UimUTi90rxKiGJAkrvaH6q+h/k+Mv8
cUgdFqmFH/aMcGSTEKhtVmlTzQQhwoXzEOzeKcK+cWYHpqh9r2Cf07iVh0sF5a1vkj/rKKWaPhxz
rd3uGKM3UwgjT81Usy7IWX9g7uzKP133ZuBtN+K0gosMPIgLpVGTHpZkeqtp/L9kn6amSAEkFKN3
yh3YYY2/F83i7vdMAdV7sFvmYfLyD8e+1FfY+c55Sv1YaX5EzFvwcepsl7W+QqcIp6JevJYTc7Ma
6AHCAP2fwngsYA+7itc6AgCLfOy5ftSyoewrhsFxfgYxJlNokZGVIJcQkzLiEJLjgrLh6s7y+pV1
Y10H32NvS1+OmcKxaitl4Q3coTC1SaOmkjhOWO27EtSrjN2kkNBz+g1tf8D7AJNKlrFOQjGO6dG1
AXqXdlYs2z4tZfZ+docMHCZM6DIiKAlR+v3ZUKAMrhZHLIXuEKJFCmM4iLWq0QUeoelzf28tkM4n
3cFfxJX0qwlM1+bGcnmTCkb2hh8YqZBChEwQ0IIiTF8Hra1G39zimDbtB/gXoA6SNX/fPuZ9AqfM
SpSUq4Ta4TKlCC0bWY3vK13ahdwMc+xBglohV/qRcnIStmJnTJdVYhkSfNlq4Xsyh3b+YvYUo7tk
NL7JJL6xa0R0ch8cuEVUo+yWn9KCBsMNTQY4JbDggr7Tg9FyeTdy/MheMa8ODPBixUq15IfvdEvC
nkcqbG5v+08r52uf1GLNSMqRl+0VAch3cNfSsgDYSE2PaQB2wTaoundd1e0T8Xkgb0uNrcCEogSn
DVsXzp/+bvDhbE/a6MwKZrsi2RXD3S8RxmyJVGNrMi4nplLBaoYg/BCUW3Zw7eJ2DfQZFZYKA8HF
09qYtxEwwQVu0I65kmCGRC6wpen3hqVYN4V2pv8+zW2dMysRSqzCIDzFvA29HKLKAVTtralfFFho
KUWGapwzs8AikddCf/rDrqpgKV83EoWvL75bWzaFYcbq+x5Vh8EVTqKfbNyLCmcg71KvA5V/VQk4
aBZBI8CL/xuTAnzZZa1TrJFknhV2jGzyErojSxmxl6AelX0+KU0tMRmX2Q8uoxDwUtRqyw1mGrzz
K9VZMM5v91mqdRgKt2o1hk9XApJjUoem/v9TzYqCBA1hR2paa3aulzWQ6gexCMhaseGnifx5hTi8
0/gLrWmean85cOTrKPsW3oHsFLtUf8l5ul547xkuD8/VR4weC2n2uCmqPyfS73FXU1GySp87TaM/
dVoYLWKQPIu7WQsRFFHRZCQkNxLZ4daY9U1rFm42GJTehouIP/XcTE9NDI3gwT9+DzZ71Ynkcfb2
fafd4IkfgrdMlBzWN/8Nv6ENrkjV2r/tmoXMjq+h7w49kOneaG5gQmZWKPaz9YEhXS+fTaOCLAU0
k42mwnPPSPr1fkQbFTLqkOaeNbUsJKOtAYFMUPnXigsFhzkX+xCDpm4NHtDne9tjtVS2TLEbvwAN
3uCEiccF80KsXZb52dPho72mtarDw6ZmycWnZdqd8OWsuuiScBXrZx1EnA48uO776TH1O4mTY+JF
wRTqrClSxrBrMxFt+Mpvj0Mr7CYHRySg5HYMQFm70rSwNG+FJt2E0xz9iHeZJUUsUGRQKPIJRt9Z
OPyapTSOMsbSPq/LzXOaaNkkNCfcARBV2TyKyYI07C3ux+WOm7xDSedSMs3XSwTiBuB6oD/62VBL
9HnP35r15WNoWme2JoCgdnhmTh49aZ6OdfzoogKJK2YLd0Wn4f3penGFsk8GCOWtGXMzLXQ5owsa
EWsipQyA6Br5ILPLxGEo10MLPeLUe4gUJ4mArE9v6jHq/hvPfRbwazaNJQqxCLVR5sS0xAXPHj2S
DdreP/UN6Gef3boa+hI+pdmAJJLMcf6YunXPh+7bY/wMvmwR4pxTG8GJZeIJi3f0IQaHuK2wg9ld
s/Y45embpAANWnyLOrPbKiJwO+SOslCDlwaCjQ6RO49LzdeU0QBarYfBgSnhYjYjjs4Age7qsCak
of/cdMaOl3vF9lagrddIn+0rmlcBCjz2INphlQ1t/0AJZueGZ89E+kHx/sqA6PYVL4x44kkttabB
VFmLsCU3eYnPSwkAZWB/XnBRiG5WlJWAgwogYVHETcK1Ud6ze5XtlGoISKhzeLUoaxyjcfmXI3jk
yoOXa5gMKGnDBccpU32vYjze92LJMIUhFlL0HAXqA1vxwztw9Qwh6zolTp/TVmbdXsLONXQYvpZR
+ayP2TgAuC3iAF+VoFBsSc2sMkfpDAwuKaMenB1/AhAcUXb29BFMwNHMrHqUfdGh+4Ha1s8LinVB
834mS9Gae68w7dkIx14Q69XvjCVTzwExx1cjuZux6SNXzHu96HD+eV9tVIjF9sZzsgY+09+FZgAh
HkuwHpWf/aNL3R2idhpVPbRySLml5PaFjGqN1oZSk9w2BVwL9cZuGTWoqAG19b36G7OZ2dG2u/0G
D0CCtprb9ERfW1KNDko1TBuhk4gm64Qo8/uggbTObTdIqCPd4VuJIXwllErfmjmqRVMcQLwnXlH9
+wNQjWTkxRQtwZIxPVGxhAvE/ilzlLMd4xVBgFPqNwZuRAicKaqOplpTKh13jC/+ktL5Nh0FedIr
2tLNmu/loF2XKMTRo7/NxoZqndXwZBm8YBneTk/rtxbdz3LjxmQNU5jN8GNsqDpVjCe2bGN782PM
IaJ4KimNjeDsQuVXCpkTcDrYYx8GKYD5/jVSSLt264diDTlPitouh+/yNhsZXc2I1NMwzpQg0mn9
rJmARUiCjLlUjLd0SlcxUP6sboYqX53yAzu6YsZTYnoWsQVJmJI0RFzG0Kqxg0UmThxYLoVZpt5u
AiHw6A5pmSohoBjmXmWB1cIbU1LHqCBGVYBDbygYS7nafoVFZZbW486ZH6qsNeFkGdh0suyg3B62
v3614NnUWVbNVABSk4F4lDmvaZvk8ZMg7XCgRsErjOZCPPcd4cWNNulmQC9CoiaVt4cfOpk0UyrP
0sOUw7ZBF30B4Vyer+5Q8mcEcHn+aX99ic6vWGI2lO0WYp2fv/aSR14cZCq0Odaki5BO/33vtaKu
7Pkmzek41IYPp08ifDlGXXqBPi/9d4nZdXSc9WL7yoBEN2BNCd/XEVMGCsHSXlLQNrr017lCGgOA
jOJbQlkzuiH7D3Zt9prQqbDa2l9XQ8VHv1o+qTLGExCLLnmpQ0gTfOVAZ4KmjELIP0WbivdxrLrO
X8dB7aa62ES8FFA2vY2gQh2O5x2nA3BFxLccYNE6e5jaGQVjxJFZpgI1QrsJTjyFd5mcwxE3//5k
Ws4BlcPmKfyK5DZsVK9I7RkeB5QmHGCVzNnGwbW5IxiyjWAVAG2nXocxVcKHzVrWTSy34RmR0Ut1
alMRU2wBoSgntZjwELtVa5a0yEu+8c/mE8T3jomCYQZbRQDJcmXTu8aJb1aipFJT/L1yikV8optF
1BJgs32qpFaDACkyZXsIPnVyhnMXXPsdI1PZtbbXJkkrMjbte+UbkRyrKR74BQu3pgtXZvgmJ1r7
l4+XYpWptMD3x5mTNiG8d88g2Bu669vSXL2dMdKsVUg1scp3Kt0rjHj2Fmf26SabWcPlmdt2sMl5
2MsS1eC8QY1kvmLqHW93Q8k+7B7X7avyAsiH0WzgB0Iw7Lb9D4xiavA1DUVsmJxfc60HFfr5Fv3E
ZG6TVNb0+RLlLGgivrd1JIQnAzwnQ2RDYYzV3FFhlpffcZuvpdPM9UUiHAmJu1clqMiFojxmjhKa
e6XICO4THfT7mruwaUV428Au6BDF6CO6D3bx3+txX17P4X55fQxU25EFBGcAxlzvEHvixKXEmG3S
0wRRoDBpQR2Cgl9oHKtB9AESSXKJkF+2xsmevLJBOAPyQOmeGg2HFkTrQQCtS4fKGEdgmXrA7/MK
c8Wtd666pSPRWdPnzVWAZ9zP23lcZc08fjBBqQI45SsjcG+gfGj0Uf5w5vL9qZ8NnJd7HcN8FcNV
f7k1uVxEHQoDfiC9XA/T3l//QrE8U08DNtWEce8p4AP0LWodA4vrew/JKmXAXJs1WmlLg3CXGXLD
gPTKXqLa3nD+lJuAp7C4fNa2fnfAgLBpXsZfZoaevucp5d9iVrHptfpvDSfzb05K2h9VUIawJmUY
AUPikOUbJI1Gj5G4Nw7vN9Xge0D8O+8DCc+XcBEwQWkc3FGzh8sNu1nUUcru0XxounzPEtZ6mngY
eUDSJfu55i/qfMO1ywBhnJGUK7zHqXSTN727r/RCPppEpwclc50Oo5/pWxHHCE3OTZ42y5xcI2SO
qa2K5YfdSqCDlx+6iDQ4rN1Auqb2MYxLmRebeUVIqx+mEtYLVcgQv8fn87MgUmmEvIdvNJQ1L+Gi
kSMgca8hFq6E3vWkwiHf8jHnli8dbJvag8yn6W8HwlXyt2m/kWOKp+i0WMcqYpHiSynhQkR3htyK
pldge0q81OM5j3RpLTyXm3OdahTbzePJ0BUMIlXAT0VOkKZ96GcCYYMPE9UDrw+qRLRyB8Kr85a2
kZXHT64pw3Y7hyEw1ql4gUD3pPJ3SbhYdDOWrnCtmt3Zq2KNjWF4oDKW9eg9Zf35OhLlNVNN+UTq
TlnOWWQr2aGpW4CRY0RyrLJvt1/dkGi7MjWd9XVuPvHUwcCY/8OUteYLfkKIcQcM0dCX/miJe6+T
IH6uM35pSN4uPN3Y5izGtyDCy8M1oGa44uuDWVmVBhXIh3hTrocyJgdCiCIzhxukCJR6uxUivHQF
B8LIxWIEYrtUY2p3sOuROu2wNSsfczcizNSAAocLBpPfckSi1DCecAP5EGCc0PIhhtOnU/zImpn9
oKgQ1nZ5W79JPO9lgz6ckWjoCQT5CNkTsuEuFcwi2JPXo7lpJlu8HBaxc9M+mNZvYCdjFmNAgTQj
elYXr22i9uBQJGPqdNHdal2JYlqfAJZh2j/XhGVhkTY8GHKsHZhAKoKWrP9O2xWO0TbT8xn+231l
vTrhAoe/DDETa1PKBejFrcW7ht4PiGHp0zjbYSppRLmXeWZXrFyKlgbI29SkUugeakjXvNhnTKNX
YdtrLSI0Fye+JCYyW3k1yGBbCGEELJ/nKo4xtMsbZnDtHpa0DPZM75OSRoHzzBy1Cjte4JUFNBKz
M4RRRgiPUR0mobE7uiN0XVFWUgguPhIKGrNe9Loqd76tx91g1RA4jOwtd7AtxLAk2Ozgxho0mKRc
5RIAB1wmm5ivxYqJPS4fz0Phz5Ur4AdjWeIpmUcfbxmsYDu7ezhqXPLJqga/cVsD+PBIyFg92/5c
8E+cM4d7so36iZPChbVWi6adbP6YYlKv/m4y04tqyBXd9teaH8fd4kgzsg7GlP+S94yH/bileG0l
SiEkjaT8TLAsMp+Pi92PPYBUTprFVgj3IT1kh1NEYs8JGvMJ+yxxyqPQJkBkgabMPCNL7B0c+zCt
LeY79x2OKbTvJi+Rs1+qdUeOiKRR8uoEbWfrV0E1j5MbbMQJzcu1QCfJTGlVypaeXDQ3HQhamRTi
efLhUveGyIle1ntSCef42oIQYItBTBB8yObpVl/VYqaPI9PNmZijJZQ91lDRoGdWseiDusueDU6Q
flOxrvMT4/z34bTL/Sm2/1jn4LLp+MeM9DxttqQHGg8EdVIA0lUAnqb2H/uDP6lgC3YB9EXqEeDL
ektCnGnBHUv76MUX05KbziQwIjwj96BQ/IXnhK4hK6byuebnuhRmOcibB0Xw6CVperr2zBKgj24Q
HhEZYmHf58nG7VKnNbi6lrtCmK36q7M6AQH7MaPQNlxycFmVFVMZuaJ1yzkun6NyJIzq4vVnIhws
TNjJBQTJVOkvwwwyspkPJStL/rpO4ZZnEQ0QMUHwXsy0+PaNAHhTN5ysLzd6vTObaYrEZR+Z3tsX
9gQJY/2utw+yOV6NshxxEmCd1Le/ArAlmzyzMPFKuC2Unlo+A9rqiln8PeiVDnMT0M3gVuYMCjO6
M02bCPXJYI6E+WjQ5cYg7n1FQ5ZoDsst0QV0UOC/TcB3WKGdZJkkdIQbVOSM8T0DfO1djDG+BGLd
X1HdSqZCmAxaInTC4OEHMz9wA+mKlJDVH0cjOGpn68yhO7lBBpSSLkU2ejFNujw0sUOG8F5DIAqj
czV1wRE4UnMtVNbBneVDQspma4NUCPfE55RTJxDvh0TK0jiRh8Z1AyF+7Y2f0oc/hLL5870rU5Dd
z06YS9P+QkfaDZ8PcT0pNyBmcIcnLF8Cwkebu8O1RScC1srIs01V/GR05OvIW2jlSh6BmnUKqOXs
Bn4/YZDrLTZfKEMbv8CLDbIgYtwA2Gx5kE8Bu5k4VdlQjueT7e3hVohaDfBfk2vqS81/zD6kb9wO
WzYR6jV9gco1g03QUOyInnQK3TjFT9VVXG49YXfz6il0XzrwmHRa9BFQVkN7k77QwYrg/aYf/XWW
yUWIGy1ZxdagOjajSj93vEXAJCyhripNFKyWgyfeaQesKWLtkCEKkFEuLLpXuphB1DOVoYBNwTko
2XSSGjj8D24mTFpCnPwnOrRqbW2G0qcT04KsvTCUcZAAh5ZjIL4K/2j3jCb6wZpbcjb6FoPs7NRq
WJ0mQByyHtit7qeB0NXp36ZuUWoIBjHz/6XNJEff0BcwemLZQjBLx7g4caZSuT0nOICReD19xjPh
YP0DJUCUMph83AKj3B71PyW8GgKYypOSAhFKRKqetZULtMbZVcpQ1JR1IjWmhOF0TnHKQHp53bgm
aZ1JAVwfOjiPIcXMj6rNC8Py/FYHteWA6CpSJT+xXLRyH167GHC0uwE/ZCWiXEmr6/jWmRHeqpVO
xh65wD5xTQ2EcbBSaZeuC5FWGPBfbbwafqss6iD7P2AVYdrB00BTLdPvOuCLkArL2E2wT/jDgC+I
O0zIkwSnjGPbPWp5oACxiWYR676y+xl2Sm+AAU5mmc3hU4MxG8DhJxIypJurpjd7f9WOQ0MK8C+i
h9QGiiWkCdqGR/78ACSH9VXKwPuZgjOn+Vqrrek31STTCYL15kXvbKfqrcVK/J1W270wiaaed6/5
THrkGAOIFnE2rj9LW+R53IiKO8YCTxR31t2GuTAtuwTtBZVUE0CmZMThS46bABaZPCQBIxXXM4kw
F5couK3b+BHjmEkanVqRnTjhoZg2kM77MFpvXnyJnHnKLB8cKjDmWMgwNfRN+7bG9VQVH/6DcP+p
qOox/mceO1YUN7ujfJBvn9sNiXJ786iJal2vlJ29CPOw6FnSApTMPYqgYZT6EaqdVZXJkixGV8i3
BR4V49xBYuZKIZaginI5DiKT5lHkcVeXhDxlW6H6F6fB1DmM+EyAg+nDMlRsHqhZ8Q02VBHV72He
0qpHKXnIiyV17QdEuKHvU/kB3sexJ2IU/p9uMg+QtxPxON6D7RpugDwTo2amhIZV5lmCmrd8J+4p
QlV3kz8AL25d454XwDwY++rrmbkvMiRUbq2BGrBRWQM5UqggtzavO9xSKU3RRQtguDHre8CftJqf
fcXnHIsOP0EhcN4w4TIB61YoS5gOxUPnv/2nyNZfHaX02JnfBOLXyqeH9Mn0QWCufOYd/wysDkEm
y+HG5GYWnDz1obFz8PH7ietT67lpUYsTCvUGmL4gDowbvrr/oegmHgKvAivSdJiMR9UgtQmpo5Za
XeN4Tj6IBmYtVhr5C8+Q9Yv4iKBufnGklaYem2xLeLZGZ6f78ZcaZ/QXCWixs0Yk17DAbLFt6UaC
AyOH9xZDWMNAjEnFM7sc4lQ4IB4+iGEe51rwJXfOLuydhM8hwas1rqaRY3uG7jGe+ZhSjxh7YB84
16nA7T2IuVIlq6zEx8Q03C0o9rkmonOqwakv0veay3ME5m1szC3kDNu0iYG/KqELGsAnPyNX5VJV
MHYvRf7IfVRY0yEJ05FzYqiXh+sf7r/JtRePYHU41EV9MLGPXTtdc8aYRWT11Siro2QsqsJKM0Is
frr5dCJvLmDteckks1qvANYmtzyfk2uxMSBDrOQ35RLYb3cbp+vezQLu2knUtftAngwoESPoJJDl
/kAHlloguzAaYx+lkkI4C1XNAUnbkXdVeVMjEH/t6MlW37UCpZObdM63TdQLmvpAqXzKvxjzCHtK
02OFBBPULc3i7gac3igzXt2KnIkHMKle61QbbiZQ8XedZLuXSSJuGZJDgw7FzzIaZVXvZ+cgX0sQ
J4KEGJ5ZVG2Yra7PAtF8fP/h21opktQR6CIbiVRMfje8B/rkeYsrEIVwyyAeaosk7JekjjXtoQr8
nm/fq+2CP4Crdt3o6tAqHO9W3+jDKu+e4YjnEiHQpIUE1L97YRUTlRYanUI7LjBQaCoMU+eienlc
FPQ87vOB7eQ273DHKI0IxRJmRN0HRisvj4ePu6Uk40Sx9Ij28rHEUiNG2i1dmFh6Ybg2iLFFhrCV
JaUCWYw3fqu7VQwAU5XgefUP5c+IlH963uEEDas6DuV/B2d2snBO6VGnR14O7eikErrBle6Wyzoh
1/pqvX//jfZKQ2iwrNXP/qlAKChtaU5JthgzTh0QERzFwO5GmX+lezNYi0jOqdZVA8e1CGJizdJ+
zo/lOk+jqEjXZdZgsRmyOBZfF11nkjlQpHI1apXO3tBMjuRJ0hf/InBCYej7KKOt+6SlLUigvWDJ
clLUC/CMbU4OzxLAGrc7P1QMH1ucXKvqTIHB9PiFIYO88eHfssid2Fsfigs84GfYC+yr94dDIavL
jYWz/RhMyv6VldvCm7ftdc/u3v2/A2Z2PyBrNDM/pUXE09EtPreu7ACaS+A8ywAIK43AFDs1V0Lk
vgmx0/FvYlYFHsBxbDR240btOX59H/Qe/wE/gR3kbizfh9QeF3QROhr41/tW8f0ljiDbCp0sL2yK
/JhcI9ZFFCAsAJj/5j0/O6C2gaVMaXfXNMWoLk7dmxR8XhoIaOoqIwebNjH40wavLSReLFYfI2Cp
2TnuMCXqnoqOYYsonxyCYVhQx1gG2YA4cBYAtZHsj0TvC8S1VpV5CJS8aaRv2JrSh+e8UKA8e+f+
OPcDhGKXSaBAyDrgozlycQfKCdQt+8ajlG4xUrN2hgUylmoOt93u/6qNIC3gLKcqJhwFEBQ+RRzr
N5nrqiDG5c4hzlXkfTp68aVSSaON5MbQxkF0ABu74+7cAewSwls3+Mb+zH/9HMh70rDrDAH1dpVR
Mt5sKGbZa7iv59BpYBMCTWQl5PxvlrTCuMQ6kxko3V8AOaD3BIW9V726cAQ1IwKH1ObkD8A0QBb3
Eg27N29ZakvKTf7n9XCqRpAGrz3D5+yKh1/eO5yD2jPMUrpKieXkOSyr6ZvNWZWAZEKD1RxNO3no
tCIVdFXYDoy3bLf+YCbHku9S3+NYHZl0VOXPufdprUUflKnEso0JMemJKYrGVgrNLxUDI9mpuJk6
Y6evkdcjrjaNM4sIItyChcdF3bvjqYRFPKK2uNkv505de6rWv+4ha2K1J2tarI0E/TDc6dvfQkNr
skbEzXWPAD+3B4lXiTe1ebi3YL89fHbjAlEQXoSg/Z9xKL8K5pLNcAk+BXIdK1dZnezQvSUd2h9O
7lpJSJyKhSgj3C49ckBKOQ32XvJ/X4ibSIuzTye+WQGoUFuMqNSHFd+80P/PFMEQO6b3+XNrAfrj
TqG7wjB3Goy/VW2lVoz0xgC5y532/GErKXQN1thTbDd2IFI1nfkUz4QP0JEtOaxlPQYDlgqD8OVy
xyDhdKiGN1hycmfJbEZE1ErE2JdZGWOZwtDi/rQLVxznbdvF6EuAkRoIDLHCicPWOuK69Pl6WO2R
bJ+4gRWhmFtrJq1UiU/yeHDsQXHhzNmaK/hNGlD3WMtdYSzzmqDbTd2wR5sEt/3ZtXmBnUnYRAKk
4VxKmOWvNdDZ9fMmtQ7dg9O3mmlcdi8NehJ+HegLLYs/XP5OmtKlFj/np85UPMnEEA55wr62QgRZ
KwO6OFbGXsddThhaZ6dOvsNO6GRKJQUcFJrEjpo4J2hrP9AxJOdvuFsbUILZ5aUCLYRWWBjWgzlt
pgQAWUhZ8fN1wqKd+a0v8iDdcyUxAntpni5AbzMU5AmC+rRWJVFhtnyPooYFyALcMFfIEgVqsIIj
ISoV+OPD1Z5YlRG9PE+Ps54uIwyrG7tTLhz1LosV70fbH2BhZLmK36/c/wkd7O6QAPQtAB9arLnU
1HLxno0Q+q25YM1w7Vb/mbhaKrom5Inj9hmpJD9sbJYRqlmA+z0cY+WqPsaRxtp4WbU34sTlfjw1
EVk8odERGH0s9iFuK54JlxePemXxy6JsYDE6umPrThhk59JL0VOpL0OeL3l751vaGOF7R94MzD1B
92++jC00HxS+llolmead3lnUMVNdb96n+ArlK/T73o4KCMj8IKWd362BrsWKSIrTbZynJoPPaGWE
c0wNMZUpFUW2BXwozMmCKPThtpLxx3E8Sl8f7FVKtoEkhVbJPtK/LxkqETvhrEsy8tJb5VG1YlGo
cgytGJ/AyOvm+ZQmku5rDqEbySLNUpe/GFj0RIyT2mvWaWGklwTOmdI5sBxhY08POBgyQzp9g5CG
e7PQpGPWGeYRZYYL12Bs1jgyOtFLWpn6BrnkW0EhszI5GrwKv/f8nd/f2dnaLlyYO5pQoIRqkZ20
mpBXCHB4pyZ4feDk4urPDzblyys0d9k+PfHISvacUd3WUM8zzVfTNs5Im7Hm0x1NtiHFDe6rF0bL
V6GCu1DVqu/7974iWcytctQq8fmV6Y3Gt8Gyc/a+Al1FXAgwPHSb1dkpJSPKkYNV9jxwzMPuysES
InOPiNnbYHJIYiEe5jP4ZFCTagwTU6c4d8CJ/BjZ0lr8Lq4+HUwGb06ZVy1/kF+a6M1MdnhLnXDE
w435i/PuhMVLanb9Q5zT3tcj2omdaKdAY2ekpOFMWWRmlQrCgfwyycRVq7398yrgCtzYeqFyqLe7
bylH9zyV6lEpDPte3SoTtoOiTzJSgFldJW9QsqyHtZ2/ICBFaSWRIO5aKZ5iVPb+2+plPW3lc/xM
VY2Jj6NCfL/Hr6B7uw/wkm9iQMppK30SGCL4LPdY4WRAT1yQh9bnJw5vbAw/45vjx4sb7+eLGm/2
ZAOhifNMf2CDW3o9U2/eurLJWMS1aAORb+DIEBKKLN0DQL0L0yfgNsA18jY4sQrSDFvcVGvqU/Ju
w23r3uWMtkp1MPpHfggA5wDiA/Px81rkx08gAfQwljHJW9nz7B8yJLKMQP4LNSCcZC9PExrNbnEb
Gz2cY9hkQHfc5uDotGs4CmAl0tudV4GuFZjCSCTFysLrj2RmgAWka0E0cYdLAve18if+7B2jVFZP
2lY5NpYenX4Tbp0ByhcX1az1XIwOZXLV/RY/B0SUpsgl+Sd5bJKJEa+uGiu5plA886WTdTM5hinL
9HHH68noMpIhgeORyLtbkUF2ubkx5r7HDc6VKbSzXGZ50707P7JLEkx80q5Ldxc3v4HX0djw6r7H
91oNZRcpoELqc6h5CWrHFy1HzGlUIrvJZYAYNvIN8qrItgXvlUUWh0HV7eibQTbNcH9hmmRKuMpN
7dK9s6z5GohOWbtonAKU7OliDOpi24galKuy4q8KoUwlRGOWSmlB2T6LaAkl2hUH/TujsbFeYIHp
BzJF5aDjYen5LnHjxqNouOjp1SjQY5CMzMhlshqjEcrVPhfHmQJOgR/WdiEfQvbTUByp9cyxnNUI
g28iusx+rxP5AATcS2j26L47ZDC8WxfnAXU18ryTtvCvzuvJmiafL/8wstQR+h36r4yEMLK94TCK
guqqHPLLeJJYHcFFR1V35eBpoFcnjB0qIaAYUSKmbBvMZC6ngpKNLZBYnLa944kiAJ64H6+NiqEP
3OUvYlqgI64YuXHYIMPJHcnUK67+Rmr+3iLy/u/7P6ttaYx5FUOcOEE5j0y5lZt6HgL3UU9ZAI5b
b+yf2E2TcON7lEiH27MTq8AZLJezD4aFbZxGPCG5DgF4//IhRYznyXqCy9FydqvZad8wC0IUM3aI
EXpk7j3EUEoJbrBCte5qsLVen4RQBaP+9wPPvcf3W+H6Gdn5Bkl+cnYKgGw79vZehjHu4pv38FeH
SqkSq8/hv8v4K98KUGS7dOnD3a7DEmRGPs7+uHLhfPSlXVWWgBaVY4AYHbY/DUI9xuBdWPGbw7yH
tLpk51juk8sQu1pRj/fjnol72K/+Z5JvikTo+EYQU+Pgp/oddDrPyrvFUw7BtbuU/HwOW/IP9xQF
bkyk07u+p6nb5/1uI6SFvcoh+mjE3HCrBt+JqANwccPGOfRg3zlZFH8B7MMrBSBi+wRhNhhz3A19
CdsPrcasJqb7zuSk6x32/WMMmDkQufya6A21kAu3x1bNFfLpc6k2w3DQroNKqZeRZpUf26bQNuCx
BTvHCt8v7JHR7hIjR6vFWKUaCbcMStvyv3/IUZHwzYPigZuNIIBOs8+Gzhyp7Yj+KSQgwaXdGsNn
hQJ/FOCwGUA7lyQslvZ1LLw7mWx3Sn843NI+lqLqJJKGlGso0TygVy4fnxxJ/FxEfgWP+tSvvT8C
Gvk0yZynPiD/q5jfw3YndJdzQERT6pdIyoJhkm4JgSkdmVFa4e+90+rmx0KtTxHipioqwhQ7GjD3
8ZZPRUW4f/rEeGaCdM/FeUe1+fYjegToSBxqAXkFYc4IzxKmA9+c67vp+j5PRmPt8N0U8gGDO3+x
T1YuDe/OtcuGUZq5xR6V49rKQ3ay4hjCtrLBOL//n7opycIi4kp0J4ZYlocB1R5vNm4oulDtE/cZ
P/0bZ0Tc4dw8ifoUZQtoIxowaFZ74rWel2WnYKwDQvyIrrrGElD52x6aJ23Ho31ldGIOFhSk3O4s
0swYYha0bBXGVLNd4sYzuXM4Y3UP9BsgJuaL0rJKWLCTbzslvuusnTud4+teAvL1VXMC7nxNpdQW
OlkKwHtSs9fLPN9jLqj6B/K6yU/zUb6Ljp5pie2zIfR8CPRc2Iy/wX8k6amp/ZcnAz+kn5BzgVSG
yCp6VMIxBIx0EN+mz5u9+LCze5zTg3TIN45J2AMViMKkpRduhr7kiXfDomGE05guEXGzODYlMpII
zJv36UGtBofXPxMZR9uHakpDF0VaKi4oQzaC7zfa5/s8+p3nKd9YDpifo4mHCPzOW5fYQ+J20v9K
3zi7Pr50lcVHoikXLUm8eyuMBIIfyB2b9XNvSNsQ3zYRNrW4/nA3Ti96MitAAh4H+eUZ0nqmYvpe
zUShM3ptKpXSHcV8S6GoZTttg2x+M97keKNZUg1XXP7NFxPH5VIXKgJ79KmVN06O+/G/liijVqA6
MwuC5mdSmY56P/h037W5r/EvNgogU0Rapb6nddeaTMAi1UMYh40ggkEDOrZppYEqPCM1eZp1gBNE
Mw92pXOBhkd/FkG3SfOpV/LWzomiP7R6kkE7V0q9yCcpbQuSHRuynHHLDDhqLTBcYyYmnHoAqYTp
lzaNYv7hfDJ3Dg1katWX4HiRCWd0SPchHJyya5AhbDKWsmJJQXExKnKHQ9uAPe2MkTR/kWTVusFB
09Vdhps44gupLwQuD7YqKhUA9L5i4lhO0vfadiChRvthN7Y+W2nGbIENCLXCjAFDP38LIoBinBQH
FFI9Ud2sGaHBVWH+yCkxdzgjffKXpxJVpfQBEzrwFEQYZy1bMI1kVCptaNqZDbJqNfnbDbwETBY8
bx8jfqpvQucsXrcqLSJ+I1j/VhjXkvmNZ5PAPT+SSfDGbkqbaEpEkgamVUAJkMilcGFCZTIsixsf
yGCrQI5SKUobZP/k9K0StZZdtjook+CMpsmPrPD79RxiesiGRfKmVVLS0HjfLFwHSIUOasoSH0+d
o3U65959szgIdBgACds7vQFtTqUqo7RwGtjSSGJfROir0rjWKo6x3EwdeykOP8AO1t7pvB7y5miM
JlNddBxbp77qulp2TrNGcOKAu1iL2QL88zbWyD1yrzIYTLrJHF4r6+6FDZqiVTk2EHxwtUa0+5eP
i+h8dY8EVY1OpQNJiPoUf4M605FCGAdFsplNDvpS0urnm8WJep8gRobB3vFx8GTYU3qKJVPVZJry
tG9uGHPuRWl/r9Gxa+DTZSzhF23D7UUz4L9hcLCra5Ko+DBSaaK9QiXqslhmfKNEhjXQbaMW0rqj
aRco6jWWXuY3LJHgL5jWxZWV0Nm2TZ1PhtJu+LrIdXYyQLHU0vZMmjA5W1uAK+U3IoEBaNxYp5UG
zXbvDnl2+Kq8Lv9qAcf1LQRci7W3Hr8LziHwXW0+9/PjatDwfNDslu7G2mTBkhf++MkpqR4/drn6
hLzTR/dBUWCZOUDtOrWZ0S52fu2lIhQS8q3DfE9qK6ggc27RlSxaYDljD6Nnm2ePLc5P/s/uJ65V
6WB8lJtpfLEdDI1taU9L3eY2dmgBa5NyWWDThrXvAgqYdYPY2zruNiZFNZwajqFMzaV+ermh3Afw
g0WIpMOy6RC22g2GLChOuILUAfAhTq5+WbI2Hi3I0Pd23xfjKSy7GVcFUBO8f9ItcJTG1GGL1eNh
WBC8mn3Pjm/kWyQrL6i4oO9iOFS2cxDyAG2mmjUdJ8IExoJcI/Srvihbjmk15FnbTEm/9qmVVB+v
xPThNRxElglKcqR3OnvuVUOccRZTUt3UgxymmuIWUuj1m60/fIOlCvmurQjeIqX8mJyl/VYHmcKn
YJXZGkTLzxlM5iV6e6FQ6f37Urs9EXPsl4dB0B/fLMtfa+54Kh8arPL3HkUj1eC3E3KLvFgYRU6m
W+09oSm7MMSMpeZAcm2/sAVrpLYf46UKuUziPtyAUfSCQDKKB3k7xfY1OHy3xUI7EYIoKJ5h4pQe
P306BqFA/ugy4c8xeEONaMhKZlh2nsEn0UeJ/lYCD4p2UDknQQ9LgViCU5wxi5Kt77AU6FG784mV
6FjCeNILr6VBXb1aCZ+KxQ7vxsxmPWqVrt7L5g7aA/pWTykrMmV0Z2yYUgu0u87T+DnDRW1xuJz8
QjuqhyFiMN45TDWtD4dS6usc6LW2LFqWcPR7YJCYgzkvJvyoI55XavM0cb/rlP2S2EDUSh9xNT3I
ztyNmO0ocLvCD7zMQfKmILNusrTMtcxmuUU/DrK3QKjpgj2lM2iftDnSWGbwlnLUKVfCU7yYJ1hd
pX0ALsV4GFoojttgYNsdqodAXuhNwP6k9jqohgxReJ4kWWkWO2avKmVgZEWU7/a99yH/AHFMB6Xw
Hj6eYmjcZlgsV81r4w9J7EzrDpcclUcoR7/w+F6QwqIqDgFV/MFhCCAE4xnoyg81W40iWk2Usz8H
TBzukSNsw41sQfsMV9UrVe0lvCkFtm7vdJJVZoIhYkOcKSyqU2zyfyT+x70yyt0X6X8wmidhIoZi
sN+LWIEEpO+Q3k8vyIJIY/ZJ96hIy/dMzjTrDZnJPyBAivnEzVsUXlgU/rbDPE6GIt7fWXEoT/ct
+TjmtZXBPFMOVgANPZ/TIrWqG+JOw5U81Hrp9cn8Twb3DEfwEqc2bewLMZF3kkHVmkzjSRsHoNtp
eJ19tnrUicWXUrgvP1Vf5VLQiMRsCQdQ4+hh0AGLwej1o3nC0g6r3P6hSBzV7PeD1+rIG9WC3I0j
HinrDvzzUM8V9QBPI3LcQ7/fhASB9qw1IVg+WaPgiAlRrt5w6j9Q3SSWvy0adf34vy0gJXychpsU
vMuIWdsjeHoS6Jtue/LNxZ3LiTdNxRoQeenKdxTmrZZgYYH3eN40NFv4yaWQR370G2+CvpDuxH+p
0tcQoU14MtwIMkvvCZqz7O9+dgbRmRk7rx9W0+LwwjT0fgY4YVmGaV+ubST2B64iwewIBYD3N74m
lWTNI+1O5ze0xNjyDlpDWTv90v7URhMG/+ZjhX6SB0dh10LGFHGTU8NGJP1tpdsO5f1eXKRqY3L1
cUYxR7VKJgkFbPSi5ABPyIPMglPdy1RnKu1u3aIANesLnot0KpnS11duGUzw+xqtOOW4mjAsx6v2
GQNjIOhsyQHk6CXLNsy4EllzAYLAdjE3D4YUkY5Ogj4he2T/DhCjiFBvSbpr708+iwd0geeWCF5g
EzFOtTmMvPW0ZeIrTolo2+F2eFJjhNuBDowMejbXLca68PKr/9uWkFoNabvpLKJ251jF8SwBtLj/
2w2KdGHU5qZ2ZozW+igDPFLl4Gme7Jz5eOQ9hE2xUSGr+1N9sUaAWIvg/OdnqJVZDfTpDBPTfBte
xo4YfMkWGPhPNvfMJNk2mvy2iEXu0WztKNiSGgjg8jphGZoU7S7n39zaWNSVp1S1rBWIwXLXRJaM
cQLu6DFbsomgEMm90oQITtEdr2Dx8xSwn+EeJ/vEXHURf+d2FwOZ1AQrO7sf8oxwjp8rT/SXN9Wi
sEHA/cC1XDvN0YsmdXv/+eFOfE799dDRxfP7tSYaMxaZfdy7PkPIRvNeBQ9HoGpgJxZE0HlNO8FG
4qcL+XPwZggnJDWyi8rFopQnIAdde1SOssoSbcZH202xhRESkbo2WLJjgNmNC03NyjZqLxR2mpvE
phQZdFsbNXTN5ozTCZZDxmrKp5tx7CmyfWzh0S9hY6OxHNQnv+5l2MSGTgLzsVbzA5+3DmKIm/Gf
T4jBxNvpm+FufzX76nRo3KUam1pw3m59at/jg+p1pvTb7afcqPqsKi+YgjM+f8kKmcsVtbjEtZoh
3bcafyH1eJH8DJgmDUNvo3PLg6jw/qJNHheGmaD09JSOQMXnQBiFXpEXwru/h2hGjhwgIpk7cpWV
qBfOkvkjTXUJW5ZC5PjNsZR9HIEMubxCvkfgrHpPkKxVxQkH5BO+a3j4DeWB8kj3whv9JXIx6uxK
vSLqv6r40Zk/UQ/AvsSI45FR/kKZgbuuYOsyHhIe+dN0vBEzMm2ieqGT96yOxHFkPjrgu3y7sBF6
GsoVXPJMtGcyyo8jZBp9lCPJM0yoQM5Loaf04JQVmxv8OZ3B89hBWrXjZOx84Im2sLSB0YI0K8gR
jj9KEGNGyM2uKK2kbYor+VrxZCVW97rUPZnIUY7D84IVrk0k65juCEBzeSRLy2x4HRH9uIweGKHT
6WY1QxTW2Imi6kGZ3NVn0pO1wsIz6iTVCOLBL7osdUef35pA+GV0t5LGQBYzyyl3shlEBQrVXX2l
QP+bVmk4PiWGsVuzUwMz4fy+VvbD6ws+tgY2JACDYtEfNy5+rYIt6mc0mBfz0L9gSOYlqmuZnes9
ZD1F6NlnMhyrGjtMoLTSeoKbt4naUA1W5Xlx3WGYqG6x3XSY6H2gKzcVohDxJ6RSCu+e8Gkr02pN
WLfpozNo5UeudoMu5TafHw8LGHLomO7HUItZonv7oirOwDGvCpBxWnemI/5/kudRQZjO3BB3GHJ1
fEB/tvn4HMLTbDh0qIWxe90tLh6beixYWxzfloTcS8ycIXXZ5B24n20/9YU8f4sr0B/U5vtOTx0j
/JNJp0MxCUimAlTiSjszqk8mgjtXMSBQfdRomkpZQbSoP6NOdD9mOkNljcKeoCpZC5opmENSyKEk
HDijlKAXCeSJBmsV/1YNUH5dBryCgAjtAsUcZc5F4DNdFLbDKNHzM5Cu81VOPJDrEPe1W+4/s/+H
fjgsc+fB/rs/k0BRJKGkNU/OtihLll/kvO8BYcdryNQ5+Vv1c6ylsbynZgI5chMhkOz4taL3u9L3
CqFOqEPZWaReu+l6Flvo5L0EzLYqnHZ780N9xMUI6hqnsDYoN9Ng/KSwPil4DT4j+l+1eQIVmYh1
U1gCUQvJsDjLaeywBw6rvpElEhPEXTOV2ZHueE8dz0VNhHRmyW8Fb9NQNtVxKVIRU5ynM1UakxZL
36cxIY83OmKdGnn8rTqFhyOJvHNGP3Hnz9fuXvCD+MnthcxaUpjUF+cb4XVLVRw74Qyoc9LwrNkT
/XvCpKErfMcAn2HAdFVcNadD3DBiDY9wCMHTTIHj7r1V8+u15zsxIldWNfWgd2tenK6J/v67P/86
bAAPTK7XU6XHPvRLxNvNOFvgnBa/Nj1n5DDVGfmSbixZshLcjGvAJYFTSqx5nxdFKzYudRRM2cuQ
srATCaxPhCoDQd1tkkNwC4ld1/2lXXfAnYVXVBlRJxbNOeyhXxEptjXJhhMd9W1njCuUS2CWfo89
uJoRjNh+oSpxkNJgIhTzOo5kVATZTIz9dgYqUa6EvMuADbYu40CD+OMcbIGM0/EcFVhR+fFr2QNh
oxTmokjaTJdSV6PtI4n3rHDAlpU4kkiP0tnAQ73WE8wP/A7Or/ygZ/VLPmvWseTxLCy/qOAz9v8t
l58H+GbowX0q5RDnrJ8HF3NWHiLrm75L4ldVDEqMAar3tyq80AbBZnJ0Yq5QEqiTqOCPXQMKfl9n
Al/IM/SPw3WfbYqbp/5/A2iyUVHGLeakeafk6vzk8tvEFsAfcNld26XYEVgycefBGlfsvo/nF7kr
blqbf/BfDWpduWyL3amDiRDaQ8L+rWS0kHgs6Vguiwxy7rtoWD+deyw9ehO32+8h8wXmMQkC0Gml
We3+PYwWPyc6HuoUoJ9CmdmdTwXL2TeyAbd9ERd11NQlayVzLT9XjHkOfPtrcTBd7QNZfhqSPJnp
xyVaj9uvJNTSpF68MjC7Gjw6nxT/4F96REGWH/R4IGT/4it4JaPHFJulIEnVj7/qzR33CxGsc1D6
XLIuyfXsdjhvRJVKixdEaq4Vm72MlAWflrX14j2v+hzn4G2K2LK5i74hivf6CCGlMYl6H+BgcGIW
yYSycS8tMBjc272Br+5CzS9CdVPpAvpKQp9iuW/2eal8ARQw7cMOM7cehiOk3Q6ZPmOf1XcB4ti/
MaZ6S2XtyLfirCExvg/wW6dd5l4TQrbN5fIdi2bA9EJzaN/5W6Ck4IDnMTGhGq9xra9OWY1cBq9W
sD623p/ETyQ2Ko6TD4LixZ6QW/F6D22vsP94kcmKy3vA9fntxDk5t0hUUjB0vcRvE78OND830ECs
zI91aGV40gLtHyDdlQEhocwcDAFqtm/rOa4lG31mwBZWcLJ06O3xmspNYFIV6ueBsR1QIziQL0fY
7kMMlyse7L9J4eipIaUaPDn/rTYjRPXFBjDOproJKQYZx5G8bOwcw/Hs/UaNEi5j3+Ab4P+aZhNY
cWItUHuPkLnVXGawmlAH++f7ddIscLPoHUZR0tqiFHnigtN91I4BFMbDQueegZHYN5HUmUa/bIW3
FJs3DNFcxmKsXB4UViOqrqsNCjXHv6P2FZGa3WoFyV0wX2O2M00ozsl/l1SXHkrAv7HvHmj+/obp
XnLaGZBdG6pME0d5z5YO3xqNeO5XkOMtVDGsDpQL9syQI4ZD1pAkusal5FaOdze3yoQFVXgDL6y/
EdQXDj109NbsSAidcZQi6rUwF6jgN/Remmaw5gwi1L2l6Tv94aZHpUhuqTHqvCO5ZfW67asq/VzM
+c8qU2aNZEWYfHU32B4IiiqQ6T0SN7Nk4nMI/T1g/utcKxxpPOIJ58QO2YF8IyZHv25GxyvqAxQQ
9vv43L5uSx8h/+qttFYcp0bsV6iH9p+NFgeEYokmuVfroScJul/AE8OwUBcUxau9baROha8CQwmk
cRYltNEmVS4Lcqeny56HuAZkDDD2Va7JpVPvQ5mw3W+mZGhnSL8VyEJko5F9iGe3OqAPWnouWyOT
EqxgPI0t26M3RGZRsJZkuZuUTxzRqJXdrqRkLvLZsBDEmM0S2L8rRZDXdkO0ch+8VATGly3x3CdG
rwM7ShahjQuNHGd4ROioT4+MS5rJpWphZrcw5aaMcQtw/c6A+RMmzn2Rjw/OIG4cNcMxI/NaI1RD
mzKaC2c7sLBqm59KfWjNIBYz4DYj3N+yXcambOTC90/y+N67gogvYRr43bdedlGGzVMSMG78/Dw5
KOqYXFo0V+S/7UpE1vtAfjSBpD5OxsRM5YczvmLFpkLmsmNxLG/JyAsPXqEcfRGGQQTqGKCo8ipa
SZAuJZDUumSC5OdwiROZsfjHtxosoQH/nbMRCVs4DQDr/ek4cEYAKoHcy6aEYqEc6+1isC8j36Nc
tBrCeIANTBH4E5+7ZrOFx1y4odd+Uo+Xu6LTFWGbPfK0Ni7PQjsZ8jI036mwm0VAdq8ku5UxTykj
8DXlRFksL+oIUVSXQBF6VCpqs5K/9VN84d85Q0vLJK1bkulzdSLsf0G4E9MU+5dDrIvq37+06F/w
eN3d8SaP2Htux05hDIMHAgsHMVSc2aguU48PKz+fb1Ylwhi5Ieug4EHhFBUQsl8A3wyu7/jTcxBg
KiREeg/9IlR/RuS/OZZYwsoIERSO3YYTlcXBH1lCIRFIWQEJnyri85pFKtnGm1zzRV5CdoyV8MVb
ueLbWq6kci3I6m2Wcwe3iAt9uYbn64aUNsF4oxfevqZdY/j9hdADZMcInxWE4/xIe32t4jVChNqp
SH2AQZPhuJimPYqmNhCEqXGREBuDMMD8KEwtTxUZ0T3aMxbQD8fQix55E2KzyhksTznPfwoE3Ys4
dAVgMnuj62gAAlRvEwdAV0Fqzu92WSoxbFAAobUJwXhy7uGosmFZVVHq4+/522QGsNVwJVOll6B8
HdHMUDHSIwfNJexR2ofKAefAqsOj0LlPgFTWTF7Mi1kZiSS3M80i7p8dGrNlJ3qPVDzxR1SDT3lR
IpPiKvz+7L4fOK3A/cbx+Sp7DAzkI64xDCi7G1pjNM7sP0kdtjL3T2mTgEroX47Apx15OW9/gLDZ
IwPbjUgLxwmCQLd/sMROYK8qnjWOlKFOHTXFoV+/JzL2sYEkGRXNbGJXO3za4r0e2WpqcG/y89sJ
3TCLjhq0CcT8MPzB11xCClFNhYYEsGfoADCwqif66LjJiyGO0XGePbpRrXjh0ZYShwcHUDNIVhcU
RNZt0KeEqG7lR/A+PZ2ZeMHM3Em1bCt1lL2/ZI+APR9ef0tP/3zZRtqs5JghbC/VoBAHXA0H3Xsk
wL9WKA/4G+3y5X+DjdS4vXWU38cQ6moFa8TBQha7PNfNWqIDVG73+9SrfSuwxOSFJtIv3vQ+AuvC
+NrDLjFRP7uXrdYsGvBR8xOOBLR+AXKJeka9tSYLvBvHVSZHjW1OPDHc4xJ+5ne4Tz2eDqkzBKO9
14I80N/JH3r+oFs5i/KEmaTviV2uWz+PQ0xoD289eWHJe52FjXcYraGVDsQEiwo4yfEGkh/LcpTa
GtqjN1YxF6BV5GMMmpeQSNT7n/gEGeam3EvEaOHuJPJY5wfCrD1TY71ma6Efd8X3HIG9c53tvhBA
NNFq5gpBnPlaXppjJa0nDboMJaTOaJd0P7YUusSUG4TI+flLh+znIq1BxvTtPPRKwRB34tmWnIZP
fRBp6qCQHPtry6b6Ax5KnD/Cdkmfb1wyMSV0isYKtSvLHZlXvvgIIVjlvnQxZrLkZIUg+h7Xuo+Q
+tYLxSxA++uaKR4IOGEKdO5WViswIngP5C+f0Ght9Befbrs0qEuQf1f0yTJYq8rhP4h/qMi2eR/B
FaLHYDxil4DGIW6TAA3LKA4y1kfQsCn3iGfLhBtKlxN5wQdhBQPA4MqiHX1Ql2LGeXIaOXCIwlO6
8trkuRhKOiJWXnTq6qyUauvVs/M2fjdl9lvNlEhGdlJhzDdhjz1202430mZI50nUT2ZICAjPCD4B
2YL/e9GLW3i15wB8F0a+lyOMj+nYEoMPi+Mm6onqw8WQdNWBkLGAnwoLpEVtpC/gImJiFR9xo7FU
VPHXtRogfglh+avWLFd+spHYl6Lpmy4wi2on6Jrk1W6LsEeJupYT7d5lx9P9m82Ifb3f/5BLMmaO
oyxUb7YPagGmkNrAHS7dcG9xTIFGVKicVPF7ySRx4g2NxBgfJ4XeDorhiIWc4XLPfq+C29XX6/Xa
4tv1DlbnQegi68gl+sHk4xa6Y1EpfQFcit8MffO2UlSQV6mCpyLI9JSHL1FV2es/MAHcF/APUQOe
i4Qw2mdjv0LlOTjRxm0VcPhcGSXM2VWJWBya1UidTDlAirPkQxeCU4KJ7kyLaxtkHP1RP6GWOIXp
dR+ltMmmTrs6zmUx1R7flqsCIHyfg9wxAzB+MwNH4uz7KVzshJNpLE/OGQWqoGSnuIzPQ11LikBo
8wWzYkYDZo1nt759qZaAgMaatGVnTOw+JmKu0PMYqvQw4o5PT8/ZGouGTn7ran1OjzDXSGEI11pc
6vV7tOaPTYj/ACidmRsrZeERCjm13la674P3sMENQHqaRWvsomZA/ZeF6lFvXhyxHrrLVvX1H1q6
hLn5YMSA/vc3rNbrUKYJ6u4Iyj85PK6vf3I7Ig5fDkqC6Jw3hIhayOnW6M0sZALxGFy+56JliYCb
xbmM4Lpq5t3FxqY46GzJ/+JVCcGf4MDZrtyNrKOUFt7VdZ8hwEQuAA89T9/a9ufgnHpN0YfUM3dM
GHZRq0zACiYXpgLcQmzeZzSmTqnArly4jjS+scvkMqt5fUBv3MyFKVnvB9p5b29MA0xvDS5A1MQ0
Aqt/V2BEC/07ILP0Zb4srZMN68i444nimhfYQY2C6f0/GkkTkVb6hML3BclTXHe8CpnA3n0J9wnc
4fVC9jMeFOAdfUZPPAUBgdRxbzTkp1gQAsW829NXFD9FR4dTbmhql38vGMQ0VPS/MFSjdKuEfeSl
rccP/plPntI408f51c62l8xa3jcQlyfFSIvU6HweO653GHm33Gh30fSqbVVYLFWr/rANvpzPAxdC
4GFjqruR2nS78sPoMsirBgMeIfHi9BZkoxarVYX1Y+lyZ7zOBi4ZJnbg61e5YfYBLRmIKKVMZNSY
yVwZg+2Z+HlkeasTFFIQkOiyY/oIiNyIvalKs1+hBLRUJ0/HVwUC6NA5boYs/ODjmeB+O9MWLpTY
QK9+K8yZowpxPMJQiQPJXb6SfzbxZm/E8a4nK1CRHORPlLkMqhM0/JQZ9WgPt/Ccz+GlLbioZtqf
UZ7bK+L4YLvIqfuOnXAGQBx3lE/hFhMpsMv2MdtA4QSZkigA9DR4wvxvdjJHJnY4W1SFBIcubaCv
66dr1BPNIeRIXCBbOMdk3Lovk6VQB15LQbIqaaDpxWzJhWT1+414hgPzEIhbX/itysDkUjzRs3ZA
KpknPbbAHN6U15TK8aq4nqdL3Xy/DEEPgNrtYb/LbDX6qqboScvV1NozdM3nUX4xx2V7U1SmC8hZ
Ocve3eOLRtKsUIqMVFbdjvMzU7+az3DSH+Bz+lulH0rfG2HtFvoI4UL7iSDQm8kjSU5CIZJyxmOB
WYG9zawgmdDBlTplIyDUigtgyPgEFMKY/BY3soflNLbfusZr2ENZP6I0GivmLba64/f57/BwM2iy
j2ikMZClYt1CviZacWMZXi8WuWNeZIWXp4ibPuc5VMbB96PHxVfj+lt0M9EXq+C0IaTDCB0doL7X
Ed0Q3MuHjBKuuyxWuPuhniH0g64yxF5i3GO+Cj17oZhXWFPfkjl7yoZwid9a66dCi6bqBsu37l3Q
wVJmrEPhuF4X/AJr8iRYUCv+b+ZKOeMv2dDo6JmSBUwhih1uMvxYz+o39axlAKD84PWOxz5lr4IY
rjC+Rh6/PzOvqD3CYB0xlMdZDDU9qhcY//ILHdzFHPn5jsb5OIlEP7FhTe1SC/AOO2uY6ZOEeViz
nVvASSGSfZCUri5eY+BfpioOHBX/MK98+4CYkUNJfUzAqGhniGJ96Iis/M7aXnGCCoqrZWIHZTbU
UYOV2Aw7tAizJ24YaZD0q9uWT1c27B5L6duOl1p+nTEyg1tP8Gd+iWb19UAP+CE8BRQytCRtDAEt
xeaiaP5dB4KF9rO0MC/45jgVV0ii+QHIVpaySmdMYl5rqSEk0Np/0s7qXe4opdq0j7iL0mNdToZR
HHjbBZxlf95Sb+4oqtOT87yjPuvt6Z06+X5x+ysgUoItEJ0tqlDjD4E5ndNzmYhWliOigI8QGoMK
MLeDYLS2qR/5Tz5nWLOKn4wwII/OQtYEu60WP8iZQbsPobkdQBbb1saEaJNMFNMbi0FmQdQjrEw2
++lRTNWxTIAZ0UM4R+DTzJWPzMyylteJBu+ELYSr2Z4me04X3fTr5MSNAmLlzcH7vQeWXDFdjwv2
PJvB0tyr++yrQcd80UKkEN3eC69fi6TQKBmbl5pFPS7gMasxiT4yZ9ZG50qBZTCSDaxpyeApry0h
NoAN+hLIVGH/fufX36F2THNrb88V4sP5dsuTY7cc4lsQFdxvl2AXynwUvq20UaIa+UqZewWKndVu
nKYLFsbW4VrYjWRbjVkUwufswsTYrFGT2bsZYVutACIqsIWq9WBV0vc8DHm/UlWUZrq2gZVb1B/J
Sy5GZqMoVwCyKpDp1fUYwyoHrzpVbxI4Mlml7P8TmaV+fWff0pZd3oavwPuEV46Bv/6CdC1hrGiH
u3JmjP1qAQmYpSjZqJv9/l6lReK6YPRnYyiiszDE5ncUlerNR/PaSkwvLLHK28aDLMXt3fTR0QXG
o2FMW8Y5UD7hG4YmuI9CXCYCem0ySQjm3RB+ImTRU7kekLZcBLTkf34xY+0PuPh9EA8fRMQOjtjo
JrdswSZqGzlq6JeDKbs81/Iy0UTjlmCEFZ4G/I8BgcWPfnG3UegQ/QSljnuzeUSDFXe7G9HJzrYg
T3tHAVO00mbdHJLr+LwFkqshiIz6KxwpzY+kV6B+DLyrBREqKCioeJm3Pg8eeBgKa+uwrvczAZ4S
E+Hq2nRmiIcAQj6nGlOl7zvLwMc+rYfYjl4UY1cK4PE/VPv4SsAKc7zyUhexx5vulBmHRj3+del2
4yWt0xnSCaJtmHlVNKzm/rXF2zOw9nmNbl+spsiTDwyFJbBasSybHfKXm64V/+sW8ktVFk4zi7W+
2ZM2hD8obkmsiegEYmO8KqOgFftaNlrFmgNbV3+AXu3gGQRLus3HvZkWO/NWsMucLMTt7RHW0OUy
b4zCKxNl7LCeu5K99ijqEI7EMOALmkpUT+diWO30Bvgk/HevtPgSvN+kky04YGaJaim6KC+0LByF
RcVfWN+ZD6YIntrlU0oOf8iyKFZM1FNsDO5wYUn2KDEUxAb9d7mItT7w09ZeEujqtxg4c4V2BP8a
+2AWTYFhIzMyh9Q5pPYbQ+tix09vKBUg8BmFR9Tp9JTMTHc+cw0lvYbxF17hb1SwmE7tNLk21iYO
1FrQYvVhAVX04pndMJHwvgyQJYpKRCmdOM9yDt78yGyJ036WujyZ0VTkHV+fsGqD2aNFPEilrB5o
LwFkgOjVG+NN43WXu7rOSWXImK8/HZK/bUhHNpNitPmWZGKsLgu+FdKEbqZbFEMpivkEu3I1h9UO
Ta3Bbgf6/CWwiB2LnmIyUNG78KP1cX84B2WcpyYoZd/JxuOR2C7uTfT/xsBo3okrMsDC6mmIcGfJ
I3eJ425iu7y+18UhTd7L4D7KRha1pv9k3HGyOrRGXPj7dt8+OmZIPXD0j/35KkxDbCjlV4tF1USR
oYX+CT/jD46qW25OY6TW9zLeJVvgStEz5YVbOSNIR5bkiHuvIlzeW3MfWXvi93h6nsGCHQj+9bF1
orOJwGIdACbSdje0BRjYCUT5r57e8SvgbGiBN//6ASm0SXOPF1C/UIveVyFKXTnezb4g4WFt12FA
XoDMvwoBO4i3X0MmAbhPmyreAhc9f3tQW9bHnaX9iIzsIXZ5g2TMGLtQ3pzIXhN1XuYH/6YSCq3T
nmkA/ZHguYcUz0bxSs8ZwnjOSZF3CitYgETX2BWNBuCM7+VSfqbWZSvtx6fOkqXhYcfQqIDvk5tB
96outEDM0koW5yyMt+JckgV14/C6qQtt16rP9Cx25csmlAlBS9FY/R8QgbYzzemJ65YYYfHhkYt4
vjlRq8w97Arvr13Z1ffDcx1U3RbGcnf7k/bTarIYhWIOtEJ85jZV4EqPBP4brF4C6R2uO1u8LiHP
xGgNl15UixSR0Mgw9yLZFgZIR+tIFUaebX50r6xtd7hAAQwhAGOUJbPuwPOGeKr7kk6k7KcL5Umb
t+3uIbllgNKK36vIuSe9lnIm8Saq/DEWN2n8AqMP/6aU5TUZwkmMfCuYDhDg3bOSkSGCdm7CQaeF
I0T5mYSiCxoVblTbH6/3I2CMf13aMBe4ZCElq1k66Cmf7GHeX1dgmDXmbaExIEljDOFMoOfMSPkM
+Z/MX5vr0X2UMChWNcmvla629IHQ8KkOR8zIL4V/DqpWmYzzm4BCg2dDNJjjmnyejKXqc+d37N0Y
U2fgwUVJt1y1d/CkTg53ELOlslZMBVOO5YK6s0mhScXgcrETDbns9k6ncum6aeHmitZabm4crJaZ
DEwW8a3xfXe5pvDTN7faedmhsH3gLhjfzJtAWxfItWIhOQ+88mrnTBbghQEMY/9nsK9qx5GaLQ5Q
sm4S7J+DTlcIuPo2klr+mIoccFO3wPVm7jTI1uhLH7qBbSJ1JzJn8ZRDsT4l1ozZIa7rw7X3cYtr
5kzHpYeXAlHGewt9IQ2TX36o16au0T19k73YyZoi7z7CrBJswIjcxyaXKf9x8YXvZNdpvnO/vMVt
yHBZrFl66aSRd3unbm8gtCDlq0kJlQoOc9T44Ue+iwQ/eVZt8Cm4BaUzJUcCsEMh/SLuS1CI3dCD
xqdptngJ5ezVsf85R9warux94oZNfEYds6QHDtMmPmJA9lF8B0GYmAssADLHw6Qr11HTd8OXBhpo
c5oL7VacxGKKc1SCG+Sya2BRuT9ea+fVyHgwU8oj7KDRIb7csZAeRAXk1kUJfajOQ3SKFoWOqN+J
P/SKtM7GYD2vIHRnw55iu7XpTGuMFiSD+gW5yPfM0sPohqgBpUpp8Ta5PXEwaHT7Bjj+P0yyd+gO
WqMIyGZ2V8i6LpJoVJV/HrOdEVKO7RfUuSPg9MVZlQNLRd6JbI8+0f2+jFgizoBtMQDlPswm+ONQ
x6yUYCfuiFUWzM08eRM5MF6PqmwKKlUOqFu5t8O3Xpk4xHb4NSy7YKTTHaDMY7Of2+jKfD0jRQss
NS64uWo1BT8En6pKM37Nc8VGLkqUz9v2hv6Rh+7pEVK0s4+JXGNzeXgVjIA6MI48bkWqFnHir+db
G7emAa/NAJ0vgHWmtNYHD3q+yMap99R5mrgTvL3HVE9gTIYtTVcb7mRjOaQ+1bDHwbooFrcabM+u
HPYuCSog9gj1i3ivJzJ3BPXdrQ5Uenu11NCkkZSyZqcWh+44P32IpP3N7mOX8nAftO5Zw4N66fk2
T9d5oKqiLWMjPjv0ZRBCPvDRh1OAx5p9iGE4fSbvMZZ0Iru5JAIP7N0W+sapkguqT2uq3l7k/NBP
ZgfDhbVXyx32szMfun5YFbQD4gxAZerz9VDH09pKluSDNCtaCmmezCPJhznCdr+tj5JU5I+qHW9k
xk1fOI7aCUDp0e1ZZSQgzAvnTJbGx4KLjO6T3SVs+CZtAEn5pLKWJW+M7EgXFeoYDWtn5SCLFGrA
fgdazZny1rrKkmbJM1nU5o6NcYMWf4HytuK1fpHDXEaCHDJgwLiHRXoQHtqIKFdRK2MCEnZiP1Ra
DfIOaxEUGMWThNtF4i4JsHNBMXKLUJ1jxM+5mrTbTwvnVJrqeQ/cpTLocHRN6nyff1moykpIKYlp
5UFq77P549aQyrbXaxgXaryIy+tzwKklKYDnLnblEZdN7YZbjnzIX/pucNvgVAYN1QI1d+J2UEB3
bj2p22RQod0Rup/fh93jyqlghqKcF47Fprg/u8C+wu+k4fbDV79UeNYXhX1EKAvmbWiRt9CYUSKt
0cOVr+BbjmE3OpUIBh8S3NydXJCk0qW842fNZ1K4eV/KyzbMTRb4lwl4s2vwcKkz1VyQl9RGi5ZJ
rMf0ModKOBnlXerOsknKEv7UdtSt09C5dQznMnUBlfyUNoDbs5UnwHAeYmggS1JTQoslPQqBnzHp
gTr2uxUB7vswAgfltL2QRfgJdUao0eOZ4Ik/IHENBMm9Awy/DqA08HTsbak0mDhxcmkM10SvEvJl
YFsCShUztpT9exbAZRYgqxHA7ztwFyyxxUpiAm+7o6+HvF5N/yOGVvjFOcqbOA0FVdv+cd3sjFPE
S0gAQaJd4Bcz6VnHsL4+XIrkPBfiyiY+Imk5yO68/RPpetX7GqEZ5wtNfQmBmUHmjg7azizvDBmS
Iwqfa6MTyL0QFEXskKMcp3Rfgw8/yfpUIT5zMTn88QWz9Iml9aQxUyUhz61jlLlweLwttmw0OYYC
c7HxTu57YImdsz91Q8B8GcGdhG8xZ0Fp8TY4iGATu8RqwG1JFRjs33h9PdYP6ksGG/D9yhrgRTuo
ruEJzwaPrRvsBkpMrWhoQChind63XvknJDwaQoUqMe5FGrgr2WktG4WxuUIeHqixoiIffPPuHeyr
hV0v1E5HAzON/J+RBSHhXw3H5zDhWMNPApxBfv2sJlKZ6wcXYahL5dCy/oKZz0Z5eMXIlEENW8Cf
MmDeOxIKiP47VSw4s2mZTTTTK33OZlvh7t9vf87T/2P8Vs6ROdRbO3ttC/rDP2BJe/lFcwFBwpuE
8b1AHxDf3RAGKzGN6KTV2wp+rOsPJmzk8EYs68B6SYThMhUT8K9fyfiSxlOI67srks/IDYtNuAKi
K87NAJJ9ZrjYX5NTwUwr9FDlLYuQngtGr1dePIdFNtGf6XUXVz+/h2FqZIRYMCuAECxJp1MuGxLH
SiqX4Dfwqu7KiDsgbrDSV3RjBesRMFCDJF50GSXGSj4cDWjsrtJ6lSj4Z0W1su1kFXjOw/GJpuax
JBbpIHNJw1T5SDsqK0u2T2g8K58JVVn26RpuKgt2VKonBv34PmlduOAjLi6UHLlwafXZhaL8wbvb
C3muo12f2tKvwmkBl9x9pf2PfoyKrmqXXK1koNX1zxQbWUkjF5O1FOLvfMNcNicyuZMWCebdpJEU
2+McHtOWB6VObSaW41/++ofAhnPaWbStpeN+hL08MWcI8st4MhAMHXw/pksLhMnbnPfHuNy3sKbu
9iikODPcFHSy/1NTfCJ+lcSzMOmNtv7jDpRbVMDI7arYezbh7cV4VQhdLAjDrb6iX+yhW4J/m4D/
Cfo9ghPhmuM+C5osjiVpcjUyeO+7RA/I7PKUbCcaxknlktUKjebM7bP7VySj/bMQaFytlzG+7mD0
HoSySXOSjlv3rp65G4Zf4ZXYDHo2XqnIK8+e6ktuFkVeWCB2zHjEA+c8zzLTxEY/g80E5jtlJSGu
xIEWZ5kXj+7AM/nrOF8twSx9JXD85ufLCZMlYkAb0QFZGGOuUXtdU3lHrJMTPHZNs1FhOZEwXhoU
GCEsgolAuMfFemW0k9Pz0LDwl+i/o3tYgv1XPQHO0J1IFFj+pKqH5Y2lrQ67kMVaoLm0JkBt5RaK
bwAG7p0YY7jjsIdJrNffDfs8JLjDW3cVW6ano5k6NrXFPVBhzdt5OA6ZUNEOAMeGMgehviMnc/WB
9ex+gEy1MB6tOU5TBKrtUJBtgxow5NY7A+JJzNuCccm1S8bQfzEeinw7xQhQFuCkPGNcdOjRMvDS
kYg2UXnvyYk82TEPJ+U44PKu49pAQJReLvvS4yHvbq1y27TQ5BbF6pw9V7AvzLJFdWfMxZzuO2lt
aOdTieg7oQ5fvwcOBZhEZlNZ+31HwY3rk9FH/+8wUSb+tBrvBsS3L13v4H+v8lRK6OtZl+XrIbZs
axwnRytILD28v0hLlx8QRVzdM/EthJIZBmn/K80oAT0jNfYRU5+kpRv41MxXTjAPl6Zsy3vGT+3Q
Cdaz2w4S89iTmVFlQ0FaNWpDBy3AJwC8krZwjBKVcr1o50GhNmQ5yx8/gws7sEjdJ6S91+7TSiy6
SQH57zqFuQu61kffkaGgpckese1W42V/Zd9CQcPov6RWAoV9om+uwVg0KnryHTfcH5pClJXT01qZ
qFugN+e+1TG955ERFLMPE0AUXRDaIg79HA5kHdhorhipMmhOdwsIGPv4y178kpVS6EnQQBxm51eo
ikWsgjp01Zz1Ke2cX2Ud8viWf+7b71tNZXQ6eqf1XMSeb+UMFTKyLVFn0zzEeu0ypC/MqwBzZjyi
M8JpCHfZkBVYkUEJKiq9qqzH8JQTT4bNlkKYIAaxHSvW1RU3MGXOZxhplmS+Y9oSS6sA8hFRyD1F
lTOb9o7w4on9/S/jFDvOH3iMgefbYwYQtJDVOpQI+Ga79I+CzqL4waVTRzaHKUaBtkKTyQNOSttV
iEjE2lfz9BwiA7n+URYECR/5wMwivb4Ff2+iL10XINnervB4b9l7BvCYHJH2ouA8HFI+vA+MxLS5
sicv6DomHszsgXQ9x+2xn2wezZb2m+VVVimPrgnW6BuGNF3Hq8QHK7JpSglPD6zsvrQjq68m9clI
X7BFIEQgllsv/+nhUj2uFWgWIzOhQ3GNGA/lQGMDT41bnaUTfjRSqLonGWLnRsGbT655VyGbJX2F
PyM9d3oOFuKSB7j+/ULv0IXjYkIs29/rx8KiY59bcpK4a7G51qwskvXVlAwXevUf15ZzNlaOi+qf
lGFKdae29xY7Mr+4yvSWJPVnvzxP7c6KLR8ErW5Zrdc/wlM3iyoLVvmsVB2Rrj8+pm/gt0/eAbhE
5axmdLWl6GLIFtU2ewB4ACC7KuY0/bI7wKs92dSmlu7OFfLAt+UVqZgNmwGhpl1hu72XhPn9vVWA
fodAgGMrbz7tJ6wszpkLW0iTyjfGbeIP0evQy7rfza7tFfDr/xm5FIZdZ5xR2EL6XupYNWs7fEtu
feVgxAjtfzSxXS7y5XoNZiKydull6HNe/hso2yzjvYk8cMiHKLzL7Go39feG3TWaX7CuMNu/gRNu
vse/cRkzqaLBDC4QiZX+cw4qmZiK008nMftOBF5n59ZNlfVzX3/cYno04prPEUgRfm66/b0LxLhP
FTnqrW+lIb6la+i98APjiSYhBB4lfq1TgvRjOvA4EAmqjmr/DpMwT2oY8qSGcgkVmuhGLVotoDBa
yN8atyP9ha54HDiMvxXp87k7/WJk/9mk/Yr4LUoEDbhie4dSHcwrWoZF2uq+rmHdo99fRnCerlWo
UlrRiR8jdY0ckA9D/NxWEAR5iJYyrCoOk7ajKDQYV8qq3gSEBedaFBH3r5JPyqOpLk9Dc43xVE5/
Hz6PBwog07zP5EGxWEbArJSrV1hcxgOiwjciSmRzfTG8Hbhioju2Ww5PnyZ1AP8+hka8ARGh11k+
1I9StTq3MHmE7p1Z9QESI5bAWXmuA8L1/366ERSOoIVzEX6gJ6BUw8D8okcE6faCrhk8gLNlq6hv
Dmp4SpknwzIrBxUidum1WyG+al6lQN3VqtapKVwyRp6NLCOUVrpK8bPZbheCD9+1CpNXbWRQQMkk
rga5cGqC8NW2iNPbs4W4V5N9C5uy0HeZeGVpl8qbXp9m4j7iglXEbpAs4ULjWGLWoh5e2PWekOnR
hvFHr9HtXuThrVYC0U7b+O6rFeIQ2MJjwebVFz++k8TsAlqFwYUk2/MXDuL1bVsPcfPpC0NnklcM
swICh5f8BjKaKJN78bnXJtWES4zBopm/N/umLpq2tbXmXaMJw5sLhC1cuIyLkTGHSMKMDotfb9Dq
lYxjqvmB5ncKl+b8NVyyFAbLXKnEvTrURu4gaEu6zxKkiRRnADa1yQUgIVbS2jF8kZrJuhHEbGqR
wayxg4afyJOQlpqdYXKXxFPX42XyhrzjsrXLgNm7pz2JmCjr3gP0SGQ3ZarIPY8a3oxukGjOYHDN
FZ3KS/H4VpSdpxs1sfI/YnnCll8/tcn2H5iVVWUw1fPJOp5JEwemiB+P8AmU8ccmyTAufIYbdnfp
yUX6FbY55KKzdJOJvj2T37GleqNddpfM1fe0K3edxIUSyWh9OkFx4jlKB6BQ8zScHoahKM/lUGnr
ecuRYzyAZioPHiolSBNkqKEHKAjFEzcvZnJPyDxrTYbb0PpCI7SUpjmNITvJG+D5c5O6R5asOAGG
NNUcQkyEqeHttfTdg/ebwLI0dwE2c/hdijU/q7AUwmKhHqtwGAXannzoEdS1nHvGR3fsAudSsgVB
B5/QLB80iP3Cf/cNoYJHjq/7FuPy6nnJaVFKVZCA4VAe9GfhhLj7A3qHp+UMJDkRo0Mxtz6pQTpe
1gUtJdQch7u9PRzJgtQ6HuOoXKQPRPoTIn7anEEdm3i2VNrag+A1odxqfFT+bfgbjj4xE4mO+6oa
P2o3lSkEHifbBraT2q6S5KMYzlg5DmZdJwK7t2l1dJmybXUs4bENrrSoVw8MPu/wv9b99e9faNP8
PotH8khuM4cFYctLi23HYD25bkj4UZKBEWF33xSq1XiyBA9W/Tu2dwjbV9nZ5dV+BlOnk+E+mjXh
CCMnRoPDrU/qw70BO5nuUTeqa3z8rrr6ppsGdl+zfEMrC2JAKiqKdkxW6iCzRJT2aIp7du1qoca0
349BjEMQ3jT+zkkZMSdesDtF9PDBgWJRBFpaioI8tRl55a5eHhHuYBlQfWLCCafzgBgdFfE5ZJa4
PGA2OVWRL1Z/iWu0DkLR9brzF+zByWrl/7UAsLYmqgWNdvCyg1ZwoFh//dDV9rvDH/FR4uKb55o+
C8iVUzxQGhRXbtDXtjGc2Fzy7UstiOQnppFXcvFAzBa0X6/96XVwQKQzoFC92M+POstFz8n2qnmE
y3MflDJHGlZbA4kq4yp58BGN9f+9Th2z52IGNEWPQAs8iQ4BM09N0UsFrqgJ+K6naDwV792bjU/A
4joBJLrdb0nXo1mO2X+pf/EK+hlV6qemRVUVmJxZYmsdQVsF62FRkYuzJC4c/fa+r8b+E7/tacRf
HanLAzZuRFWCQS8JlZ5GDchNBReQOJhUD1/sbM9nyS91VtE8F7NjKd7jYvjaizeEBMMoORT/hFsn
naEPW4lKR2p6CGAAJJK+g1TcEAUmj2fjOmTJ9mD31iEguNHLdJxLbsZO2tyWU1oLRHsQjga1pmRI
IB5LPZRdClFsZP+SP4fW9rcUqnW8d2OB27lVb2a0zFH3zan2Z9CqV+Ij8kkDVs0nJX7nWuFHtH9q
sJx1OuZ+Nk2QBuNtVDcfzde625dD6bT5U1sIZ5tvGxHh1ldiLMLa6EIMDQwaYIYqQCEhurD1TNE9
jf6B9/O/eR9Ml6XoWpzaL+vX+mrbCDoutqT8fYD7Hs4NlCu+Pe6BtROJq/HIoXZQqkd/kOkDtNFl
7qoRnB9sBULCm0igE4qFIp4+i027gE7jIozLnfS9SE1nkXCqWZh74ZARen1+qNBHxdDdmPdG0HKa
zXxSXCUI33OWeSkh5aadsgSJZfisMwFHsHnkggtGiD/vNilxDhX8cz2kc1VRewDVKgzJjz2huvmQ
vBddIFrTJsDj2kRqcosozFUZY7Gc39oOpk172iaiXFXFzyQcmWKn65vX2Yz3Z6pF8+IKI/5qnMd+
sOI60rzhl1GkQNehg9CQWOtQmwfCuzs41yolCCb+uTwMe/sLb+F+RF3BdlMBLeEmHG4Hiwn2nGqR
59mNahxMP0oJrIM8rN3gbczK7BRM4pqJUqjtLGknibWZEOhvml5s/M+3gs+sW8/W87r1YnVeBEdx
AzQx9jzf5yRxQ2Z1V+nfybZbTZpK4nEQM2s1QFSNkKWWsd0MrDJw7xcihLKmNGJ1s9ZtEuIvFAAV
+3icZVArqi9dRR3p1/Mkbhaaif0CdpE4lQ1PqoJp9SOImEa7K4bes3ew5YEFBGp7tOM9bED6pNjz
4NOPvxhrL0iVUbxPBPj4HB+e6bXela/yFf57Mss5NWKScwD5pzPT5Q9JR5IG4ZzOBeDiOUj2hVPI
DSWVgolOZNcQYgeHVsMF0Ln/wTTZnTFvnfdGX2elHeOrgGhDCFGy8aF40WFqx0bEqwVEAiDEHKtQ
FGrmGBqY52tS+E8y5ihKvhoIKcjCog46xqHTJBpOBj0p2EYO/Ns9GkqqSjSSp4KAZNDUFSoi4rfg
y/+eHMTDn3BNPKLVQ9QQdi+N/T+9YkfTS0UyY26AGGaTgGBUm+obDua6y0hM/kNsk5WHphrxXjJG
bILoyDzq5WT3xTCjYXcsbAX8tzS/aN99KsLg6RWB352mNl/ZpsGNRWoqv0I/GJiTevdFKldMvTsF
wO1berLSBkXEyzDWMHDh9fZUrGmRsnt5dU8pwPKZItMdQczJJmkCizBi4LBYJgxchpBCJVKbiqJz
jGB2QtPrSqxYftE84cbNthHW/7mL+9yVVrQVbrwyq0LVnb+VyDj+ioCEzDznShlxEL+c/KxOIEcD
/RH2epVD4toN1uphnb7jULsPJZVXG1KlQVw5GcCPyEqNeT7zV/AeB5fymQk5cebSZKOmgUTF0Jfc
JS8fd0SZ713cRRgGxPRV+5UAxakDE15R17ZJ2lcmBkmMl5V1naggKptCEUkWO7v87HJRO3ZczzkF
+VXfSL3NGAopqTwOhRgGU0FoL00u1R9B8UUWFr6TD2aWaEVQputScUQwic0APZGvFJPwmhAlZ5yp
u4U+FF7IsADwRvRr9Nkjl05UOAXu98NQe9I9RZK3eAnH2nEZ26Z1SKGTWTy3vWdJAOF3bJBCySMB
fx8STTmuJo7zoZ7DemOFhejfiMcSjconCkxdIxmwwxyR/J4x5hYYG8j+LaCAOLEyB87KLEX1/vbz
y1crlhIxGWZAMrKs24D2uO1GlDO2sXTD4mjb/EMFvLytkvwiy8PamRTO8WSrEhmY7tyICWHKH+ME
syv18hLOUDBU+fVMV9yX0pQqdyq53LFnMk8jvHyXv72a2W/+5NxrHu8oTd6zxD21ECKF03Mnvz3y
Uj+04RynY/MfBEdsDlMrgelZ0LSs2lU8qL9uSgMEgKzh44otMry0t2Fjeq9pJjDhwhVn5zSE9a2F
SOfl4R8AljTTVX1JPWMv3RzMH4d8heVEQWYjWyGHsvCcjyqqedBcX0ZE5asDrbsk4cBpqtvAChEF
sexl4a7P+Hl3ARmVZkKfIs+Do0tMkhfct8isvgEdz2RGIrGiKVm9RgSTyrU6YxagFRHtH9s1avpZ
izJKVbATR9Zxx0qLY3f2mMKOSi+fCxhjSaul3vkSIcGT98CsrY6thdQYpIBXJrWIyUaT3eHzKoQH
Bm6R9X3q5JB3VfB/DhU0NePMbgbqvfAh8znieO5LUMuVip1WBNQijLraI6kZvtoexU6Vs5ygYX3w
cY9+Bthp3paTwjMqXR/ZFWNSx1MnHXhznWyzJQraNqmg7sLRn/lJqCJfSFcl+SuUx0h3FIMl6dGX
Lk13jBhIbo/aZkQT8GY4Blnc69C9CnkLJEXCFx4ieH6XMDuXtKt3i4JwTlacnzWsvycevj+owMeJ
1Ahe3ulG6D7XN5/7M+CcaZDe5wi56LtZcl1nIWYFFL+a8sBtgVw/hAOcXHgzVLVZM8Ym497GsIDi
E4tMFZTiJ0uSP10YoSiZYtHUgbigNSkxQovygHP8BQNGlwwvjeLUdD459/AERRaMndkK1g5i+9FU
pqCqafp2RmG7Cf2EyWfl4IWR43LHoSm9T2vhCg+nYnu/HvrTZRhJ662D3t32e2WluLOJWgMm49qe
pWUTCN9641RIAS879V0BFrkDbgQ4Gh6Hvmmba755UvQHQg4s3JEJwDYb6ZXZOFnALHJjDArQCPT4
/+W/dOID/twfStomuH0/NMLIfU/d4nmCBOW15SlqyDcbCfxHSkALTdkz2te6DYl1KoT0z6IHHwdQ
GQ6aSdhsCtMG2X6mwhhojdonqWq5e+kqqUbmnBksmaJBlpRKWolEDx3T32WCKIA1r3+fdtCcuY5D
vm4L4ICBD7X7K/8H3wKCETWyakHEnPK8Tzdqc9F2kTMWm4FyUVy+ibQAYler9jGHsHa3ooymTmDP
ZC7/CjFoIe7JBAERZjzzV3PbK1+By+EgXRnswFxuEl1KmA22e2ZIYijRH8fWgwaB0V+KGqyMGG8N
GmiCXTdlm1ai0XAv5Rb43s2F5y9Yzs5YTAJVz/Z+GxFOgPdvgrZEmsYrhPJfZr+VLG/R91TLOxlR
09CM9IWAym0Z+TE891gtTJSGpi5bEOsnK35w/cSkZY8QKkvc8g5UqzfKmPZ032y2AZcHUjqHa0NB
6Bkf42tt3EbwB6KipaUbm4BPLQoh+inObZsYLd/yjY+TfzOisdjqqX3Jcr2t8bAyyzyZuIbS6t1x
xZZye4HGbClNhU3a9YXFqeWANXYaJN/mLToxDif4NxblwXYisCSY46HPg5MuTZ1BeWaJWAhlQlIR
wwu+18iFKWEa48Tj/kngdxQGp+S3KYKw0h7v70XYkpQnfNDNpyzusdiPvs6Vo92Kc1mnuJMFARAf
++RmMewN6frHuL3AezZ9VDRp+qhyFCSp13E54+hI7qeK7G48r2fuqNNVqCmHPVpc2l6h/HlWNkk6
lFOY2B2xDL+5QOy2ilq3vvPGMvy30rnVBOAU+Lw6SfN3VJjXOdABAXAQjPFGZMS5hKG/5jSs95R8
qW6f9MYb3WL+AaeNr0Z3UDzq8+LCVC4EResdVJuoqgapN5YKP5omW1s2d95aO+7D66S6xUjz1HEj
VYTUDwIOhwZQL8sotRKoaXsveVpQ2MEeOWcbj1lUezblbqsAjq6pmCYQ3z9+uXD1EVT74P8dWsMT
V9yrxjU6AT0DaRa8BJ+QkVXnMueqfBKGGAjjMzzeljEcDLfl0GRsC7jWVg2iB9jkYe9mihlp4Tqq
mdl9hHeNWx7HxIqASU/iRcISCkL5l0hed1WOxcM4yXJS+Uefeye16gKM3EjPLtpDPKbgvXtFjs8M
ggxA+Vwx/iD2RHDMedadDsTnujPSsZnnSCKgfDgqSe7GChiak9a5PbjNve8rsP8bDANNqVM8xWsY
3swsLxgrrEHUNH5/6G77zdZuVxGjgq6dblDpkA2QGj4PvDhNMIQnmPgS28vTW44T6ABB0gEuMsJJ
sE4iMhwrnP3jv0AZWIFZgpGwqiFr/lXJSJmgJUwZtPoG+f+2WrjiN5BwjOja+WKc4V8u1vh6zaiz
WAlT1DfwGTvbf2UcUfUBRY7c+xcvwZ7nRF8s9IPrik7S/wvfbp7W/WVlM4PNJ5N3yNgWQgJrqmnY
y1Eb7T7BkosVwFX9n6BL39eLv2dT5uVvUbv9c+X5mEL0B7DGbpWVbjtqEJEFaYFfA/fIk2rwIz5s
mr+CJFTmUkCBJa8eiJmL+ddnFq9hzDFwGIrTOCEPmnseHRXt7BKoO/SCaEZcDXuGLekoSioGEHnP
tkItUlEzqjNoPmTr2D4aA37NuIQF/9g9QLdj1ME3hIuQ+lKVIG5Y7uSgwU90mhodMqT71Z1tkhyb
wLFRhxnZcsDIn3XdUEzQaIaB5+diuYuUHFJ7RHmlVguSXW6OcoSDWRkQA/Xp84RF+MZ4JiaW1izB
CaLEoowArbCZss1oYHUjv61YObpJ2mve2uwnMtw4kOb2m7wWqZpHO34yRwLLeF9sjDxXjUDqgDJZ
kDSn/GxeuOc+4f38lq2eAlKqvYTU5j8ysNBM6K9mmsoZBF2sJpuoeJFBCUOM+S/b5LmmEgrcBdwg
8kJ/e+HinNIxEFz9Cl8B0jwQ0Zcs7BoxT/55Rd27nMfaFzMhCbeUVXb0MKq0HjFzQVrzZfdZ6Bsr
NR0+wBMgAuYKSgAJ+944/ZebgYDCeeaIT0ThZQM12EEUKprDWGx2aY/zvz83nrGhwIYcxVzaQriv
GUPj7ns8rqsSkbO5/lMTrXEgs/FGyaigpUsvE1DS+pmY7JikG3U4LUxsDaM4t1D/1AhaFkZRlx95
qlE+T1KFcOtGxUopdhl49IwxyjCFqHkxg3zAwyid6+1Zo8TMR9OqNWFn56J48SDTg3axdHbsIYqQ
aGHA79uRTTcwopY9WDt3eLv68cKr7nPS2k4qqQlSuf4j/wCh4/bn5v+mh3dra5OA0/k8ebmzX1In
YG9OmORKaffY+PHREJ+yxkkPRUNqly0ThKu4pYFqOUf3NcTgNGqBQXeR4eLVO6zeF0uOY9MK9YRb
1gH5Py3dlD1orzJX5CnRHMlIY6MV+AGqYIbtzoWbIoZLAmvoOCTSirHxyjKqoh5Y+pyn5PGfoHUa
P6gqdWkFtIWRKeTXOKvlERQv8+y7ogB0mOGyob40iu435BgpNCNNnv4y4YCuHDTu/Gww/c+EqOia
839McXpnDSMFqaY4w1euE7UOhxJhl/PsQgLQlJHGzUiRbg5XfBSe5PYfGksWs20teSnFGcyht4em
GkR2VBFWs/ZFw9XWNQ3WBBGZNtt0+bt0HnBqPvYDJRQ2FVae5XvO9rMtwfmisXlzIiJjujeFkI7n
9ZzQ3Ef4CURoBxYMGtGU8aom4gawuR+W2OQNq637HuVZ98uGWiL25wZMBzX6HCxI3iKUWQA0CD8V
qELkA0ytVhOKA4wxEA9znyEWk7bXE7WBkTL8zY+o8StmB+tAwAxvtTOWjvTz2SOKuHFuSvo/rjkK
HTh6AIKCbtSuq8XDCZJPbVyBzR5jTqrizgHiZUPVqbv39Y6i8jPruE0IN/w4JV0osux65tk4XUJ2
Rr7V5yF0B5Ku8oR7Oq/tzkf2SK7cOKPo2GR9ePZ5TRWdneLHPBapX6RXZUGGlpo0t5300OONfcuj
Wl8ql/ZY9547QG25ma2Me4llBfOZBgs/fOcYLzWKOBt8lc+ChakhUJCYsTSnY2KxqooAFj674V/u
ccw6dBP7Fa6LrlMMiYOUWNdhO5zVrUOWzPvn0mBK+kur7ZI5Gxaxs/JsR3cM+oidsFqADaE3i8qc
gQScZKB/P0bhqdFV3f1h+URSlBXtI6/jzOger/3w8q8SiyCc/POg+JvZs39fOaoRO8rW2Z2BMOk+
XU5FOj64hUvamxmKP+TGID/bM0NxViMnYjoJqh4Xk+YiOFWDdr47EjuzIvMIGjms/F7JPrVsjXag
M0M1Zw1akbpAIwX6V/loQzaYqMjBjO5lJqUWdj04Do1F4nI7v6r6syi0OZgrOURjRsimPgag2udd
T5tS84c3dyAFjFiXAmqyUO0KYobH/MGVXlRes9vNj0CnmzBFLsT0nS09lXpVXzDpPDxTotozGegK
ISAQh9ukSea12Jm8fWPvV2KXy9TwUfVQfi7ZWgtW4GSzS82minZ+9Bvv/3C9DydKv4MVZneS2d+X
f1MxQG+zsuND8yOI1eA7UsEh+GXh8PJMRdl+UlntvOghtJZIwl/ZARr+0wI27qgs/36R2sQX6v3B
uX3RE+Q4q77KNjcqELjDXWHHVHj/kDp0P+kkONNF/3DU1GEBr3D8N8V950gOBOngnTNNN+EErAEm
gXzx/jB5IsVUF2cLaueuLsb+QY2YkPSCt8OSZTuRb3l8mwNrDRuRO5FyfoQCWB5MIcktSWIJFrMK
K3GjmzB0rINsh1/KF4sAX8n0KcpA2xE61ARo4V2d8tlOOfssljiiE/RY7XPQbQ/XS0J/ifiT17Vs
0QJ9bgXxh58TvodWZlGQZ3+fUSL3ee0DNe5dpuT1fB3DMjylXw1ha3VSyG+6OEesLgw8ZvoNwW7Y
00BMTbS2nIrZW/i7zlnT394HkHHtaQ9wQZr3o+6qgqvGNKks6RKEqtsT5lUj9rQwemlGGaLymKoa
eVWgCSQW3wTv7vVcfhWi6aqzD3K0ZqBANULAlPtSW+Jm/sji5n7baJb/5giLwCGbx46ap7SnD1KJ
OqViDxjqY+EBojQ2ohmyyxx9jBUzN7XIMZqBj1T5gbM4VjJCRL1z9wuQYSKwIv8/V4zEL2ThApSS
3DjaeDO/IX4qEzw3lY3NCl8sFeRG64kKsZNvZyO3x0QgHqOR2Let0/z+4LYkXlHwhhUl5qg0/l2w
fRCJw13a+5qxeycLG5+33ry9Ar8yuNz8ppvoksZb4Nj558KpRLie5SbxGchnVdbEqgx6rmelKn6g
wYrgPaZO/EBEe+IQfDr0gphkOp5VA3mDh04CCaA3NUB+4GgrWo2siTMATCv5uWeWlb8Ku035nUX+
raWKP/FPKEqkDxL8Cr24bYULg+Di8GdlXu3rmAP23tHNE3qvPHop7pIErF8xLZswvBB/xWPJ9z+u
6tXahTcvlSkVPxaf6Zvx9bNs3/ORxsJ65gKMivhLO+PHQq6K0hfCDaZlAb3f9hhKF5OlC3yNZZKs
Zp6evPvaFA0sOcGqX+nx0zVfOfWZnYs1KmCbo13aIqsoqyWRBk7+lpWXDxLtLPB58Y5opQsRuz+I
wlByfaKJNMBWADxGTM2Z3FWutAA+zBM4ENoIzOoLjOWIDcBdZHGzZkAeTvmbDWAoSB9/aL4YSsYH
EmIDzok0lrbYqQN6EDeS7y4E1nZaFyzHVmRg3jdOdpnLPXUeLwVpDIgu9UOMnVEGa2W/TQveru4A
ImRHxwOFSvGA2Q4oz5xEh+uRjjxO/K0wCFQaoYMBhGNmWiZiJYbaWeOdj0ouP/iSBT7knZwBDsx2
ow3jeYUJvMROp4MmKnhD6shny/BT/IMA0dWMepSPUmHzMoNY3SUcqExP3KKntXleGmU8gXU28irP
mGpRMZx809dF8TcUm0CRCNckYglGW8NVgOabHkJRRJMRUnuru31HM1XsETlWvv7ynL0jNTvKNF0i
9sG5OrjPqpJDYQrLnjt05A5ix3vXgpMD2lnfVg1ezI6jbYyJkvB0F16MW+aIIY6bp24+eZtslQ4q
RKHxMqFPwKpirdXEqFuESCG5sPKheEvJolZPV0C2fNPFzdxf2pu/JDUoNlONvcSSi7hJ6p5Jz1eF
8Z9YCNUmvSItVPukGDt/coEOORcKK5yGOAIg7+UHN+eINdv9+Wq2M+A2hrxLgNGrybzmnKrnAbm1
xCVUIVRsuEY00xFvJIWJK8wkRFrr1S9WiGtKPTYchahQq4gVcDa22ongSPV08lilx9xSYU2Y8VtK
6/tHqQv8doQLAQE6Sym4IpPRoCoNQFwzHLE79EGV+TV4wpysmBencDn32J0hlRIpwlqM+h46zLjp
5ZATUEFALYQ1KKF6QIP+phl8JpQZK+v8AttEMsdvL8Ob+b9O/lgdHztGZcj3vxTxQAoTuXc7h51Q
82z7DY2ZO8SUFT24MpE28MLLncmY+hW0l0cU8UeAWf7OyHCwBMrL240AypyOXQLlAv5Cf47+JgUJ
eX0aQUIWvwLiWiuLEnqCS87FcXs+DAtQ2KMrL+2ft26FOpIJQ62Gxexq1ZNI/PUGQH0AbqCogQTT
9pH3+wZTe1P0nXcHbNSi8dvs/oyolEKKh/3oGv0Ee9+hYUnOxhgXsPM3QpDbKKaQMJPZfvNA351p
1WNJhy9x56jCmoFS097c8ZJWIw/3oYncF1jSdWVy0mTaTATYZIwvlEJbCH0P1jIumeis3aQRuR0P
taZtyPSl4Pe4zQzBxuT362/6NndVzyWb4zcOCQBM+DTOuMw3FIN/wx/mamBdgHNZ1+A4fUcJkV9B
yfVBoasV/buMPWpw5d/Ua4mkN014NX0qspLUbvprMzoobGQlwW7qA77YvTVEMjEVUti+Nl2aK99h
j0GzlspEYI8afuQzM1aXQGvY1REYxPo1WD9QB4yo2xx1K1mzlsDHTXKQx5RIsU/E9926gduMqfw0
/g+ychp/pxUKuiBQVYqYCT1ocgsRM5hTjwTv5E4ozVfrwSj6dDk0ra6o1U4rHR5eJRHcCfFK7hLp
F7M+wqiWirehNi049RrS1gbucpJR0qHZoSF4CA9a7cHTVpOfqIJXh/6kqlomoQn3S8+y70AzB3Le
xTW7Deer5Z2rvfllQaC1VVRtA0AbQJI3VZilZNr6fLoXGcjtFgv9wdW/z6uqjN7NxEw1rlMmaEfQ
o37OG2GAG6jfY01D0trBH8kdanc/dTramv1BkdSWObjLJDtkrkotaJxWRuxn13aI+Ykhy6WAU2Yi
97vIl5sH42PeVazuJMlMKfOqq0Jz1v8to91PZhASv7rYLhwqqIS+kP1d9rQ4HY54NIQAqe4Lnz+T
WnTDGwvihdZjgipk7tEYam3pSQpg8Tt2PU8qOnRl4Rg8tByhfuvo1uj1iRuyAmfSgoa939z+EjbI
LT772NmYTHbzhBJcDP0fquUe6KGubYXknbxqfqFQIfbBB4Oi0WNmiOSPVtJktYYiXnJCuACwk3Pe
U2rBI/pduuc4KSQVBNcRiAHMy7f2CQDRYB1+iNLt2m5wD+jZm7C5xNl2myzLfMg1TiF4oRnB6cJt
SKAM0UHE9EZpv+j4MCEIKEYZL3kA75C+seNpVBQ3n454BFJVm0GU+D3IjLCMK7Aac3x4nF35DAz+
lDE5HHgw4vQnUXJaUVIzeGABuUmOxeNiu8BfZz2NxixkIdZOmgNkTRvnbQ8vS69P1nmyO7YYYzr6
pOkuWCbjz02J9wNPkl0H1Tthu5QSf5ki0TA+cbxBZ4pS939xi5l01AqZbmRApnQtc6m/htKMhi1E
aakII8MiB5UzNCCUIjbs4zmFyuDS3IFykTAR4tOKMBGCJowt9YR2EiGawzDqCTT99KTOizz5MP2z
ev2MZBaaF2LOOpzsDBGPUgru/E85Jq9Il8viD8VogYSlS3cylquJ6CCClJQPl6E4k0Qi0wzhG/nj
YZEEsU/+BF6r9FO3E67lq3lZDQX1u1l/Zaqfi6eGJzUqDbdAz1VO/ZjUEPRdOMLOzGF7Iz7B+7Fs
loIhNbbagp3VVOlHVH69OLdpV/D6ag0n+NCk5RvuP9LLwO38/HxOVB2dbi7ymjEMC7Gu9Zqf5kYs
39RiD0iaf0y+pmxV+z4d9gDnQ33huNKnQT1X/FfyqW7DXiwKy7TlpZHPH/Wr/wfwM6J56NqlpoKK
OFYGVDPKPZb6D1QKZBGUFEWXpoDDfrILi23fogy5JPRNyABYm+UV861B8sl97eL5hy9iDXlcV1a3
CfgG/pCA0qFFupk222VzQ+I09jB9xpvDEHkceifmsvpUzWS7Bi9xWuoDE8BccTL8pAS5z9EH6nfm
EYTlyEUfMVx1VAKmDs/q44ogGIWkCQS46vSM3Kh8ZBhNosUMl1q4KnZv5PnBDFlcHTreCtWYY14T
jzw3wOaWmc0B+8KNbA+ddRNzW035BV/QaP8lYdUsTB0mZymbZMsqD0QhMxpiQbYQn5KDFQ8CyZjz
RpbuAX9a/SnT2aO6jzg4BEX34ePFuvvD34r1X//5KBY+IW4oQALjfC8tSBnXaW5NMHRm7ltEgUYd
jubMX1jyq+cZZkVyyO3k7MmN6K2EYFgtJ3h3MsO1kk8TMTff0IHGGZ2EpWsMQS22T1wQCGdt1on/
asTZ1f491aBLGH3BBHV9sBpukKnFo0pGyUXmBF1sOj8V5dJLpvESvSTFTo49pj26YR3lu1z4srRK
/nXcnOgsKMEfk+6IKagQmQAOlXolZDAXM2+6HIIf82nci9ziu6Taq+rd3z3n+dKJ5zQwol77IT1B
CfzPz2/AMe5JOmbUJzbRWNvl+ia9U9VNDek9xcVI733yHpSUou8xALDYMoX2hLw98RRa9L99kvOQ
T+LDm9Q1ddCeCdfpRT4nqT4VcUKB8vhoIaIjeiId8XwhRvDd2RBLLdtz3Al0i38s9YK1dcrBFMfq
yafSqTBrDMkaSCnLVNpfdBTgP89oScJhMhTY7/fQXMbBiSJDEXTonmLZPCj+RnliVpl9e5iHVYwR
jCPCYvS7mxfyoJRGrTs/Z9XtN/Qc+g3JsSbsdXt291YSoWNKz2tT31GucjPYpAQukQ8LgZ85PVDd
RAGhxOrvM+Seev+mc5EdA3Sr7J8PC9S7h9Ra9zHz0+MUjflXphszCvde2LdZ0Dj0/+z7mGrpWmtK
CNVvbDgSXXk2zIbEeaXTDt3sccHfHuHqVm8vlUE1yKoHV+8boSk2nJ4nkkOLmUq9M/bITv9Rxt8C
q1kdmOFiveTcoauJ9ONrxX5+/eCS3F+1gOYKQeWx9TaYK5Ory5Ltn2C2v0eWBAjf8J8Qn2L4CoDc
eQQL0RZtev0ZjMoC2On1XAtM0bFNB4L/xrVEWWI+3gbeThHFiWUwQYGi760yXVon8+fT8GS3G+Nh
ot0vwqfVZikqAYd+TQMfdQXxX09BH3Q+Ez5GTktci9pzd4I1H6YlxP9ZQWr9NcXeTVivO7W/BJ7N
CeBUY+yVRexmYKdfipwH+jL4v/+ddQqRpLsuEpzuFkpeegjsLM3bpIhF0Dr9d/lG3+04AahrS3gU
ECd2D8OGrhn1M9qpt1eqsEN//2G9qCQSVctyIT7N8X0O+SPaxTs80cysVOf0mnxiOyb5d2qMdmeR
MyLXfZReUovdb4FMHGX+PAOpwF+e5pV7EtI4oW3E179oDvE6VU0Q3t8L8J8CVwPybmaspnVgPSmk
6RMFgVnsJBBoNuxxX5ZuCnXBc7V/MOdTyzY0B9ZzAxfYVXIBH18k01sEYLvrIgnSFofUskj80EcK
gTwjHcZErj4tSD13XQ3wMq7RdUSMjCjNYEYzdrQFw8FyfRD6KkEgDmrm4+kh3ym5qQyypm4Jy023
GwBifABdZmiLU1qQwH8pEXGAXUFpK1pK2GQdHmYn70DfgyHrMzkphtIehh/MFWB69MSRbF0j41Cd
FOeddeeceggKzktYZP2HHrNpjWT1oQCiT6zcQGZiz1SX2rtNjXHHyjy5wgBRu5rbkcWY6313tjew
WEf6jC835nJqntpyWmoAU9mQ5P4zwZ60r6G+BD/sCaK57LHtt2TdSoqXSkEw7MpN8P3LYX9OYp1N
TDckNr+JQdpyP6vjhGpw6Kh7R/vHTMPs1EkHQFtLO+1JXFi4VNnJeMz24tVubPE2L4SpG4ItKMj1
VRmxi6juA0C4Zbu6GWjh8vVBAHqfoGLcPuK6RX3yM847d72LnEUSmwz+frMZVeZc7fsa9FYEqOVa
c+Y+X3lLie2XLkJUx/HbOyTwwp393jWD+4WBtIjzXJBJGqIGKd/+QbVdQh7Ixmf+B9vX8W9TwvqT
+fI0DvnRpEl7Pei6HeNO4wLKWjGkk1DgYy/JU6T33bITCP7rtlazekaEyGcZ6uTbTl59dTwup/w4
pOXz3KHDoBNcOJpDd7iTcsdk4hbPvkiudyqaBIS1KklvSStKLj/5cs9NDWhgE3fUxDPHPAOEhN3j
vLcohu5RXVTBDoiIUAnQj1lbtIprJ3H1LtE7Oe0NnIoE0ZaAx/FDX535Mx402jiakST0PLlnU3T+
dIffWY0V8xufwkcotaouKerMVUxLEe5rNbXGSyziQCpsZ0XkNHP57ZwJztzf0Jn3hUzoyT+8kD/L
rH4gzwDR9Bad2+hgxhWfNpBp4R5iuBfRC6a2jDxiqAe+31qWbrc+gbGRRnmsqq2UTZSApaCVUN7a
HAjMH9yL4OG/yrFUsDbF4nfUej6ch2Qsmk7zz4THVqe5yaWZz5BuhElkBqLFCrxnTNZtIHfCegla
5kogIpb7bp3o6q13pCn9JWOV3qUDob9JaLZ7zgtmv4JYohcUkG2iqi1zRSiGMU3TKwIW12rhWqDX
MwV98bsDm/pQQO1guhgRDTJmCQi/BVAzzxiMgXMHJCMPM7B2T3u6lW3fmDT1ziCnPv6huC0P7mKq
5StH3DOQfaAiDa5/uQsXCzvB2UNG7LEsi10BcTDZ4J+5Ev5f+/kDqQi4NHP/me9k9CU49u0Wu4a5
zBCXM4hQcubAz20Pe0IhkvSyOfoMwdDpzplqoQYg7kSthfFDOb2mDO9CAx4xs3JkfOQqdhLfN9sn
5HnYcpFrRVUCV9RkkWrn0J4ZaLuGd5MXxWmnihOeBRGhzyu00NwwEWdHSbraeBOzlkoXjb6vm6en
4XYDE2OuWdKTw4ba5NuAmO77sX5zCksJ9jnOkFIqkiFlwKQGhaxz2xcJ5+tfOmasEi3/RV2uDFTq
ycBYG7FITT52LwLAPUl+saG1Pa0ZUaWGQkBYZ6J+Zu+oeJzyh1RRxohHOQqtP/U/VSp/W2hYIzLL
+C1z8ZXpa8uQNQyu6A3ZaedA3MqkABuXfb6K1WytuO+rSaW+keUcacWDJIzWry/ISfI4/gQcylQm
F9Og0PfPkId6wNBpHQpjLJM2Qc7vVm6FjVqq1ZaBTw/0Z9rwVjBZutBjixjkFOK3uBnJcAxDXqOm
ioFoBDlxVYdkQR8AfIZi7uboO5zR4AZBtS04j1xYQAsUr2r8Uvm/yoIxrL1K2LRkyj7O6f8dToJ+
J+rQnVxfpGw+zSOvrkLJU88l2P+bJ97Ipvd+Kkaq4WbSyiXyc5ZhaxFbsf1WQcNGPIU1Z2HHrNAC
xixtgsKxA8MJXOSHsjxTzcsnw0qwwjEytz3YH7QdwApz5J5vxrpXdh+x4NO9oaDouVYCw6KB7lwt
7n4LlJ2tlJypdWgR/C1mbZEuIb3zVWhAPXkY+GHh7cJ+Uoj1ogL8TI9yqMgI2JzWN8S3Yf0sCxzP
1OOT/8R+vWsjWVA514CCIisbEzilA888XflTF0ew351jPqjxQIsYJpbPsqX18wAqSOeXchc+Gozm
+4+ZkF4ulDXNoQxMpAGUVHe1HSuV0fjkaOXJUwG0tUbkCRhSa1m+TOJKCI58fD3pNe+0f1r/9Rjm
8Cq0qwkY4Vd61iAO3mpOeIY1w18J8jJgMUYi58aSkFJTUaNbvWS+XKq7eUncTaPAUAcOq/ADsV/r
C6bSN6PGFt96V1fHOZSaTtM9/3jqKavK4XpFdXy4SN0udBzCkoMtz/StS5kZAOAQ7buNPJDxfV41
brpG7cGpNHMBgFekH7sO7B52OKctH+t0vbBFg7bvJYmj9ACUDdXWlYyq6miuB7l3Hu3eVwec75N4
CmCeOKSf8Lxujtd2ClR2E1JLEVDu936pm/IXF4Tv1/2qngkdNeLirBrRwizYJj2xt76t8i3FXSyn
JN6BFTug/QxUvQP15zTd5W8xVc4/KNEfkoSaodtuFl+mx7V5P73xm+hvjp1/eTEyQqzzDcrin1Rp
gWyIJBlDpYups2PeE+Mi9BsP54QbM565/9A26YW/W5V36LL81e/m+UCbdWeRpZP4xUV79SinrYBz
vG6L0FfjSU8++HMw3cTM1Pd+z4qphv28XuD018ZZ1n8eDKkpJFrr5ynvy0cX+RZa/TkZO99ynhwA
+WyBUiideduFGfOr+Ee+QCZH1/Ni2hJYVCQwWzq+5emqYRPInrXMui/GpJPkmYZSAuiGbxlwNEn0
EQNaIYfULNKlCzuKIOIMRRSKDRTKglkuSltRRJJ++g0FtThaEg7ii/DV7mDJq/PfipL3LpYIJHqU
mXvd48+4Mrz8jA7QEJAOflQW1Nf5cud0zpKLsA6cn/j9H275JduljUc9loxJnUmamInwvRyZ0rFs
twNEqyaA4Q9zKxo7ng4/BrnomjsQvs5gRAwSvKsIJMN59BGJSDAdBSDAd9MbWEZhqhoSjTcmX+Y+
4qZ3x+k6lM2/TGD1r1Dr+e3N8gRZiRqt3U7FpnKGmVeqSAvmzsNIlLZuQoWsiS+ihYNSsDyCRG/O
ZpyjwGeL8Rp8CSkmEZxhL09kNiZlMmz7kwKIFnfp6cU2ruRjEUTlYtiH84GuX6zi1XnmNE+coynW
2BVu2YCF5tiNaBz8g89/0/sxy3+13yREzuSEoUaGpOEYayuvtX/NrFOISGcn952Oa4R9AnQ1AUI4
78+vhUS3vr44j/oGAJxYPAchp2NEFevcutQYcEZrZtqUr7QE0T61mG0h1rPOtNLdWrjeX7d/wJur
jCKC5Kf6wLSMbjsrBxWNF04a+9P737rzvHdydbqRJcY7Jzu4asTTQqief7HIgh5umb9FMbYsRCw7
QK8WCPPK9yPC4co7dhZiY3A5KhDef1HnyM0jG/UQa0NWpII7mK7EwZQvTPC4ATjyf8MwQ9X6u1Bl
MV6iMwxaflPMQiPGr7sn0VtA3QkPnWJIxuacokO34u3R6KnTNSZcAiC6qH9Igu/aOd68eghPTISz
snSJRpquzsOJnvBU7TdxmorBkZ8PedIw0Vwu3ZqP7bU5z15auWtBII9mIJo/w6LBGl+UogYSad3/
e1T1ay5bKxBAsJcJRNdh2cwMW5BopOpicEHIPWSEZxlW8GTJ43L1r8jXf9zmDE4IJAUYd+j1OjOC
q1vy7UZlDZ4J7aaqTo+UjfXdDk0RKGiL9M+zJU/fXDF+94GME2lBCEyHzUV45mviELO2a2WQwmZm
qRShKOUwQ7mBgMgv70kIaya9viRXM1mf7l5LgaaV2TqwZOl78jmtt7t9++7PptGOgV//dYqzFL4r
uQawcalb/G3JA4rgi8rYRWFFFflha+GBGRqHUh3q220n1dTxnZ8HUKOx2wn6HnxvE4dYEikW4WCv
zE3/tcSLddm2IbJjNLNB/5i+Tp1y08wlaN5+CRM2CYhQfeCw6A0MbYOdaoeRMNdFpM3YGzLL0UOl
pRECLCGHeZpW/wlWyb9IRl9++1Nd+LQDhkLcO1t+iumMk1taCeSTsFdjP2B5KY+qrrCoPtlyPtV2
Po5ByhiquktF6aZq3thy1tKPk2Czxii8KRjNaGdF3rCrWfjCAtVRrIfZN2DAbzJeRxfnnY4mao6w
9YU+IEGBdBCax14bgHQIOFtYGVR//j5aPWAFLf+p3/zvH8jEjBU2wQJqPUy1YGCFSqfkbCYBCy1T
yQh0ZcS1bFlndkOj5INTrq8Fb1zFUL29QupNLxAZ9g6J976JLF91B7ThY9+ZRpGqXUUTUS+yCJAj
yRrIVbma83J8XDOwOe7kniGchFcxB0hVS7idDfOpjumxRsno3xzpBO0o03zm00WcmZfwcBp3f/c/
O9QOkc3I6sKbaNrW+NrrVmKvumh3d5vDdOpgt5f1KxfSnsl5YqGPrkvQWZdcU0wCSUu/8cfp0udd
vhhnoXMm4Y+75huNjQP1rn9YtJPGHuLp3YoxM+nxceoMFuvZNnqYkpoFwjrVnnW5QRdAZO78ScYl
X8xoRKkoDDsLk2vHZiRDqdLMEzt2v+o2EYnsu7I+Sn6wINB91wJhEBvC/ebWxQh4pU9Y1CrXtmys
busp3maI351woAH7+AThZygE1PV38vjyEIjLJ2rcsdoLbd/iJ2qFzz1DpWGdI8H2PW3QZxBpyPFz
OOU6v0vQM85rbIB4TAuKru7vYwFtEpsaGbbPiO4V90q7Az6R2K8nkSoum+CE+M+ZtLUIT7tn2yDn
OvgiPqG4/rYCTgdahwJMAfEXaXiGM/gge/pb5M4WRO3P/GvwKpZpqsI5dk5PwEXjn8YiTPLUzUXK
jsyHHyoo+T7OHL7aJ82gGV7sGqRezUgieMLnfHzsyfgFm63QpKTZCQEbi89hILc2KEvKLN/w/jkz
rKB8VSPv22UipEDzxsDK0rYGDBPWGzrjFqAVaoxH4oYLm4/pVKnYyPLtpfblXpQiP8MrVd+1s75u
NvBAuESLbBKPWf8alldpoZvu/K+GgUaK/o+yS+ryu/m0atzoEI/DzknvwVlTRBcexSFVmzo+81y+
JpXs7WZ6H0Rk4Mhjo7H/wPYnO3m1m81m6AfujLP1jJNPg+ua/GkWA7M5rOuh9WnPZ005Q5zaFKvB
W43arOI73JVYgkTlSd8hE3Gr4bHTuQSGvXLDS6PvYlUify0+AA+oyT/3fkgWcav1Z8t6SAAwJMsL
PrOgbJCRuZo87yIForO4CMB/NhTMp248GiSIiSSIBRV8ue9FfPoNz+MfbDpcgU3/3HRrRA5pm0no
qBQabofEfvFm8LWA2VIgCLeGHVH/ibh9aV+wlbaeAsDogKVQuNqMpC4vmYVyMZZdB5yN0UcmE9rV
Qdkeip46l/CVsG9ewKI3sn2Bf2vatikpTphglgf8hlXaRXBmZuFyIFiWeC3C3coAj8eyYNDv7zxl
qb9J/3V6pyKHJB2ub38Zucn0E5fkKyoREC0HQsIhQTi32J5YZCvHnHXBIlgkIc3Dr1uUafYM7Y6J
XAOVN0FvFrKAp/GczZ+SZUIb+qJqZ6SPQZ3de/X2KEzu3hK4evP2VCnKlN168QZl+73pQn1nL8Vp
4BdGX0uYY7I5r6hRIwwQzMPUnGG/dyaFvwkO4m5x/3dR/oVT9pI2Z1TXcXnOC8Adp0SLBWpemlAK
ru29YW4+ZM0hWBXRzotBNRpEZsbSJFB+E2iITPmPSEeHq4mBP1ka4n0WntimbLrAce7hvMmKD9cI
46j72C4yPOf0E2h/vA85KzMH4Hlhpdgvi/2t3ELebztsqVv5GOecHG4aqBEddUbIu5+GwLEGN7Fx
hTlgaK0IFEL5jhur+xbHq5JDUM3ja1tm7VXpPg6dH1g1N0/0UBMkhr1wYYaIrbk/f5pxFqBCwZZC
KdLS4kWCQZXf1+eXxu36Rb90qUF5J7Z5HDkwEL1nw+7oGqrzzr5rcy8qb35uNDh0OaFbv/w5iPhl
JKL9RC/dtFB5b1jI6yeaboFqnCHXSdai0oiDTSSgajcf+WNJ4OGB1XvIVAhqqKSxqqZO5Pmv+Pyd
yQSoebf1CAEDas9jhhgL2mruzIB8+wRy5rbJmCK6JRdqFmhplO5SYrt/gqbayqF04FzI+2gTF9hg
pXE/6kW9MEHGUrC3hjBcveXf6S+V4ZpUiZP2favcEZOAwxHraJIR9dUgCu8FgxiQ4rgx/P+TtZVn
4VRHJ7krgMJb+vyHuXdSdkMM0TY19JMr/nRHIkRB9yB7Igc0Q9xSP0dHvToEVS9eH4MHtbXLXQjN
ywSaMcebjPLbrNqWbjfZMrUUL7LbzoeTpB+xcK0AmhxsKXqXk8kjKuILJxztpG8RSUHHxJJWJVGZ
juVO0UJVtm+XToNuLhz9Deu1HAEIV18jNy4s1OjxxmpzPfkfMdtZ200MIY0XYs/2Y2D/5sDIqjXW
Yc4SiHQWULxdhqgMKmJfluugfsfge0SO+aJmq2ZGcYkXWUBlASiDxdvwHNOJv87RtLdWdPOlCbEc
gM3HaPo4uhiOoIgforpgH6RHLGKW398rsCJwBmtnMBc0zvtIpHVx9x50Uy3rze0w/7QeVdhMWPbI
e0RiOdg3ZYXow4RlLmJTd7z6pCcQlJJ9p1l937ka/6khAr8W5SM5CtrdklwaMs1ffgA6QgRLw2P+
YLWu/kEAPV2YWaZyJCvXkRMjzw3f2/BozE8w4t8l8o2JAaS96MyU5XEzdpQpEVOpzmz4qTFdVOHD
EhmTG50MHhZ/5gCuTja8z+WhyzRxNd0HZj6T8ofHf3eb+4YTGQkNKAxS6YSie5cZlLXilEgUnqmI
xDijz4SuyblIP3ndpRrx8M1DM8yX0Ld1Ve2RFJiFWT/H4jXxK/3J8crVOKEkye4zx9MRJuGbY/1U
KWsQstKlksgn7ZqmvMdhnYV5aTQ8p8szjjh2y6t5IMC7cEr+x0G6qLJf0GvOe3/LSHDwtyliOEpB
VDGAt0UHc37TPxNxQhbc7eKDmR5SbQ/uTl5PhysuHt6lPtZHMsN2ag5iap94a68GWPaR7GI7X3tA
frfHyuJEuAzX/gPg+4Tj4hqc23EqpRjnfh95aIGxu/MRKb4DgTapvFJ7CPjiWQwToP1RuZMCNSuT
5GAqLSJBMhF0t92t5sE04oMHaFBaSQoNy3TN3xdcoKu1NybtD9GjhcZNt0xkUsyoX1XZaRxNEW+9
/HCxSyKlDV2P3XC6UvYIDUJASSeO3y0LWzilOBpB20qzQyin1k0Fk65KB+gc1aCNrSxgvDAETDql
gfIvYUFkBfmEa6kexZOTtLfqiiX1vTk5NGGvjTuKIOlp9L7eyjojFAX7zcrdDo/3ulYAci7LmdzU
MYyDxy9slOs5Au8Q3CN3DsDS92fgKxhawP2XZE5PRjFyGrwf841kQojVN4jMKfUKfAeAnrmVkTzM
rOHoBs/9Q2oYft0BOiBaoI0XnmopOvLCN3X5zJm3++mROPr0bWQMsl4sqCbFP3yHwhWirR74293D
E1UESXaWBAkhxjFTFEkF17qVt0qZecQc4MwT883DlXjt+BBdEUYZharqSuuXPhJ8Ibw08ceLZ9Tg
PMnofCWfSEzUDVxXXCgs0hPlhSXKrZKHHFGN3A6CbTnZ73WYSNIbcR1Wy+iDTgbzBdkZLAiYmTqF
8XrlMx5KAv2PhTP/in8NchxoQmZfg1STqAuz+pP4tHHc2FlyDsxnswQDm8IIABTpKg6s5NsTTwht
4IYAMga7VH/uBHZ+D5wvSlK/PwNPAFoW+ThqKg/XcAZ7W1LX9wCMQSKDN+hy81B6TqvLIAeMA+Yl
StHIrK2Q619Qlu0XaqHE4xl1Mn+y2GJp7hNDyJAGCBUHz0OxS9q88+QWdh4tZJgNIhtkfv1t/Trp
fLVA699a4oTd9PUkuZbUI+mWbKDu0At527pauMBcNzrzrQhmmjORn5YDIWtcUsnW0ZsS07tZHMti
K2nkApEin+z9vLaJ1a+8gWnqbrXeeDgIDIWqF3qkepNo6WXnCv22a1Vf9PHckAenJZALRRcImRgq
aHsSw59YmTFv6uMTHTHPaNGPxDGKLIAeusngFKU27ezsRQbWxCL7J8r2BDPXowZ8ncj2Pp8wplLx
gX7PO/GEIt65eM3RXmUUssts0e16d4STjlfLY6UHmodpLqtszbv1cGNMT1lDMPcPoO9HTcQafqbr
iOoNf7Y02pmXyhJYgW891UtxfS4KiullQabEO1YxRUToVjTCQFLvEFpezfMEKmVYFY5vswXhx0ZW
K/uToiofOPcNehTdbeyE4oh0wrm7Arn8yhqR04g5Pfb3qWbfD2cq6q2i06UlXLWY37P/hVsH8Jfk
gSiMM2gdVgt99hsm7i1dfXl9zNVmCHdOqVgXxGAJ0Kw7wSRKDpdmMNkwQOmBYJquhecZht6x75TF
EdGJRjcE38oE6X1iFsSBNPeClMvnedJ2QQGlX+fHn0aLV0iMEIVu5f0P8pJa1GbeUCmtDxYMVXO7
KYH5QgmuZWV6HZbnax6sJL3l+8Ff78kUxpWgizbfnnNiP6y99druQF9tCHpRpvIMPdF4QJ3CYAcA
ThXsGgx2OJilJKQhBH9zjX7BRKEG0Rr0JhZgLkJVQnf1jNv0qqFtVOjrEE/E7v2gDhBw6gxBogMG
akAvuzsDgSaNB39l3GtQHm40z63Asi/WELmHcuB5mdEyLSWmBUk9M+1HvXTh0sNdQn9r1O7wBzIJ
xxk1hwZd61Erkas0qSU7xfELb8UcWOTDYLDQS0tYfT9qB4QhWKDEirX2muceQ43HblVvyLeBTfYL
K+85VaCKRB2JL8jYted++65gclLdEPbXdmmVt41+SH7tTvyDq0EtVqjGKRdJLsLm8+x3XeXO7ag6
YwopebLBVib14dgKJZs2lgmbqJUldvJkAr68VCb060KUC+cBLVsHOf9dV7PBwmw4RfKxsY6m89XK
heu055N31llbowhfxqVEDxXP6FdlotCiUlqZBU3eFMttcSweJOblHIFlStXiiYmLHE3rU5a/fI+F
W40aokfYDUuHPa1liFBAGvEZf/oRKe4ZPQwrU3NdnE4AVxqK7Yq4SoWPsWoY8DTGQevUWkJMkmDF
hjrEpvswDvB7laxoYJyqjQW0qQ2iaBtl1uI3jpVf4N7V5funQD+o71vZfBVkbb+EX/FqEnLp3rUM
L9C5NsXh0dwgAjNRNqBmg/KYVk6a4Z7KSrg4OjLulyV7lH92AU21lhxc3HzLUIhlALmowZAEMJCk
yxkD/NWhRx34lexWr42Qxvt0nU1LWK6geTOQIIT6DHxlgullAl3NlG9ahjGqSMtecrWEp1aR1i22
CF+mA1NJdEKLPR9Pa7i09kEQrjtiKobCbkHNLvr35abORsIghXd+NqHjbLlQKw3EFtxYa5fUeryl
Wi+n8WHGe9kt9yojAR9kurzFcK/b2VJfN4LZCcMV3KEy1vgLXb/kwu4x/ZNlktVNCiHmg6Dxy37e
G17tzdx6dL87yWuYLsCVBqdxAUnWZuy/3qPRMJHfFYGvR8hQ9qFwMUPFRGvFC0xg9WdSBbo5yPUw
bDpk/jXfNRuq2aozFa6GncRO9vo/0XhM2DcphmxfC3jzSroMWe2J+hZ158mAmU7Vs82SwxaPPU0O
6cbAdz7EIAptyNGlwXH98Ig48YAJ9R4gzaHx3mwGZwSSDb6yf+jfju+O90V/cs/d+lr/hK+lTCvm
JFW+gjXt6rG0ChoXs1DwN1SYMY9GDyg/TLXaQxBHBm1nVBD3LOaMazrhAbRM1L/wGDGlqVfmDI0J
SoLBMrnmKGqM0XQrYgT1/XrNc7Cn2g7pALISXmMHPGz8NZYHF75/NUQPC5QlqZWiENkPZHdiBGhS
VOhnZpe0xnpHtvCFIuv5tc01JPJLu0Gd1wLVIYp0nv8aJkiMbX2MHPGZ8f5GfdQzEVQnpuzR+5zK
mODZBRCkEW9EBq0xRPPx15Uv1KIDGCCarScdJw+OYO0b4AsfrWeq52DpP7qhvB0tSVB7QL/9x7jm
87FaFLK4i0U4qnaTf5pjWNKbdjT0dhF4yXwFekRIf7fgogBCRQhkC0fprJEZvwH3T96R+aC6gSPO
EFmq1657fgn48WIc4p99glLAwBWxFkrA+9tJ0QSQo7MVUFq/cAHgTCFkR0w0TQN6+5IAYffE6M0/
gwFaOrdRxmSG4mt/htD27fsV+aIaj1VN0KuWEVlzX+UGkY1vEzUmlZ9S7q136ZuT+T1KcSd2ew9q
wT0VB3Ng4qiL5sUyfZu2sWIy+18YUo54qF1mYxs0i9g99sz11gUWjDzEqLFRH5s5fmuHNxSrpipw
yue8iw8XV3Yvi0zEogeoMW3BQVd3fOeDiVfTAWI1WUJATHi5xvz7K6GaZFrbLV0lkfWJtAN8eXZg
d4lWsnZXC4Zes15gsoTHfyU9X9xALcnvyEL7HIthC/8+fCzHjgf7CLapt1c0TrWzbqCDhi02KRqF
56kHhf/5nEHASsNOuH3og06ovmuwkO4qcafv+5Cq9u711lXJFD979Ky28y/gXlCxvmqN6s31/e9h
dJj/N2ZW8f2LD0zf2/tMXCMduQYxYPTgB6XFa6fcYhlOXNYNeycK0sjMBf7OfASORShnhl773B5c
KjPkpXBAnTAPdUP+WIgCfjZNBG/YhQY4e4s38E6uiDVUFLJV/mTrU98tp0wxtPiTneAn4DYMP1Fo
zgqZrQYV3BEf7Ql5FwtPS2uqkD5u/iSJhfNvbZaqrYkCmXbNPdZNuA5AVWqa+sZpJPxJMejPGq9v
IoVdS70Weo4osfWUrqzOLaM4xuIOgnaRT4B74gMXV+O1sVaZVaiKsJaBq9laWEFgy6VRWV5wK+a7
BtBEoxXzvzgeroUEYWkDbocAgRIMBhpm33UgFk16hJKv/eqsk0KzTKeyByK6K6j74gdqDvMbjtR9
TCd+1utgFFHJSsxwysdRAxU45xyfvFiQmDzAHms032UT+T0hQEdTKPGVkq66+JICKEhwrhEqIP4W
w2xkD9qv2tb5bT7jenJBG9b5+W4SjJ41XRG7FCLk9uZ9dUCOTGqpOCnYtbhW9QImUu1BrHrqm/ug
W2k1nQf9tJirnK+ugDopJUYAO3ucPfjOJYhpOX6gQ1IGSi+GhfdYg7qi8kTpG+3S/2hFjT4XgoC6
20ne1Bntzstp6y8VoYUyTalWTZ9anD+2Rymi0HM9njRZfqOHRlfiAzQyJCkGXoW0XIZR6XiEmivu
HfB/9Qv6s8vB2PC+txgrxDLQKQjuVT0OiTdePHyauYzqLh9L3dzZ6IqyeZQS1FN9W5jfECjBvKBi
/h09+ei3TjOo215F6U4aHGUsHVwa5ipmcPtdwiDOQeOqiJD6MXLurbBpKVSxceRESXRtfLAm+uXU
u0L89ozMhZnaPljAPKovez4EcHGbmmws9K06iphJ0Ls+omJEYCmIUv/oz3AUtI03SOzfcSwOcc16
Xp9aqItP1uoUUK7LR5+3OlxtEnXLAZ2k7k5j89aQX8RpZL9/EUGiKOOsfdwclC6hStErFlXCcIIx
5Kn8mS+J31ZKDoEDQnJeqnaJ/khNi1NtBvoG0Z9qij/Fr94zOOLwA47qB4Xkfw3/7cGbR/DTi9wO
B8F2Maba/rAJaqrOZ/p+Coi/BzOzY8vUZVNwnD7DKBVXXkURbyji15UrMatHqLLCHIu3t2GLYf74
ghCL4dGfvVkzzKS6/ZAROELhXXtmeB7klkEk6xFVnBSargjts2h8Qdh+LndR5bn/23/Pwc9s1U/M
J3/Vm8DtW84IKHz7a3whPV46ULgy8PQeM0c6i83e338Py0tNUBRkIwnqTmjVCLnSzOYLHxBXPMkf
KadBxlpi2Jd0b8lX5F/YQIjXlvKhKRTLPKwGiPDVHH+kncZ2n1lvu7ZuGt4/lEm/ZKv732rJz/Ul
5xArlLG/ECcpJ2F/zLA79DywvEvqpfL8koMHCiJ8YEgWGRgnHTX+d4EK4CNNWOmUeGWDFYNEc2Kd
k/PGXojlDonTQnza6wdKCM0cGQw0P8W/nXXrExRQjZm/Ei7rfJmoaCSgwi5uytstQvHyuxPpf7hQ
8JMGQ3DuC5nVYtQuHJ/pW8OS7Yjd+L1uJpjHAN95OmN9HCo8PTez2tA56Y+dY8G8QjLRKme8mYqO
EBBNE9ZvaBhbllO9hys5zxuj0McYklGIlzTlpW337Z1Z/2ccFXn2rVDee47zTjbUGFLmQq2uh0Ae
m91DUOS9yhVkNYj+qKqA5Jma/U7QPNPNuFDqTq8Gs2OFBfWdUII/C8wIdQNmKHOIcxdzZ2gHoti4
ZgXW6R9CEnVUJt+ient72nZ8vRUOiC8mzlMr3nl2nZajodpr+jzKsLU3L9kzGTgt53o4zm5jq+R9
z/01/MFpeK2ziwer8NA8Dn5oRiyARWaiSTYabGTGcIkhX8AJPs8clzNQz5efresdeS2J2SlZPb+5
SnVNT8SP9Eu6sDnreWDSTWUOdQRN60KkIjsLc1cwPmgHHC83O9EduRZaEtvzWtTbsUEqaKy0vMVO
+Xk7V+xQI4wbRXkVskrHFjuPZ82i7wJDejSWSFtUy7uZm4xaqtalHDvBfoxUP2DyuyWThS7l7kzN
/53GvJ9ktikId4f9T0qBOiQ6lL8nyRo3xJkZQVzQpyjzk/I3wsz4xz2+HF2o/0dGJGkbOKv9i0uy
Bj+1iq36DzyZyyqZ3acPhpKeLzzqjLKNfbP2f71gIgsfgujwp8sM7ZVNN20TabgqA/vPNZJA29W3
83vcxJ/sQwscefPsWaqV7gs95hGOqkfVGbwc2lNIweR9V43l8KIWtxH7MoMf77eKB7K5ppt2x+1/
Qa4ZVjY0lSHGBq40O4pVS2oDdv/2IHxyXU/iYEqbHPH9MtUdBQ3+VYNKbNq5ztEPfMitBM3IW6L6
u51sJLEbMdJ3p34VITrkRMG7+95jYo5eGgPWeHuMAx00PV86714H4ahEQAZO8WdVzxZ+85c3o/Aa
xDcCjTiYm8Yo3cHQch+qtzWjMPCOzHmWkTfb3TzLDjiI0eTbPiYbl6G/GMQucUzXUBIb37QPwfUB
oKYNeB75AXV3bPA5gWXjn9dtcNSTS8liNbf4JNozzOlr5ITZTC4C5EamDHDeMS1zSQ9o9L31XSSP
4nv12yoo0ILGlZAr6o6u7Ue8a+MbrF1eMHXj/Q+wNpdKPRn9omweJrjkw5Vv8DJj76U3F91sxuDu
Kg4/KFe5nlPojdF+Ue4zdmr47L2iqjTq/I/bTAIMZs0uCB4TuJ8IJkK7M/AU9m/HcMtLPmJZh/Li
5l1PpvYMf9dEZqWy431SdRqeOFSBeHzwhyZnEstXknut2upFyFySQodGnAC4Wh7ui80iR2/sVmI6
rSrVzYCOaVu8Az6c5veuihLMQ0+7GZLopZaRTmuFPvjpS8M4eUveTI3Wt8AuOKFJ7H4In0BNgSSZ
C8dnkuFxWpv8bvuTOnVkqPSkk8kpJ9oFTTjlM2W4+l2GMnPvuA3q0BxP9t7vL9fzg630gaCe4IF9
UWnZ1xpVbOhHcLDQVwlOop6PHOh8oLdwkLgX2kmSnTvIDZEAurzQG7F6lAGVNXWabqerpxy0OuMO
8V23FtKsumnVnkDIs9BbC9BmJi0xUuSzwUHEu1I23zKm1ywYRaJf0NGDhHx/Pw2EyO2jR8ZqsfwI
cVP+hOsXSLa+rfRH8reOtZtrC0K1FqmHY+tW0kdlVrNoAD5V284ma9kmbZD6WO8cc3ufaciljdkX
CwMXjL3hillWAZF0peSwzBSsawi16XSZxJona4EPr81V5KwSHXImZ98db1avQrUb5EVRRMF7VR0A
mr8aiOzSaYHu3+QCM1Cor9xMhvxS1l7rnifuh7N/f5vKUhn8DOBr+ZlX0bIpf4WMepfQdjMoUMEF
HLqspn2R12BpaT7AZ73TAlDBMBwirwodSvUVOo9+qtdxIXhJ/YC12H/hEq1Bttn1arvq6JM6j3NU
C5HOftfw/O0JuzmLT/xtkw8HjtLlrqawxqH7BLvYBV3XK0dJKG8WO2EKkMnPGMFqhlBDuC+P1Vyk
7DlQ3Ax6mDlf0fJlGxSxmjpNaQcSPT2GMEtmlMhuIpqklpbEdIohgUFw0rUHMIIKz25U+ePq4RER
m3d8OKXL28BdX/8EHPh75WMwb72wbN46UlORg7MSDbho7gm+BJTaQOzbHw272gKYvIYAeXHffI5u
GD7w3XnFjQPS7jbZjEvNjViYsd4DVlGyIFEJMSPadbUagRqyLMcehCnxvjUx0L2OMrbNxwEk9X05
IyMYYWq8EV63ebCcjK9aaPGz1lw12G5cURcD87tfl4uf5zt6jI0UVGCui6X9t8129GG3b1noGZ91
XpZdlgUbGRqR7uaToQ+1O+W9fw9FwEesCLCXi/cgRPUhpHlrMRd1LSa5sgWyrEQqVwdmJvZmRcVT
lNTGDMAk9FcSGQZBClCr6qM9Qb98ID+paBgGd3WYl4S9PPwhHvCgIIleWC5/fo/+0aYDXbi/e+y9
pw32dQcRBFG/LJEkB1LHcXRAfS2wEIxOIgyEOSoZHYcNHcKHvl97eQYAdYAScHMPCPnhbHJmUDes
aH7NW4MNCZ+YxvkUVTowBJr+m+MSfI1q3HpbeeIqZuas7ytHsz7XDFirXdq8BH0rrNfI3nOmDoYh
3lLkPWatPQcvU0KuLz1mh/4CwBwCux9/4g7emPPgLRYCCUXpapQOabgvH/UI+aRYlSY4wXq4p9ss
kwl7sopCafweE8kZutuBmwGSmx8WiD97W8DzsEZwECkkdfK99lupwwDrplbeMJ/XVpsasj2WTfdt
MZjR75sSY7TYxOsiyAMU/FqO2vGAGEYMPldHw0eam+pbQwRutRDhxBUk6Ptol/NK/irfCdB+CZTz
BttYlnQ5Ms4NRsatGeKCB+oVIWqFR1PzDC49D4kPiODOle3oD1/KTPwxdxE1dRBMDw5CAXb585qX
FgDaLZl83nb8xQ86xdXZ9qwgSYJBE08a5AEwPxHWsgXAL6j4luEDL7WR/1A3ps+3bvxrAoIUGN2f
0mXWwGMcG0vy3EG26RFjJRazCNRWlKJPSLQTO7F6i2UHdZddvYzHKB5tRxHhkMpkt0KrH2w5o0r4
kA2uT4SOVNZhiylRZWWkTBzZZC10jRJSEfW0WfI/v6jsEnmkxKr48h9EzkPQ9Ciz+EQwOi/b7LFk
r5GGlaLxJf26EtOA6yYGQuObMkX+JPp0+wT7ez/pbZwvIDmqYtv/QeJ8ajahODjCs5QunXaeznSQ
q43Trgs0Ylg8iNqLORGm7CpK8p8ZrEzt9TsQLxrrenAwIUhz5Dst9zCLcaTi4CYvP0q9aT5wKJuc
VV+b1Vh71Ak7TMdlsX7/tD478r9Mt7xg3hP6axkUqn9kVqge3LEuV7R+qhcu3nJM34G1VyQEtQSq
vWo4u14Abm9e5MlxfHafFbOJgrBExsrexXTdRrsd7Qe79tScoINB/ZDShMxS7kFv2JKEUKUY9bR6
i5IUD33xgwOh595SZzmpOvxJBXoQ9MHcryIOrsCZ0BWInVgWV/c9E/9VrvpOfPX6B7cezJv04S8c
hH0JzawnJwNi56iiI0wgSQvfSp+2utu9oGNi9BFb7fumaGlyppjOC927xc/PNmxLDLTAly0ZW4mE
huRxcqiyTaF/oTULtkadlxJpuUHfSlhwfl3HdQSJNvz0QWKspZRZ6PNfPBXCkut3zsRbDXUtfVwZ
xHCZbtXZqcPj0BgIf3Ft9l845EVqElqdgLUWsDqRU62YMJpSZeBMXIIZTAnfYVsQJQZm+DTxwx1i
q2SZTu+wIXwsLGcPcJzmw2wbo5ZzacjZprkYg4eGUujlArhNC/rUXSAtxBYa2bie39rEXWv4/cni
V/uaZDWdQ6J/Q5Ll21fzF+An6FrZ4LSndjKU5vuzKxm7qvXP5qxBfieI13DXPejJ9Ns7v8iAdkMf
/eTRrKREhSb22brsnZtcxKQUBBLCZSikYkm/6QOjtj5hZo3diVeqZX5thCELWIujL1AXlREGdgK1
sq5DO+/pv+GDccYL9UnT6OwsLRnTdZrOJwX9b0hdkJlbtvNHHV7PBuDB+bDb83oKx8ZtcUfZwNnQ
QLfsQ+g1dJutmfJdb75LJTBSl5U5Kf/LiII0xWeL3a3+71utVXFTpjWJ4TDE+9HbZlE1V5mayR9c
/933m3mArTbTIjcTBM+/fAee3tckoKAue4VbmMQFrirqTAPx61O12GLYSLRJxZjzvIWeD0xkctQ8
smiYLX1B9lpY0gqwgYnU+ApKcRjoUU4RHQXnp6lUAaPjkJawYpc5h8R7hkdGmNudz/SyjNFm9H9e
08o0hmZO1cy+ZpMKL1fBp3JpVYjFvRgYeYUHI6KRzTqrpKDTzXM6/Dr+sTb8S4EbnyaUwidsE2a8
LHdVlx2dCy+TIe6IgbqjNlFeO8E54j/+yKOhiZDGC/NWD8G2aE0NwA4nX66U8a40vZA7bpro7Q5E
QeQOHrOYJe9Q4ZQbBYzxHS0ivY7fajZI+LdFtQl0EiE54zu2/qU0+VBfi+4Jc9Om6p/7kPT/mVfD
NZCgziFQdFOnccPQIRAXSCHdxYwYzLxuYYal4YZ1TXEL8/LRtxbUVg5fLOo9Z5CmLbiF8cbq/rjo
HqkxeY+wjRnTk+4CAIwzSfBj1GB++hLwxSf17H6+4kc+VYbDv0eMRA1T7baMLKCzrkBX8JQwmX9A
YyzrDz4BwTu64H8aXL6xHcT91w4JUfoERFjq4DeTeBa0qucWSTjxfAPj8sqMfLHOoNrNXrI8EUSs
tR8McCHu/tPAweibfo+D2/1nEuYcxd0tnwY3c01hRPA4cESYX8fyejBtofzdOk+QJv2K1rexkRHA
llI30X2iM2x83v767oRgTbIFXltuFOxs8RZvOdEp8Xll+lGTU77u7V6oSDx3CZBHeJ2FZ3Q6vmk7
aYS5di0vyq4pzwSYl+6mWhRwUuQEPQNBqqmV1ATux5KKUbd6URIFrAaosq1mqx4phGVMLhYLYvIS
QQWwFwATvoBD9CpwpEyRpJ23zMTYKMkAdkigcjJ6MC0BBf8jae/q1rv3v6ItK+3CX3lj2ZVqt5Nj
9zX2NG/hbx1AX4e+Cug6Opx4V0qmqM9yhy1Y7X3OCsZ6506c2lv1pcU+YlScBcNVWBA90pC/HUvN
hVgeERTnNW+vl2ek0BRZbWTsEYcCsd7dpailIwMjJkFfVPDmh8YQJjuGZltP7l8cUY3AlCWudyeT
2/13eo9dblDgLC2FNS81l+CQfX56Qx2g9TgXPdmMI2gVJ8afy24OHum8QUEEYUzBXD37ARygJZHX
nSsYbGmUJfxi9ntuVxFyqNhe51/ICg1On24nOVTkEnFdtMMiwk8LquL9+vGtUQD+Eo455treYDod
A3lE0MZLPTbaWw9WwVaybFWL4MnvaNWB0MrHuuJ+khM/vwDatakxbt5Sr/gfXN/zyxUSbQe/qT0e
nGYtPtp6YzicjLGmUWKyKZe2nERdj1XCiG0ptsQknnPmqOSc4JcEiYLG4ujAoPETnBbKsRV9aXKk
rsJN5B+9L57DYI11fxECqpfw5R3k5b3nNBUH4xupcsTQzyafzbwq0khGFjWcl2xqM3RS5Nsh9s0K
FyaOLmfFJ40nuGn4wEKC3QUFkbtiEQMqjTvFMWe7rp6yGBqZVEqfRGigejNNO0hQ1ZySAg+9dyFD
OawWTlKv76EvmXaipz+kI+efTFnYGf3/GOYtaFTbMqyYV5zLPT13CddpX9HgCTPZZCBF+pxkunvG
dc/W5b8JjqMrHZ8JSORl8uMqeGFI6X2jMU2HnhnOcqT8PX18UAlc5VXEWS2LT0J/aE6EfDVJx+b6
7iaDGoJ/cAJh4pTZRgYw4dRE28JYEl8qia5JX3HPjf+Ebgi89piWpVuYzpYX9CY0z1tKRNtbTSW+
JRD8EQWA09gv27rSQ/vXc3t3j0E6PTvpePqryPE9RQHCGWg89wJfFAcmcKkRJTTpSfThEVtkWTty
4moKknkB/5JIIRZ8a2pNftwnQRDvvSKz5wqpeLiQ0DSXa2TxplBG7Fn6Q4LE9b/27DQukSt7LHAN
TNrun6aoQl7BwIgokJR2u7wvRSq6a2pm2qKatgpFS/RTebtoK85coxOKd0Vs2UxUhV3PL+0b31/t
TuDZFFkLT2KQv1UC7/Ss5+5Gq6KVblytQHYcPlmK29h66MRkOEyubgyT7C2qnM/eiboVNESAPxCJ
6xxcdGWDS4vEp0xkvlsWurbpjTfAynPr6t8ArAkUykhONO8pTBtmKLAKcAp7JRejoDQhlCX4Zuz1
thO7YQcTsnfiQs1KxkC1OHr0IUHYVqo2ZFnkfxTAXdiBbySA8xsYcHDhzGouryHsgaLIEIRQD+WP
0TpC7W+ym+fwOr41uaFGi7cxP4xwJacol9qidkt4PqH63gqN11wc/8cbrF5vC+I0a6Hw3fnVlzxs
ormJPFx0OY1QYNYFoQshyRgEeGAaO7OOB/U0lkw5B+KUwUzi+iNbrfRynXSUJWcjT/v73MJzCub0
qAkut8q7Y26gQCTWqJ4sDI39Qy5VzZzQ713LEOJMY8OOUaI2rujrSPxQHfOKJ9RglxYhh0lBikee
mPdsP0s3AI25Oz09iinjkdkTS7yCxD3VReCtnJ+W77TeW6krDn+BMZiMG62yHpOyQ4PMEUGG9Uq7
MUHs+Uy8/0O6QdEIx0wmKbzgPuxm1D6GbbHJHYfljw00yO0EDtTbIJtq4REIp02x6EJQqAIUbuKe
NKMMwn0eJbCPmJMBfpxOO5QEYuvVvuM89D/E30pftLIWwhA9H5oykKnZw/DtXPEfqsNygRfmNU3U
jCotoE45KiXh5nQEoXmZ7BuQQA0DS6pq208+/KFp/JzK4E1ovF1KJOkxsQVZLC0OB7uIJjYwXoX1
2gXTiERGc/c4rxv2/EF1aQlfVXA1Mv31W9EftKJ29OJVJLxTLdlERzuuFvMGaWloxsTc+Gl31uAU
b06HzrFUfg989PrkMd+pK4hI1wVVQa4uDrhXBj85RwxvDDgeZJwnrI5JgW7O6NCBEuBSOZJotaQG
0S6+wd3ygAx0FulbCIQ0YAKeTsONRNs/KKxmBzwVt7UGVQR11fb/S8mqbfR0f2YzQhEfXuSaQDmz
0uKZsUiGU7NHqQVOplM2KB9Q0C598HXSqNA7DEY96INv5+nAlAvPxyO9om2p6BEev+5GRuCEoC+r
enisKbFWQfvUwpe/J8xAcWmDIeHtVqpEmjXPGy95euI6SVeUKaOvuVodQbBd9YcPwtGAKu0MUCiC
ZzUMoVMGkGK5XnxYXAHOQCvFsqHjGI4ED/O8YKdpy9ADfWUMahtN8f0eCXYZoeobn99iLcyeV8Yk
6kcG8mRvfmdZryEsxVBhfapsxaHo+i1Zr9gmyieIongabDY2DiXmjGvqF303411VMXX6HykfM3Zw
w3DDqa1j4+WcM8OHQI70M+ABZ5S0fIsGqnpE3laMcW92uYoaX2yezhTaEEabov0lAC7LjwvHn+zP
vd8tZmjY7oL5mSiVWQSdRnyfY87C7dHhR2WmUMNPGlMTB0m1uqZRCsU51jxiz2yDc/MZ09Uwle78
DSKMR4DcVFgTcxipeIYmAhj2DnD6qtWoeF4oinBZyQcGU4E0U+qKpUKwkvhkDYLaJwEMnqWVqvk7
KTr8AABQ9fyDNQX2ivTbtoY/ssTNCTvlJ8qysM4zJBXyvg5kzlz8X9WxvmSLBJC/Bn65128E5W2h
GqAajeKxrghPGDS5A2+1FNHG10C4TyJsjEm1B3fSuS8gFDgPmIOz9dknyJPVVVuTx3xnCs2c4WAd
GZlBekTxC0C94zyM5dkldNmQfV60DWFJOCqP576T4yO92b7hKqTlL5eBQ6xmxGLamXNfDPXdFrk9
UOKt9YIIfk8wH+SUFuxfJ5D2nxxej5O+YaSadaRBmp6N52tH1zSVS4Wr1tdVsusRRLCXw8KH/cj0
jPm0AVZnx9lCOBqlg0As7TSqoK0OyrXCXFjfunBDRWL8M1bjDFbyyJae6BMxlqFwRtuQuoA8zEG2
L09WQkMZ1J/y2ZgNI51wjdhX2MDeQStyWXCRiS26bbaUm7yX66hyfua/BAV079CXl6cFZ3uZ1NLb
DVrUB2vcnKSP3BtrRTTBmvy/mHuS9vC8Evm20qO1ZTa1LpyOb/D4IMXZ/1AnKfSOx9Xh2j76i2ZO
zgONMq/pU9FLzdynyGDy7coopKx4H4//QfOiiKahvLzBzlLa+ljKXD+eO51MuujLs1LXH7tstLuk
ljyxjcjpMDvc6ya4DbLVmY4Q1S7lnhQD9IZPCOMK/mpvCOO1KNDjzIFnHw5Z62FmjEkWjuJwQHsk
3BRaVnUYg8cahf0wX5S8Q0+1HScso9x+tVN3izk2ui+FKJdqI5/gqZ6YyZbdgAWCRRDKrRS09OjC
dPaiqGrEL5qpjqCjd0b6+8ZDogSHiKW9tpV4ZA5Uy71/y+Iv3bC4fQu73zTEnrCqc0kwz6XhCQ6R
+wC9GlJvS+im1qezS0hY8JyAiYFG2TuPxw4mCYf65CZJhzzZPUh+IJOmb6YqXxdIjqXHKnbAWoNL
7FTEp6p9XIe2cgLAZxAgF34ScPKoJjxUg7I3UyJp27IRhgLWq+fG/QicYYcx3wzYSCwoMZT3t57z
4HgxhbOlwg2HNClfvcnWr9GIiqoLl+8J2hcsF7ukPQUDj9RGJPjwVuaP/6uJfl0jnYrNGS/6p2ws
6DQ/xRV0o+R6SJAV3iN9/fZEeCWFRoB3OzZHqIqOx7P6DZK/Og69NX6UTFho2LSsQYvx6mXR+exD
Kvm8xuGgrTEs1tlDlNFL1nAiN6JMZRcWDutQm2dL7SOrWV46KsuEBkUSsze8AL654U/Aw8r85th2
2rU4z6GGJ55HrId4pBtvK2DGkLT/RP/ypw+PRbnPvE4Gvn3+v6z/2yo+Ck1rlB07Oy5LBBqlD10H
9XTyQRNUSGujtJvsR/BAO187rFKVK7z8IgrPtQf13srveZOX400qf8eM1f5mYf8iCEXP1oeyqBNq
nQ9hMko0qlgVUDDjkgqYzdvCWHkA2cW8mC+JgwZIuN1QHeektRiUIGOwOdJNp1pJpDkSQRpZ+gOx
1wfbA+PEa5pZpLNU9KF/nLqnpW4P0P9QnyxJZVMAJSMdXrjln89MtCB2ESKaXVkEGQ5FWzlfEvwG
KXDYxIJV+P2pht2kxknSviGN+3uPbjqwn6CUN4/AfI9vR4X+zRB/YZdaYer3ZYjoErMQABC4KQCJ
wb4IohzAqeKwM/VfNODd+ZERAdYqFFTFszq2zBQIhum3bkCbqDSD2/jJyg4Htgukckm3mN40+5sM
hiuE/kv/HdvnSsfQQ2kpbQiNCfCiEUS2lv9ubOiTx/qd5YiXo2WAL8ixlRjtLDrFEz8GTtEvsM+K
Bc18ppU6usY5+cp/6lCEVjND9J5MAP6Kv4HZP8Mq8lTMS7r0bzOw7PNOgL9XP9BCgYXz/idu+2GQ
GV6Q5ToMJIoRAbsVXnIrOdQeAZw4/eQ7hGj8OSm/Doe8Vm76DrR1LfUakXDvJ6OXtbpd7mCBP1hl
6Q6Iiwkcp+aT8UjWU3bMPyZf73QncBFU/c4LFhUeeAB7ybgr1OwUaII8PxCWah0CqrDI97cg61Sb
DRaRH4FhS6hq7GPk6HlEGb0Q51Px9VYD8f6JrTUlkCWROu3rGWI3pHaKgI9+4Lz9XnhTNxY+In2P
Kv3DCzrQ6RAFZ4pQ8lxlrDU5k8t/C3X8Nql9t13E8i2tfcyqxy1mNRkDNaTzNPilItVesKpkbJum
1c6I2S2+rkQIAAxCldTCEQn5bfEFDHlohLtto7PJe8sJbjh+UbIf83uzDuZFYUN6khqlaVjbr7T3
QnuMINsgkgs0uVtPh7d2xNagieXJ1pOmzR9w9+kRxNNKG/mUrQPsLKWpgqi5Ve2mT/6Sy2ZnTs8b
Xu11figdaWfDHFOWsNfLkgt9odfryTCveU9WX3IPioJWZH/zoc2ETg7GLl+NzbxZEEOzBD3z6lCI
uzccIIN7uXFHdoqRdxiSDMR8fcnDW3nO5C0UUA4lDQCd7rRlSCt1YfvLZ30v9WqRmkjgaS1Why09
z2eaFI0TZIMP8kxsXxQpvhY4620c3hvy7UnPQye9E616GUfGrriQfYG8OJyL60j3xs5pYg6QDroP
sMCY6BkrtyLkP9u+2a9msqMu7lN94qpc/ZcF98hvZwEH6MGx3o/Ut1l9PdIJ90VtqO8wc9/JXSJ9
xAAqCpobNBNbdxY/YSNFY5OY5wLaCkmPA7hcKkp7mRvW7u+kU8ZotG9cepwJyjZjA3KldJMwQt66
nqxnmJs5GBiXMuF1TY4AOEkF4sTBL3GuL0iCOk0dnGKdO4Q13W0fo9wqanHXwm1FaO2p0it+VmkV
fdvYReqo26hsyxVhhNMl25cJsNCnIxwrMRTAx1ZqXEy+h4PmWofkI1OqOGiMODjoOyTLgrQI/RKR
xkcRjF3w4Kts6H3OKA2CWl/Og7dKQf0TjzjWHJwSSD7MrlYGnC+bFjnzwIBVXKKrro0o079pUzzz
L0OsCrfuPvKOXV8mnxNcgh+P4Agn09gHQbjocAypKyPYVHx2WdSohW55Ghf41XJn6muID6tOqWx0
tXNMBnWAcRok3jRPDnSkTpZEHu6+4UIamkL0DCwlkuS+yL2Tf4eSqxY5Q9tNaTX61eN+ZNXJnJ9x
Iw6jDZHfQSgXX1nSsVwOQrUFRpNkHjyeP5ADkd6ToJ6sowni9A74IB/VM7PFnlbMz3KjoKg0aF+f
H0kf5HXTV3JPhvfoZBw8xI1pGn6Gy64Rvnyfb6tudYYstfRNbz732VyvWWlhYCheuANAPp3RvbcE
Gw9e5A/x4y1SxE/ku041ycYtnlpZTCoyf/0MKMwljbg3IUDt6rw0RHvUxUJwaurK9pBB5xX80tSv
AZwrzWHHW+sBdMOrssQ82WwPoBopQ6SXujhp40ihmFL6wwUR3W/fp6vGG5Hr2vMHde1vnaUqAVqE
OF+0iO66RaAJLS+Pb2kXU1LJveB5FwsAGkp0jKktLqS+rgg5aG/qvsfn2rcHJm4rZIQkNIaMuatc
0gej8HfcM8RoscO7Bjfb5vwnSM3lO57DKaj/Zkc+xEThTeAUE53/K8X6dlSboffeGCFXTK8VJBA0
/THHbgO678+33cTQy8XaDfTohARnPcolFlEue8G6bFwPATx34WgiDwC8mQlQm4mrUhHS89o5lZIt
QQymg4BmlDv5dO1R80Nzu1ozzBjVJhTfmATwTJvtstE4C2rRKM0ihleNvqN9jtL47eDCVTlGY9Fz
wG84DITZ5noW2FWRy6L2X8wKOqJahgCZA9216nhM7aDWdItLqCZC4jnDzbWaZr4h77sBIkFD/SVv
VPLK5zEwIzaWxVHwJGuDgKxOaLazR2jhTvVWQVssWlQ8H4HWq3OxmEItrIDMVgVmEWHb8+9Op9Lp
Jx9sm2lFr9dAcIhUDB3qjeOuJhps61q5UiJU4NzZkk02NGDDaM2PBnQ2ID5ivazeZJ1KPxUQefg2
owKirB4UANBJVVgFCMps+efVOS8olS+I3xP8/CZM92w+h8ZZyRRaphI9RpWswj5fGS3FEqlDKe/Z
KMx/4Rt/sCqHfBm4/asbd7qvkZK0mHHGK09UaKuUJkS1k/tE9oPAYLTRpfB8VwGGHvar1maHTrdD
avq98g7X0uklxFQsyt0KBob52jf6x+C6D91zZc9vcdZj2LrpSaqe8bjXLxxlsrjgNIemkiHxWvBV
BZ2oAbCKchtu79RW7Fkk6PTWtf4W4KOsS0nIl5vnH2UhLWoKgDuBd6uxo/Jgy/6A0vXfN6ilwsga
41cXu0CrVVUxEM/MbnD11Gnl2xcQyvLhl5fHnp3C66B5EhqZodxwl1Pz9/0B5fLP0GIvj1Lwa/DE
ZtAfT7zDA8ERWJyk5vMavw1V/5a6yIsQ/+jtnIR7McHeH3nkcPOqc1sc9f3c6P8/D32FS/jBWBub
v9YOtg0RD9OjdWSBvvS7eEoc1yE99az9Mk7jQ12+JeXtsvi/O2MAeU73o7FmL7FCwHruHL9jcObG
2pgWSYICrCLuNwQQC74J5awzrqOgFmzhKuOEwMqTIdaB8Wf2lCPWHyCkcVPk33QcdC2HwAYGL/S6
aYEx0S0328siV1IAezk6/5jXwNIrBLXJMrGF8o+/f97rmb1yG0XFkW6fB8FqtHz1f10ZNhMyqbHw
8KxGf9z4Ym1XX3/AeX/HjwGHvEQThFejTqIDrJQpWU3L0WclcNxszuRuAa8f92EnDULuYzDOHvbO
U7RuIma5zCc1FS9zF45g41sYY9FHhPSHqyrWBktvQWcJrGbuhbrHPUTl7VWzDqTH4P0lM2gKhUiL
Ks3rWo/AFLwPRSRXsySmcj3mLDeGNFasIOm2feRmmIkgjcairEaT59FsO1BBUbXB8IV5DTqhRvyx
EHnqivqHEhrW8xbaoHo5ChrCCkZbTld2INCIBQqo4ISzCLq1JfzOkO3mcw9qXS4aJl7jSX2bb1Kc
mebezmSs4nzEhmVVie49twxoNAluXXCn0r2QrQd8X6CN6YL+fdAYcxy/g/WLsFiYo+DYE/CvO5F1
zftpxCWU2TNH/9+S59XJzbTxMraCi1cSEzGMTQEno4xbOp35TBso16k3kXS/MaTlkbSYG41sw/7Y
mV4PoTRNKgJ3xWFuwpnQ5kya7+bl7mVKuVMkaYTrVZSR4Jf++kqKsESaa85lBD1CkuUmXm+Wof36
6gVvWwOZ09XnAHS23r2hxn6GIK+k/TMsBK3suCJj0Ok2JMOpPkezZLpjdUdKwcBRvlHP6W1RM8dH
1QmdJVxsu0PFODr5SpGMFpixP5aNuFOGccR6IvfmmmOsaKdtTfJob3HvW23BfyEL+1DUCPIJieOR
K+wFQQRrby7rAQ6Wwl/imEAYx7LFTG5UM80ZhmxhUxp7Eg1uwb36kckukr8c4pxqtbqjjc4bo7A4
qc3TrqqZRlqkfWrccIdNBjAcuF/sB9lUaom3qMl+idSNdJ23fy5j7+mlPZQjaXslN4b5/LXxbb6l
wvclxawyrc30vOUfBP0vZ9qgfBkUUN/QHbVxzQWLnVFregofL6eumHbEnZfaUXT22Z4nNlwBMthE
oGU+6LkM+iaGzqkQsgEXzMUJOa+tqUezwGw8THexlAaZDYsfmLbtY1y9iH2JGLlTL79MXF6OkYhd
mfpM/ZYzmZIk9iCwEtA1FEJTGo66BobZW5orAmSYTWwDMs9RcsVgKjoK6O1q3JQn50bXyUudiRZe
7PaZrdIRU9F8melafoZzmKgs/ILDmd5oN/Qnw07jdE329E1D3n1WTvHTvdFBzKqR3dqQ/pSLVixn
uHYyhjmRt9zbsMtlQrFpM6dWuwDgN7eBIt3GsD1gthi0qRt6lCfylRkyFGYxvu3n2MYJEaHT0nzE
vDUouz/owCFxhuLWLeXQFUwHBQwxEWYA8nO6WKwwsCsHDXf1289v0HnB8qqWpHHkU7pdPIhUP6sq
Pjg3bIdr3MGQvEg+BZ3vXAJiAaSRdlVxSMyVh3FYKvK73LfdatBU+n6mE0qmoCqDKfd1NDYGXEHl
U0kC6JV7Jsyty+Vy3wpTyj9AiTKQ1wp/mZ81fe3eSqaG/tsJFEurShmRDvBIuWh60uz9ZtvFIWDg
LWrnGrG7eIZbL/P4NSnV27q4VTEGbezgsZumGvOuILHR0G1dxAnJhbyDIwnEmd9L6tly9GN3uKux
aTxcUT9Ug+d81pkdxoFSMS+OUwvZS2ZgfIjL9q0Da4Y6sE6mZEfZoMN84JIsoM89MrOTviee70KH
9YHOUc3f30aZSUOCllDhn28l6/R89vg5+Q+okCYDWSyUpZOcNVZAg4q6S8lJU9ldId2Tb8ghyUnO
vTmBe045yo5HAtHxye+J75t/CAATv65nLd8r9LLheGyQABGgOjF6wuW2pjJS3i+1T2T5Xa0NjdXB
7aCOLOA4xGgV0uROx+G1C95YIlVmw3rS30WXnaI1g4gzISfwIQMpBbffGmCHrMYb4/j/zhW9uinL
WrgdOIUP1+jpqwvlQixRCYIdcLygMkBkOm00j28jzjVxO3TtWhSFZvgODvFEOilOT/qp3G0hUUWg
hrQ2eD4H08dTatjIV7fXRKizyKfHWvHUcdPgWVbFvO4iVzT9/koIh6gmdmtRvSddEVrw1jbV2Z//
xmSa5N/eQkEQdKPl7IQALdonk0wSHaKw+HDNc3N/Z5dbJj9dQtVrHdyGmE/pPHn6o0ZFQAtYHGIp
vO+GYP0+Lo/6fp1dA9KjKdK5pJbA4RSDjj/juxGExE2kLf+tN9jyiWtHTZHVuLcRND4CA7AVGBhr
E9b2zs4Ebd7Nmuzn1fpIAWK9AGuzqThK/5n7DCKzpiqKC6AeXrx8O6zR7At5iiveYwgo0p1MUOPg
IYDxOYy1NF4ntsqnOoPldQetowNof1FENc1HW7Ixq47IjXFFcXRR5mWk6tDLsWUVDGHTWuINwl2c
ujrUVcv9bzR6/+cMKiCfS+TzdPflOBfyOpyvZ4psqDDEY5hsNd08wC268LYGiVo4Z6g63VhsBkUJ
S1rVc3Tc91+1bTzX9uZ4/1/EoEbK0B7+ERbmsbe4iP8W1xeG550dGoT80sC+BKWJmt79ynOf4TSj
YSdkIfQa7YAhIoQjl3697Kh0oOHcbwciquPlCiImp2xz/V1Pjb6jiuzkt2R2JgTiBJOS8fvu+K7k
QHVZqbjUvXvdnIt2LNO0MaKzzCSpxl4vCX2+nZDvsZwWzCV4r4SsDWzIU8Yz67Oj0GLdBFd4abym
4B6v1aSd1jXlsDaQlc4odo3K09XneyGqg0FVtw+fYG2MwhL9nE6NhwZDouBR0rlFPEi7JneqiUn0
36lnFndpEWmJcF2/UBJgj+UvyF/K40M/RxVgKhOB16uAvvSTVjJSObzdGWfxnQzjlre/p2r71A8u
lgjhvZ9MbKWgd6bZLYBtdSzDb8MsDWJyCzJNA75B9aEFUdW2JKK/zUJH7k0w97Ef1WnrMgkGlF02
dVnwFmPqw6Eqf/njcMbUUNzUlt9+o3NIrtSNwSp/C63rhyUDoY3iAqgqbWoo65L14kA6VbDbDg8+
qMlel3AF6agkIkZ86kKXgaOzU2NCF3q29lTCtnSbCT/du/h4EWLY3QwKQ2hocb+TwlZL5luiQHFs
V4n5A6CifAvyYiBYA1mj1CuMYZ1PpAduKSHrPND1LtlE7F4KJ3mxGPoZwgxajwujULYUPipilrCE
1XXt0T8YLpNpYMR47ufKsBcC54h0qLkW8O2nLpqi/NcbX1eiZilfaNRQXcItHXhe8T2yPUJ3Ziz9
Br38UQ1i1ZGkC66zMpFe3Fc5hCAtFjdYz5PTd7GJTEaOJ/OF+uQXIoimFf6bYHadyNwwsFtDKKXp
T2ggvke+7id3K3oJfUYa82FOWjWIZUm1+68dq1x0CQ5xnRCcb6Kxmv6TAjFxDq11xNh/ucuhRoI8
eG6rs+eQ/8GaXo1AM3La2LGQRhDIYwesxY8I4T/KU0j5xMtlKpElMI+0Wcs8z2SOp852mMAwL9DR
mGGEhBrZlFQSSsTH42npmE8PpQuEMfyePfh7KnJen++67BRY6elnNG4zG9FEnVVHZmYp2sBkxs9Y
bC1o17eBknhe0htkMma8LYElclaYmY5XZjKBNgZAzOVEMjMj2nATOY0f7YrptVu8zPItdGMyQBiS
hRcRH88P3Plv5/5IEjPesqIPakYH0HdeLq1U/DQMALRM0kh8UKDtf3BDShiTLrgeKhUvJl1zvHhL
kO8AMWmFUpnN7E7ZJ9Tp1SlG7CYwaGMDjSs+2BloPwqFKYHpRtZH9CBzg5YeT3UWYwEZc0Xrzh6u
bM/wU8RDYIgbrYO0nITtbOeY6vpvEwtl0lJ/YzwBGklI9pQGSr2TJqrsEthBKZa5iHf4Xn89sC/z
OJIXRqu3wqW6q8Ga9FEzdLt0xqBAw7kpLbD9yEMZzOqRD5PrZoUNGfckSoK08dUvu0AFNC0I1f45
QB9/4IhSiTBABGJpiRBBtSf4aUzWmF66LmtlQte/q6Y6BcC9mnGEZ0YrPgWVVBGS/zf7li0dMdib
ufIasCkJWMWSHq7GYRcJsU2yX4WdqATVF9v0yfE0gp/sq3nMvzRqMwRzG6r3t1+Q1bZoUykr15GC
faJOZnCsJZr1sr5U8b74c0JqvOurq+Oejjdm1LjsMwsLYz5ZhIFYelz8avvUHUc3c+L4j7wv2UXU
x0hzcDtKOA4wzrzvqfimiiQxGPKBCi9U0XvfVavN7+uN4oBtOePzGUVbKZO3qpAQ92vUx6PHAPWs
SwS4UjEqwU2gWT/W+37DOiWmVnP6gcztqaPuBy6P7FP3xHmsJzbt9UJneKberOAiGtUeenCwmOUt
CZJGc6GQ5pRaB09aX+5Gk+smm9B4qkOqWlLN1aPvEbcuzBWURF97W2mxJZPagTl2y1OrMgrtG7lN
9pA0FdBZ04sNXwoq98G6NknrSWIu01P0SQSOTnFpzNYvQ0e1jZfxR+O9fyNVVD2xBujAa4eDh+ub
oX4cfeJJpew2B63/pAFWw/U2CU6q5Fh7P+GCZbZ104V2L641hDUazJn5fcwbTnswLMjDzASGvdgb
l1AJXHaDOSgJ0UAE6TAl1teykUyE7qc0IDqfW0J/8AExywfigsovpFix6TAjLKKgVnu8HJnZnbgk
ruUx7FaqAiUoGNR21OPkWmScjyFEClFc/ZGRdpxEkIq7mwT5hF0GuaZjhE+jLeQwiD5CJ5I6+3qi
K15ujf0qNR0Tl2Ih9Thz/baarTLcrT6Dv9tNrI80sVYOCWxStuxnRABf6g5G4NgnuPgJwHwjn1R5
zd1en5OG343BM4XNOJHOw3WgZpuZcLMjJC7KPwAdfjqgPUzyMfzM2ijOMsNjpjoU2vkA8X+160pL
1CMxAmKSkW81UA/g64Xb2xWiV+SmkvwfSnzDXIBV70LPrwHLtkINyFJL7Mpzsa9gMJztjqdkelyC
oITyIzKhkZ/YeMMlCE0pGwiLukCyKj6IgtiOejFncQiVo5m9mmlEfYfQeTpc8nTpTsA4oWz8DNCy
7eyiuxeQa3wQ8oQoiJpLMEsWWVKSz+cbWAhcRpt6YCx7rT11Xgw9aOyYnjlsTLuxK3e9g7ppsSC3
35rqX1vxjvvtGEmB6gnMgGfuUm66d+ftWaebv2CdyzJa8lOgl54Hz1lRHFy6aO7Ms0R0qkeCe27y
Hh5zwjdu1a3HC1bmwQbHNkupMIGie545a9/16aY8h8Yl/HiSDi0oU60DE8ni+kOOpJ5duCyIwjmL
30NqjXR1PQAuzOKg1oNAxpN5CSJBvaGUcRBpfneygsvwBjP+rZN4liEymLhRpA6aTnr2yWByaY7L
5goFbnLaXYgeYWUYYh0l5LCE0KDN9704dg5LvgBaYh2oW37j2dJRgeskjVG9eLxTFIQ4rsBdNEwK
zNwz4f1OvQv751ISBRqSYQQnT0MGRXl6L+YrIRhFlY0LF9CZBYi1hNsviWQv8694NyPMPqygHWMZ
zibyTYEIOXLOwvVHz1WTDrYyzxiRubcAXxnIYFjOVJchIncZym8yN3Tpyn3YFiM8R+iON3uPINI1
70iwlly6tzt6kf8xNMyPXy/ZYEuGGL4xvlJO2MgRJxOK5cMs13fVsHZ3F2s3BXzKXGvMAyj3zBBg
cyKkR+ABpCJG062ZMliN1CrG3k0fs/vyotzBFgmZy/hR/ryrr+RIS8Ld5tQWgureoPN957wgogtM
GEIhTMV5vIasClRpJ5v5DLPt4Ii/uw18boRrgBbh+eTVI5BtkGj+Ib52GneI8r14SFB6rZ0PBdyT
1LGwWI1f/ukdtAsFy/4yej7f7c2z/UxI00XSASozaa6zQDfEkQvq8gRxkBoytqy+uJ7pMWitgOUF
S9k5wGJtN3u5uWaYPpiveJbCBdgZ6zcgv5ENmvjLGL1mtdt+wN9cp9W8f4YWm1o2oIJgXjcijBiz
dzLHlzJjCiDwAubJRDB9zAVzlYOy0Gn8zwOSOaMmvVInzSuSJKphCpI4Nw18nNZRVbHLe39IdkFg
X4H6Nr1JisAm0FFyqKsSQGAOIy1aR4ewBPkSJamuB43RNce+vmXhdI5DTqUov8ueEDalkbidqvbD
5CHTKFTNs7d1D43qUZCqlpl94Q3M8hwTaeG2OYmjPloRmb+3yslaKMwfjJlWz1RtBPJoKbmwnPLI
DNYLRfsfYc+bCx8uGPKA0Sax3JJwdAf2AbV4G6A63tudA3uOL/Vj9fV+WtrUmUywGQyvoCkHiHmh
mASYbgGeMoyrqkoQLcN6OK5/HZPZHWOluv2A69gVfOHc1J/fMBqAQ87nrOGz25K/PIyHapmY73NP
d3WlOJPDRQKuIW8SCf5ZcmCKbGVCll4DTKSiWsaI6XS32DAeuCkWcOHjd5Cr3cKirbD7pqNJIUIG
D5xkMElah0HmPoN7nggilqfkG81gnyYB53TgJyjqrIVJLuPvnii+AHppciil+70zbTl9jBaP6GaT
4F97WuEeqNhUgL08uPVKkvVTgQAvqQ8yqcUC3Wcr7hFx7OPG9iQxvXdYESSKNH5AIfnBPI9g81sQ
tF4h4HLT9NtK8OVUnTdwYeQZryoJxcUAGhXSs7AExUcfUVdI2tnU2ySGvLypNrvKxo2NQJpgLwgx
b4IY47Jn6yJJqFqT74BpHycQAFDlf2I4hTwhsBT9O8E5r7X/BhZtpJYgObps+3ozL4n0wiRJXka3
xdX+EtIXaVOhKOngDpkmrKRnWErUqs5M7GBXvywE1xDiVO3NC6O7wUUAV0HqayVTovtLmPBqEAwW
yZeULQnqIA2X4R08Du/8gnfFDaZNS22Y9r4k2T0DSyY8zvVSQwNiEnCts0w+KQ4LitoeCJSU3jbq
2Id4H6KvSxSsSBQN7oSKFawTDs318szY3o2Ti6vmJQ3/CsYQmI6jzsSYBK0hMnpVJFlHuXqL7mtc
IBhzb4+Gm35aUe5aFU/IjK9chwBotA8Lq7CzoCTbHXFIw18uv5LObBijiNxjsn2LBtf3UkGEOAVg
1XUdjHUJMQsMJt87tgB0d/auqD9RFlrPb7+/wvhxvX3gJb6XygjO9eRe+isFntpWheCsjmWB1JDJ
AirzTdGevZLAcAr04+5nKvCfgyDG+zykuTQuUsPy7WqkFrX/uf/aYvQWbo1O3UwnueB8kYh5pgV7
6IuJSeQr+k4btav4AvpXsfaxjI92Q6UZss4kRIgoYKtBbSdWDgrH9S4v3yHYiQbBDu96J0NsXbKy
Yas+4YbLKOl/AgDb/yGp6iM9JQwYPADV6Cht7DaTVX8Pj7DFcZlBPC0vqmamEU4tgV5T7H2l9X6H
dnKroaKnWXx4PmdLJHtGJlZlTSF6xUD6DOhkH9QQtgYC6yNVGjI6wuwZf3ixWibunIHNbJyuXYbU
Xu6DkQI0HIaTf3PUOSgsZBXcvAfquv3SwWMnUM6tlblATG1KSfqTu900WNep3cHNH7mSkMELr4uF
uI+A9LVrP9suT51BpMb0d8Okz4Bp2jhMOQiEqgJeQoiH78fg6+sUMbe/Ix97RmrxQ01DDVjNIhb3
e6uinJiQxBUJv67rKcMStzvZBZmHzOmkrPlvy1RBmzBhxwLviTd7M9E5vTy4gLrEkXTuVykAkbnl
v/AB77AFOFjWOq3aAgbEzgNzCzPlUYcye/UyHG+kHZvQn0onpHaiDSK1U71An/RRWo0g1b7mMI2b
w5j9x9Oz4LovAkvs/Qb9hXh7IUsQo0MLC/X10JExISnjqjhcdLnDC6to3WfyV02rcaEvf39+48bE
YppIWRkNbm+LL4uGyKax8IES5egdtTIbmzFp8MTixr+UCmemBj9fmoevGq7RP2ciYS8ebt2HQ1ps
pt4tEf3tDSeiP0h8+vdmhWU0jW32drUpmoh2hH/iK8HBZHksHP0j33trXFiVWad+ji1RyO8zC9ay
cbPiu2CcM5colMhcPiUoAoRBZxcv4vXSmq7ltuGHy5NVcD5zl6GmqtLXV9tp1JXIy2e+9Gef1jGL
9ZLOWmaExnyxk2XC6rugv0rNGkGLAEciKf12jPQ91Ui1dmA1zZCuLQFub1SRP9lqG1IXaUffoQmB
wmcEofyWLtPUdu2Z+Cs+QV0Y96DPUpvMThZt+nMOeqExrRU1cksuIJENgMCBs/kxbGsAdTJFF+3y
K3bkkR2z4bmFCY3ZjikdIHEUsWTd4AdIUX0i+JJ8ozm8VqYm43nm4IvYmrQdYQJgJv6slWqr+C2i
D6AYT8C37ozYcnacDXwJ4iNp87tC0Rq552oauayvgbvJuXphHA1+o+Az4w9YMwHPQumfpO3PLS9T
k4RwFHQK4UeN2oTFQ0f7lxBxsGZp+rCt0snMlGsS2Vb1l4FF1IbyJivGEjsjph7UTFXXDLtoyJ0Y
LyM/DV02hMcOuBCVnpOV71V+ffGteId58Jx2VlvlNM6IT+3QdMN7RbBbhf/9sxgV74Ej6JLf+7cr
3h2jDnQ9AdpH6ebFMhYdm2RG5K/PF5f1nVtmYU/LtvWMU18VXbhF2/qzzmRVs/nZAFn1YlNvg/1Q
W0AVMLgOrIN1R0rsw6yoTHfp00xKvhcIZk3PCRiO9JeFet8q7g24W72SoeKwpK1pDz7FjX7bSx77
yq6kKIyqrhZQNkDpUI1hFm2iLRxh2Acyn5LRMdqGz2z7fOaLRDyO3ciK4U4GRcgCYrO5mq4M1MHo
Ki6z4Pr4eW2jRZuGkPEn9qwPvwz0bxRpaWW3KyEvcb6vcgovO1BTFoLxclP7m+ha/YiFVkXRyDSD
Dwbm7tLKu/yJONFdIR6gZfl10ijK7fbqJ4jxURanpybPu5YB9bxUzXgZJa/2nkOzj7QrISojc6+6
X6I+o1tA2Tb3dAnvlMfaFHCW3N4zjI3yC90RnjLFRNytQE4PEHryqBJaPJaTeGo9psUN1nl2efez
L9HWjfFOS7HHKdCnTSi0zuELg175FEZuNzjSceDZiMjqI9QHpa9ja+wLK0MSsTlM8s0OAOSJxN3f
eR0A0FieVLd/rEYkqNNdVc2CT2Fk1Jcr/VUCdTOmTsKDqH1w7h7q+UmrJkH6Rw+8seTqh8smiU1E
P4b0m//5o2ZQ3UR9jcOeUgA2MCML9NmHYS+eRAnCBoiFq0DmjpNi/Y7pwMT7SVfbHFa7oaiT5/X8
DiMiPMY0Y21Jedmeo5PoYJHx9C1Gxr1HgEzs3ljCEA9RFlNuLgPy5JqebTQ3C1uNds0LhcFNwhWW
G+YVYFbxnjlbetmKUZ4n3+WggKeVC4zHotk/x3aYKX4jfRmQc5t5BTy3NJAgXauETEpVV3i45uOQ
vlDm4VHkPN0rTjwMpAlN1AlrAAc23hJtSucX0j5fOCy5xISJvTiIeRnNJhuuNh0QwDzorKh52z8S
mBWx887jtdY65oNO+aKg2IrNF7TtmYt3DOEIlciee0uq9A4NljPdeyceHdyZQk39h7iKfAxJeWUW
wroseZFItC5tuAruFtNWk1ODjbyYAcmIzfWZjnDzfZPxaDMBovyiuOC5BRz0rtO+o15dw5pbtU5s
5pyXyx/xum/zUTJ+/s1bpSqGfdivMz/LK6I+uLBE2K47JCMxq1YsCsjxMCwKL8F/DzZdPC2zALKA
3UFx9nmgXVwFbgEEE0O/TiemdAKweFkY99NpVLEoLtBsBmKw5IU/NOyt9dDkHg66kbmTEzM6morB
sOqBebhYhrxl0ahNQULfxcH62m+4L8uAxZydYoM5m2u/uZ7ycjMlAIZjLooVtAMLJVR2y2nXFLPG
zBGeFd5GAQc1d6/leab+U1BdEE/znliXRIKYLaQZAG7e/eGeZET/T9bFhFUq7YtMO33wKhP63tu4
rLQ4jMU6rU5K+iXZnO+ZwcSBHBUn2mZh/bSqyk3cIhMNJhzU9VER6D5f1cxqZGmRrbh56mErIHGz
X7MZjVELkycbJVldcRBgMpoFY5kPVY5zVcvCRibsW5Y8wCEUsKA1q9IOEvo7Vggq8RVS6U2Y2XnH
M3YghjLznTnjYHCOa9Sk9G+KTG2QLiTrLpt/COFiQn9EcEt1ULK2RgDuJE1zj1pWnAYunl/SxBe8
y9xDXpkesYUF9orqdi4v3sti1xWYxVGP02R/tDAfvNWfdfirGJt76hNcHPTgodhq916TH3Br//fx
kxTAg3/RD86KMF5aFRNDL9ahNmB9CmS1lKQQjv+c7AS3E7MDuHRuTEV11OxkwYjQ0dGMx8nCHOZk
7lu5SNJFKM2WwcwdTno7zzHvTSvtpGrBY/13Y6OI6JxaIrrTDJYD4j7l47K5fLM7+PFHY0TW1/Dl
C4U6x7HFHsogd/DxHOhM2GcjfKKP1AJVgLMbwjga+OYl91iHnpM7sSR1D7PdDzv4atLobIec+6dw
Cy0+SUUtJobMGo+k3GL6wOBIPbzUEIsepcnk8zA9tXS5wIYCUD/Oso1Umv365Fc9cId+mCcY/iW7
E7GlLHoLHws5H792FV94kPdSmUl59gDlah9KQbjH5xMsVDDmsTgYDPE78k64c6QyALWZafBwvtkD
njQEjLzdKt8Xz86U3GUanayq377Gr9WKGw1v0epFcuDGeZqzm8xWdKyrnri9sQz9Br9Y1t9yO6fR
umqISz+HPO2sUEg85JjHmH44yc+nEJxvIfaiX0n+MCXl+3HWdVu0mVwsfGddjBZoPd1KHW2y6847
C3CCU4rjIIuHIrYN1Y9nhE9eOuljoes7GXxmrfYhZVH/f/2bOhfL/p7tBhL07qOCIXgRi1v+5ohE
ZDfWAvNlc4j4n/jnE3gc95FkncHlPQvcOrKDH9KTvv2TyYt4IgVPCk3ZzV9vutSjiD6KKyrATrjX
nGh10W7XFrfzNGCmckKSB84mfGfzEF8EiLUKi/abp+YQl01RpZnFTUYDrGxXMn67Zr3+vRom0JQL
vuMVW7xXGb6KL1ILArPvx96x0MYutHCgy2gJs2AF4WAYYuzBOt/TESKx6Q9lMNp+G1Lf90eoL7Ew
Qu8hQ3sAabRAGkdwIo8N1u8dirQyiTmBoAIqfRsfZ+O+WYxP/nfe1vPBqjNRGge2yV+Tj4m/Bwkf
AMBnaWeR9EYIbKY0hf/oMTaJGAeoeL0lzsEOyYOM9CkVdL45qnn529R4lhPClhbPbtGBEn2lNtNc
v4z5SfCF6n6H4b7z1S6DTsG/AJrpnfFFYZGNFp+ySbxrtzb0OdOb5dqv/rejptdbC3W8VIXGt+NI
AX3Wcve3OELpQkikWCp5Eympn5drH1y5GknpRff/hsO16JjKuEzZRpA9PIiYZGVfmwJrDNxiCa/M
qZGn99RZq5j8MuKCnClt1cvPHlr2KlDA0P80KBiDun2GdHcccLFm8ON/HImZFFqKiKtVW+0xdYJl
+uRiaLvOBoIKuQ26VEw66ub/DeajCHENirgu4CgmqdVuMVODqS2+zcyMqur+wyXnazyddfPSCPc/
bfrV1rPquyipphw0mFlBjUAi9pw1sYyw8rUz5FF5iIW3K84w6faYHHzT+Q1Cun9UECIVMR1lyCK4
EA1j6IojVgM4biPhn9CAwHmZ9UDkEMo4gv164u7zWC0NDrPjhzGzSh8POIDpqq7se5Jm+Z5e5eSX
QJtOH1bwfYZjx6RVV9zL/bhPfgfM4toHXXJ/bc6xzluCDRjP2iRB8t0mMMlKnIgv49aEkPMTGflj
Wgn9z4QOnW3s77kXhZqyPJaAV7POfU9MRnCBLuKHgKxmRZn4mPmNJ+AT8o4vo9HgKHCQB1P3rJkS
RQE/xKtdzNBjmtOpenOeh9b0/tW1dOzkHt6Jb7QgX2dKHoyLqkGkI2ikphvXN7zai7PdKO7TdGmM
JZhIhEJTeQfEEbHvD4ZDKN/nEhkzWPMmGXExSEBDXYIAycuYjJa5qu2Luke1ycyguYLU6AK/PDKj
uyN2GZS+BFFwc3lvfY4XZZi0EtXV9It5Qk1HpMdoXBdiawsp4wbiTD0oRylYzQJZ9XOVhqTuwUvA
e74YMFe0GyanQkWeOXCORDbbXy57CBbAymYu6xEr0tk2aNQiOeBvljxc/8DGkZiMNL25IFEMnpNx
/f/N6lUQwlGSMy4xv2QHJBwC86N3SF3I4bJ9RaI+zP7/YPsdxLG7VQUfXOlBN6amZ3ozLUsWRtiK
FgM+1eeS3KxdNQBlHkUQroMwvzpV93krUqI4M1+UXghJz/LzpCTBMC818yFf3Gmda+Kkffj7quVf
qMeUvJ1yiSrtX/f8MPTaPQWOYMXw7KCdOU25K3i13VgJMuHhfAoonSjX/y53pF3QFb/UWBZ16DJ1
CR13mez2vIbtj2CCG7UH++pH0K8ITv9I2uVvMyn18qkULB0AyAi6lDxCugSlQvG26o9mvmk7K9Bv
rHkQm9SgUgstbkCwRImgoBN1me1cLGKc8TULzJ8EBfs/+SzRI8b+N4gEU5GnOq9SHjrwi/BCeiaA
bPJPr1Uol44N5iZj+6Qzby1Kud53UVezxmmTxhUwH5797KprJhoolGQsZLi8btbzOAeM9KYv51nI
88TtEjhHPEeWMiFgtki/0GcXR2zoK54XCRscHwI5CJhAxuPSzKo0k5PK2yk+aexdCfIXgUg82w1P
fd/oSPhLl0fztYbIYzqrBV5+gw7eCHy+E8JpzIwBoMVBoOSvgketYdjeaLQF+d6FFqJr/6ThEFaT
NFYJEx8F5lYtVlyiQenu80Ylx0GtXH1Rmq0f+bvUtyWPrf+nIJ3ijYMNmVjop7LSWNooUbjdMa8L
d9dfLAyZ3XWZ3ge16Pj5RH6l+MC3/JpAHbWBq1WB58JWfJoXAJZ2Fo+NuvhzT5fxejPS7O234FHE
4MnvY7sZgT/Gk9LW0EWYtm+/gxianxtZSfASLafWaKZoCniUK/f8vvxlIkW2Ut48S20/w2dw/qsY
DkIgd9gwbAmOsSJIpZCB4hHNLgxffm3xC2vfohskDQthHFKatM4JMd0hjKiLKlN9xhS7UiqTMCGE
1vYDf5EA5UlPcz8jNvYcHbRzXY5qyipHXG27TT+acdmeCDDpLytd2J8siUdcBXD4/OnpWYu8zO1V
R81YS/1oTBTsemZiPf2xgsymmI3uqNlAqWB1xPTMWuPwGCIynE5g+ojAiuHhoY3Fxs6r2DEx5xLG
eLz3COvB5EN7e5EM7G195NN0ppRZYjpSJhcC5sZckHFdo7lL0PZsr+f2+kMFTd3mV+SHe6VgrZzM
mDQwkkgfDmGDgzBaL93Dc6ffdLuKBlyi0gVBGDHMmw6UBAYJbP4kGPYIlV750wHhoMXRRgkYVA7b
bUc9mll1y9xsLsojUd6YM5abcrGRFg4YWVoXSGm5ztOgkkPefQVH8/GeyzgVTefL72lffX7DGSGL
XkFZnA4k9v5z1rsUQNGbVcVON/byQG7NwJUomHiR9TxdjWFhwTT3iI+FCAki4DF8QFWYPrBHE9H/
7QkLZjJrTGu10rM7geynSf3uOd9ZchEjhhyFURYa3/fCIcBTUk/+Qy+yGFhQXPH9TKz/4b4h6h5O
r50T2BGsCL5w8/ZDMwvREDx3ONgmI8IMP4JUMhU4cjhYxqIXyHdTixoIdWdOHIxydIx3ebgQUqGe
ZUSRrYrOGG4aq9C5sEN64D9mTcTaHaNxdzqs8XVzXq6d/pieNKk3+qRot+Q9dXwz9gzQDJcYexfl
AOQch+pDOqhqF7Ux/w0n1R/66L50sVQOIlo4WrFF9TiO1W5FcoJnmP5/shKfLYecNV3sIVKLCIZh
u8YdXC5pvYBZ48S7Tu3U/vkMGlqAJt4yn4pfzOaTVPYP10i/lpxFhfXJKbj0opN1g1EgQ8fSQXYf
XheyrvIiPbLazBUHo8KMtCgd53gvtxiGMzrEyYsFEA+l/+Rjo952MjfFCdhNSL93v0w3I4JbJrvc
7K5FnsVkmmBvyoOnxQvxPzbLbF6x2iSFXx06ijOCDfqxpswJoh/oPK/hWKmjgufxaEtfFplAGjaA
jDC8oVd5NO2LOw/zWkK6b3412c5H8EibINErNv2lDryOwnLEnNoJhZHuwcM35Mc5UwMOhulqTeZL
i3QuKIiiHAuZFtwK1xiX0Qe/jIyqRPRsocWe1JEk22/OBBYOQyDL2uSzm13d7DN16uR0nAev/eFg
9ipnmBMEyFSwBUaVpVHaQnZ0aC2X+koF6Onul5tG98RQcoujh1kwSeGV4ZEY69GwzaxM/rEbLVTU
rcabBqUSv6x4nkJwcrYRO91d9VyO8hn9N76IcmnVgRxParOrbtp0M4qwYx0gnesT2BCxYA+xtW14
ZHa/hxSIZH7szZ5NrMHlKv7LV867GiiuNtTeKA3mYtrRydm0decnt1rNQKGVG1LoA6t4bH8HoMzm
Zo+duFubVoyy+Md9aWc2eVWzrICDsNB2HK3gbxrKh/nv067UG/5y1SxWHCRKVkipkUvXt5kfb4lE
ewMozLC4qcWX1RYBkqb1E5G/7KQ3fkyqozvkgclUrZEG4I1VYMgkD4Ypb9WD/S9Odk6Vi7JcJisk
2+1Of1sirIlCe6HgwFcaTqcUu1htRcIOOdoyHFpeQMLB8IgRPkWp0HEMsE+L6LEjD2BFLCd2JlDN
RAXA40Vr8hChTHvZAyR5agQWGRIv+Q9MczAKdfNBwJWoSBaxvN92pWEKq2DiBOBfBTnfC6NAi4sD
BmQHQP/zy2JT8rimIyS+28LiWXMBoavGQq+Qzkxks8KcM/TqcVxGoYzNHnP5ogx5pN7aovb4yNCX
5dyFuf/X5luc8LKDWpEujNRXJd2P1J9Fop48jm27eS3Fg5k6IKVumLCwc+qJjYMAlqFMqnDp0U+v
86P4YR7ki4CcYgwGrh1wu2PAfCLuB3C6u+O/z0avaZVdTpaI9F67/ZqOWy69E6eVhmm1IJ3LTgI8
VBk7N5WoMmukZkTb8ef5cM/HXZPKo/wNp7Gc0OXlmtZFqcewxLqinT2N/C1udqULj3PrttsGP5PS
hn+S5OTQFIqBS9xrrTTXJ04j/BsqFK0nQcZRzKLyewmrSb/Tz2jOX4e2w9bJYTSJCHbd0oc4pE/n
oORv3p0Jlkzm42EiKw6S6F4D46Y4tj6RlW9XaMCB/2yo9gEwYKxGRXLg069szVfJFSTFfFceZw1c
b88rj/Aw5gaBpUT21/tvlnxyAeM2yKXt+4PuFLCTgBQpCPyDdNkjjjX9oxaaRDBM2b6nVJ3csT83
2TVptrUchvgeBiYMLU/D/384/67wfVBLfbr7nYBn11Lrk3k1wyT4KzJYiceHWemjvZw4d1IqbaC+
sk5+QdayGC3lpVuG9C5Xx6gN84xBdXFqxHfSxt5oQgfFyiDBwRFpn5pcm9t/EKJwxFZpzrmOd8En
N17KJMIUnJZxBIm8qtebKxj3iHTG1bAHqL9s+UjpF77p2OFCDdR6zKRPflxlrC0cWFxzL2KZDnRe
hvoNbWDltyctcpQoEgXi04o8LQLioDMaCi6BFmF/2ARISpAEQk2q+61xjmZHHZ/9V4jfMP+gqx6m
sRlfZ4Ix/r+nPD1gk6Ni00fQyM07XFVRUp7qYEyR3NG44WlFHzs993AE5hepx7lCfEQ4U5TFK8hQ
e7UwHy4OfPp/V4k4EOEPMKOdQjK+O/MY6iBaSZ7ocdhzCimAYsZspb5bxjD60oI4lVWw7XN0ouoK
AFj86iiFUGpqbdu5VkihXS/uYWEFEpy35/cJ4BXMBCQ46BgRIy6PaVVRaFWXI+uTqqb8MKwUGbsz
XJYA7SW6OxuT8+KojBN35svUPfXuHJbsTCOv11ax7jpSS/je9Vjer3MxV4YFmLyg1s4pJsoC0KSo
tWtF6qZxtQB0xE1BvQ2arJbba492GIgr2IZ8i6vkDVFWOhSzAYYNTaEsdxX/tMijdWyjpM962swJ
WiilZnklC2MCyT3dNZ5SBRzWU1zjf8CtGzVvyW76RQxCQDGhsyzatboaHHAsUSYzfAHLdB09Y2hA
ccJ9x9Gu3V3eJ32ph0KyqSW90iPlgwtoljSzgHYh4BNRhsuPS96Ge4prx0swT1JTRBOzCBAg0tZm
+wmyCCX0L+0BGxJp7eHnyU8pN65cJTuC3hryJ3CycbLW4kitKFZs1N1CoqFHMXAYX0iHBIGLDxkf
Tn7xhOOwjRTf/d0gIB3fm3q4bS0OZSwvNH5k1VQ0MMC19BiwPk771ovb3X9fN+zm7B/baB319dLy
BAtWgUZjGRwFUI6DBUQXOiAUzeuJCLvykWlhs1FkqxUKNt+bpjTVy1Np3p0UrWXLDkvx5n4IM7Ey
VE52ky4gPxQLiAjyHO5nTydbIPmWOym+mnYrUTk8znW7mkmdGIPxssc1Sff4W5eR+vA5U0rgV8Qo
o1bYJMP9Tc2EKoFpP7QhR4c6r6RMxTadk2DGYx6vT7E5yvHqBcXC3jkd+L/X2w+8Gvk+Twi2f6TE
sA8mgSNft/13/B+eFgy5lHvv/WpCharDiVAj0Vz18YySf5g0187Hzf9T9Ss/JZVhJpZN+0LcaVt3
33jFq3jCxMiy9dGSfgt1hktdgxc+AmBs17BmBvzK9fb/MDIMqKdjEuAvitF+oodgx515tGeQKEUm
Top5U+B8ym3SDxrF4RVt3PrIIBAPEDSoVO8I9Hion8UcXHbNRQsfIaQcXR1USa4UZMeci1ws94F2
8jL9tvJTikgh/DBAJM+nrsdZ1xbdmt7NUsgpLDQFQPi5UTIKQQswZR0pyGmgulC99M02pNVKernP
hw02LeOdVcLGmrAdaCQEBFo82+q1y9v7aO6p2qsX83FLfLjuNX8+qZxJhr2ca8LjptT7XGs0JNCh
7N7b6Q4cSHifGlr2PgAH/18hbAEEWV1ycbqZlqimcy03L4+JK6PWt1VTR3//XDZ5VIrdf3da+/mT
OzU7VU6u0AHOYaxShI38UZcOaT24bYPj54gY5Su4JrxI+XO3BOc4gfYJfXOYWWSVFhl9bWpYw4jA
q8lc2ArembMH6RXjFpTZiJHVPstOeYbPGvoplwsbobZF5M9+h5dQ9PkVXlpSnnjvb+DIlzbHzfjB
vMp/W+oIK9RcncKQVarWeEvCn0Gg2OF4OxrR8MyKaI2sbVZfQKdWsKuCCd+G7IwRS+28hnPN278K
GF9+B7JtPZ90L3c3hqCG1S0PfrySqEdAimMpsOkoMIV27C8xQaI9p8wO2m4YtG0tkmW72MwFU61g
B3UvN8kF2fUjkt38XLiOlJuXbpxvD6hKrTYvgdferxzI5Vf9lfna19xNdPHhOIRoStl8rdrlUf69
NSvN7rPg8zdfmDeQGVT6Tjratn0aJuS1IvF0lNIYcw/Xrnx3GxD5KQ1cURbHkT7VR6P4V+MSQaDZ
0fbCuIpWXuZf4ueS9VygYiJ4BIzR4BHlSYj5oTp2rdSmhJVO8vPZvsEtKAcIxkyzJICpL2NvSk6P
v4QAmua9hOytqNre+e3CRtmods4fuQGFyRZBP/KiKLShCh47YpIfhMlheKd/0A5aU/lZoTmQCaSS
I9UD9F6bIoJnBXwE+YbcM85OTpOySozWi09BL7z4GjiH/VsfoA/gzZ/ienvwApDi6ya9SQGec4Hd
2HyMmwUqSGZM3hPWW3W376C/3fgRF+IJhyahXw1wrLJx+Nyly2b4zx9FWKFnt+4vJbvbH6FIcM8I
NGC+Vk4CkO8xII5a6gwTtwG7rBUJQQRyXaZSAFDuZBMIueeA8bkVi3cIivXNjDHCD3OS2hhG+DgB
7L5QR7QrmAvxUHNLLlru/43xEodgbRWhzk0KJTfYGrEyGEr+RFEWkp8tghh/XVrd46TAbLjWMudb
vfHHZfua0R88T5EgpwrXU7yh+4BYzjDvC//6kLaQe0B6rPmWiRi/OWxqyMmvkAQtTIptpX8/WnLZ
6KBZ4maPf88s7kz1x+CZsOqz+SdDp7woUlsVakkJho9RLpsKrt1BM3ZhSaWE3kX5udKlYET16ppp
0TttA8s+uuBq+vHPFsZxY35+uHD4MqFsnThICT9naoa8zX0GyJSnMt3iL/Fgk7c1ViiCCcC+G9xW
t29CzGsQpV8GEKTSfggV0upMf4cq09JMdsFENqYk6jFMIHgsm+KebB3R64IF6+e6z9JLm4SLF6Wr
Vujpd+TPGwpZ7HcsZOmc0PMp/RQdMTPbtme11yqP7QwqY61hTwopX3ws1zEEq9GNMJnDjsZVXEdM
03VnsuYf1KQzUXdCkf5WuS/L9sFZLaeGWFh8KXDhyOk9KgkZg6agrDVdiyn1QaejzyHukCynXvhm
pSjJJIvBEh/FSC8Qyn0N74/8/XgwO/J0edb1JdGrpOXnmsR7LfpTKYn9goUEKps6o9MIXI7vbhA0
MgSCPXMpVNiVEVZ82stl8yonuLnP0hGUOT9wVgIqgaTXmMfiqbijjD4bpsl6Nh7Cs7xZ4ny2Pedb
QdCrDHtLabqArCMZwnBoTQvuaabcuyL/nKJd2wKHnB4A6+liHFYMmZmh/DW9K3db9EZqWhbTduDA
ZzEMW9b82q3GDRp1PRSQZXviYgHb5qHpQyGjGgbsEGVZMqE7JjRIgwEX+lvE5lXsiWS6pS+2mdlA
FJw7ysxYyp/IWk/ui69TrtB/3Ni/JtQXKPqFSkbyJjZxfJBfJzmYMKYH7U/TXYrQLZbJgOrhetTp
U5G21UWKm1UXazjLdXmGiUjjgah3OFjvi9N22QRZUtZMTGj6Y+fYLELI7J9pXtSQn472f2mcGiha
3aomE7e7i/wWZwg93adMqajqkO+vEnayAOzo4Q3K99C3r2woM+1wsI7QBMogxvOOQGXFkqbF8EVg
UmFAmrBIhIT7weAjXnpZXRExtPOFjQ23hCyeqEvfZlhQusAOBH8vqR0h2gOlmQT8fFqcaG8LP1Mb
XYskAcKyW2+pZPNYfxHmYEJLLLcfnCVi+qc6QpRxboy9BxhvIUW0XCVhgTTV6pBCHuBJam8fHSA/
psmkl5f+3zz9vcOJQd72e+ECjGa2yLIHBE8V6ZXyFd88eSnPWvIRZsRGuMgHJMDhRBjObKbCFaxz
wOiIDTyY+/pRjRNw3rHqhSy49//3XmzVRdsFTi83bSEGlHcr9rcU+DqPp8UY41YDafrppF8mY0yy
EXdWDicVMhCmGcN8mr8bT+LLDz+q3y60Hw/kqvMhlihZtDmG8kwsivwAwcKeowJwg4/EVLUWFsCQ
YWdmjfWyjfE0ohLzb5qSRQ2aAvgZ9ZA5lQ57XkR4WpiAmIm46EgHcevJIw9s35On6RqUQWzME1HR
XGxEeXAu46nm7a6uYQR4wrbLAxDt0+6zy63jjuSBQEdFhStub2ZGyx+wSkJVs4vLDp0Ji2dALbG5
dCwg/H3MuBGhZs3I3J5tfQSzdUA19yBlsY9VQXpWEwt4dfKzjPdt0EAiksz2zxsNE2W5AJPb+UiK
HIrvhVW/1LrKBOiPZc2lsbGdqT6xY5/SrCkJXjPNDkVQjvcMQQ9reKWRe/46De8Gp5w4bMBg9kEJ
PoNc40w3ZotuhdK5sxOjHSC11/G8HcKRvWxMH46iZlzMo6FafO+f1lg/HlIO6UOLC4Vx4YRRO2Oe
PZyXdTM2V3hMU4QUWy5obBSoWCsiAni8D6Xql7AQ+sz8KFWX17A8brJhjVM/nLBQeycDDQpIG7SK
W1A74e0K/VO4LCpbOdzHQ911zQsFYTiIqFall68yUqBSTZySGSqwpMDnRXV9Wrdi3mBllS7cgB87
uDIsorPLoQ2fCLmZk4BMgDkRHMCbkJVM4HQhLmORFI334T6quRZ1l+0XcS0q0XDQsxWCD9Pd5dpr
SxpPIvzsQAPtPKVbEgDGBm2nx7akZkYmNnVQt4a1WZHwFYdUadSGAWRriZJ0BRPaYMhLsNyt1VRW
zqQWECOkOKsebILNy9zpOj3rJkPdFAAFOIe3oLQp1zExkzDElDZNinNWBIhefKtPb2J8TqAHKzf7
q0n+ELNJUCse0D5Z/hPpx4EdBwooyHkH/5bmLy+RKTHqowP3mIwk/samXMUlY21XqKIPZV7Wwn0L
/0Y8Kqo6Zjdel6IG9hGXMx1izj0BLlF0OKR7QZ9Tg4JvCK6oAyz/Ti36lpDXGCgIHwm5zGyRrKIy
db8HpZA1feb3BE10MZC5d/OWA6cxrWtP85AzvtCDOEvKdPvBV3tCKjLOxa4T0IE18r0xCCJjD83k
V3B5E4i1PFMuCMqfUCohSZeT/d5WZOxzz0kmgoj7nWfepPdrc7jDyJXweE6fPA04dMm2Jhr/y6eH
nePpmiGwNgroVYlyvXaNxDJOIvxAGqR75eOXdpkm2obbZNR8Ih/Ucc1StHCbxt7htMLTwNpr5qvv
un9au37XLhuaz64myA95N5iloG47KCR0hLsSuHa9MsjjmylhneiyglAixI087U0bSngrRIfMASxv
nq3RqGcKhFsWUl4WHt9KwBPhkY6iLQFIH2+vzT1IfoYxU4nFVK66ScbbOOkuKR75/4WLqkH07Qxe
uuN3KlqIOjZ7Pb5cJxz0KK2P6g1LJ8w7C3JMM5245XQd+IPbf1BBS/mW4/myQhgUynDq8z14GX4z
2BCwA6gztin+ZPzKjJPjczmYVmpJQUYqro+Mff8iO4NRr+SVVWMdFg9M2Gr1SyA4MIbH6AfdJMJT
ayIrDzb+w8+JAgc+tXKWckvwvzIeXw8R5QU3nR7Od4D1/gKd1MieW3xCuqEwaYWkqRAw1hntEPfh
z2T5zsWMKg03RJDjgx1JPlM9kGP9Np390KPeVZjnNBvlej9IYc0/nLmiTW///GVDh0KlWq3irIzZ
MsB//swt6JwrvQie3Lus1rvGPemDIhmP6978DUnUbSgeOMgScu6HTPk4Sw4b18QsD2YdABCWvqjb
v+EF5EQzncGUvB/xay6MWFCH8p4IuApkEbeV3oyptk+5aZ+gRVn61jwYr5zm/Y/W62uStJuF0+eG
OPvhdlOlfrgIFIZTNqkyDMpXB7e1cptdXba65FYYSHLGqY1Y6LAtrp94LDPpu78XdW5tdK5CPtxD
cEmwpjIPafJStBbUExEaucbN18xAUKCLb4I6ftyOMdxLlVIblIpJCrJGsCB8axPieD4wcaEdKlRl
iztJsZjiQKHoNWbingEVQjqvxXgJxLw5wE8xgjUDVjMnxZMZoUt/E05vEK8fShpCfw8FS8IlffBZ
1Ah2PrEUK54LWfNC/Axygx6cv6NkRP+ZKpi0WM/NrBbVG9wun74/3/BylFtpjSay6IjA4jLlQPGp
HkutIDYRzU6Fk8sW/Rz71F+2PRWrWX1OatASLp9qHpeU0k/lmWk+zdSLDfEGvDOz+IlvB4pvPDM7
ewS9ZMmh9KLI5GoCTXrdaVS0AcnJ73J6ZkhdZ9MRp4uujb9LCmdyKYybN8jBxhGT8te+2gbi/acL
zHLMKTHfHDw980R7px0MfG/Wt6anfiZXBCISq9mpC9ACbDJAmcFZSMmdWySLPA65VXLkYUvWp2ld
k/EXDuMBVW1x2+85aPa/TlLk5CrkbjJkmBCnBFxoNnlQnshKmTAkHrEkDBLf6Gtct4ZKtaNpidxw
JKauxVqxKPp5FmnmN8M7VoeJu/Zf+wuQL6zXRzr5VO8rznLIm8pXX5u8Dz3wTjBoXjTBaWOxx9/H
OdEiTuVSGwQguejlTJuAp4X1SWhFslzyr7NOSXfKEFJ543uiUUA0qLB5lLd2WwzS5LwptxdI3P5M
K/0JlgIQzS15AFHAVXw93SuCqP5ZhekniU65gKdyUQXTk2mVzO0yqwg4hIUmKZ35cTdOWQPCPzq6
gmH7F/2nGD9PBctBBuaXOTunOccUiCH8WAULzHoA4TbOWL711x+LUIYBEX8Vd7xVI/VjZzz+pf/m
hAFryp9b4PyOnp5/WNg79IhnAayqMxQPkJPWgmsJv9/IY4baX2xN+h3oRqz+jXtCHF8RFBSKuQoS
I2oKFSudOtor76nIH5oyMo7T5rpjizcMfwINRafYlp/hyc3eLxIwmPKoCKWgN9V85I/sIkWAk7Ez
gZhtnRJ9Ga31jdDukXQB4lULotzSdO2vKbm4yul7303DuhrWHY68I1zObSrPKB76c8qbBzIadnuE
VcbrhNlI7uzGAbrdSg45JjQmGJGOG0rlRQ40y1fRb8XHDui2qnc1sKniqVIAQsTrkH9HlEboeVnv
Z/6mhj3nMHNx6Tu+1W6ZrgY65dNs0uM/15cUMdqvMmOWy7LAm4VGaPFXFxP2f+UOOUMFfxxVoxzR
QWS+vmKMsN+DaMbBVZcb5qRUAtN4ve8cxjcZ8uWmcjpsv3dJzXWVEn1yy2hrF/3ImWNVtarTBebE
E1DmBwHUAjOrXuW7h4ica72vJSXEGomvHQLOsvcltrSmi/2GBsT6Q3k0xzUgblGg2sFWZFlzB3sv
qSAvEZQo1xAbtxu+pk7C1pyrCQCyGC/AQb2FlivjQNsDmw98P7n0UJG7BxdpB/adkm/094X1DFT5
4U2JCmoGN5/E0GJAtkbdr4f23nhImJLizBvRidPiXGu84ONfETf2rDSrEQDwFcCy4om1RaaucCnc
L+tvbQbkCv2/MbAL5jF2EJQrWlazE3PpdGNPURI9WzaZD5AB6kRXAOtGhypOyyARfUsOBRlauSuU
iBFDTW7OXqfvcPaGpvVuv3rWHbOWtOpig7jSVBbxnrdj6lsxOOwWDd7m35W9JdiDxQnHe1UF14Kl
ClV0KCSrMSd2sqnd9G+D/+V5oaYrQewCEItfpOEkhDFFF6BX1CDrUTei7HymqA5ivWF+U1iND/Dg
MUYM60GNyyTOtT+GXAf4oq6s31idUd1y/Vnzxh89AATSedJreDA1+kSm3MtT6KG8OfA3r7bnT2zf
C7UHKuPrlYWbDLYV0S+ik3nx7I0zvScGiyQINQsFJiPnY3f16ztcrRfK3aJVG5ExvCudoq3AlmPt
WTS83x3orcAAXnAguA1WXlSVflLJQnBe+tubWwe4QQxgEeAJaweZS1YainrGQMCQiNJ5Ny1AaLKt
4wxxWJ9g1hIGK5YPsHk4YOsNXHrrwcoODzH7etAC0iMRizuam6KkWDbXo16VvrIEfuEnqEk5xesJ
sJD66Etjmu7TNsNBozs2uiNj1fsohyT2WwoqmcNfhrHLtVLQLKoVGhM0h7k1lHUlUqpDsFTjwNHs
/lX29e8UdbLVuI8ULfIBWCgjc682uXoxyy608l7nEUNvyCJdoD+RwhkgaAOQBGbVLOfusJ2wZueW
3bxjs556qKnMi+iuPBZUtyudVxJ7mK9jm6qiEdbphZLDyhKrM7ky6oShV/sQtcAQyAtWjPtH7Utk
7MTMgl63M7F6rKpFjF4RvgUNA8kvoGTDIcRk/Vt4QrKk+DGUTfZu5kw0wI/IYGbQO5LCob8VuhVY
Tl6zwGBsIj2cc8Qoz4RRKr3aNpqucjbDyMwBiVpr7BJzhA4xd+xkyFvYZDavglUFGOgL8Ta4XLIa
o8Gf9E12WoUIUGsBAqHAC3mmHTkOEiqgwPI4WZ2bgU6fPjA7QjdifJWGolQCCNlRdUrhpFdqo4WD
P3ZPljpv3DZm4Cr9TYD4+eE0yUR+4g==
`protect end_protected
